`define BINARY_OP(out,a,b) notif1(out, a, b);
`include "../.generic/wire_test.v"