/*
 * Integer wide range test
*/

`define WIDTH 32
`define operator xor
`include "range_any_width_binary_test.v"