/*
 * Integer wide range test
*/

`define WIDTH 32
`define operator & //and
`include "../.generic/replicate_any_width_binary_test.v"
