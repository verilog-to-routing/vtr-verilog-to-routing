module test1(input a, output b);
    assign b = a;
endmodule