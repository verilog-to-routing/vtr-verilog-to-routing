`define BINARY_OP(out,a,b) nor(out, a, b);
`include "wire_test.v"