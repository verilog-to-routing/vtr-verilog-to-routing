module top (input in, output out);

assign out = in;

endmodule
