macromodule my_adder (in1,in2,out1);

input [3:0] in1,in2;
output [4:0] out1;

	assign out1 = in1 + in2;

endmodule
