/*
 * Wide range test
*/

`define WIDTH 3
`define operator xor
`include "range_any_width_binary_test.v"