
module top (
    input wire clk,
    input wire rst,
    output wire [1:0] dummy_o_out
);

    assign dummy_o_out[0] = m_axi_noc_rready[0];
    assign dummy_o_out[1] = m_axi_noc_rready[1];

    // AXI interfaces to access memory
    wire [0:0]                  m_axi_awid[0:27];
    wire [63:0]                 m_axi_awaddr[0:23];
    wire [7:0]                  m_axi_awlen[0:27];
    wire [2:0]                  m_axi_awsize[0:27];
    wire [1:0]                  m_axi_awburst[0:27];
    wire [0:27]                 m_axi_awlock;
    wire [3:0]                  m_axi_awcache[0:27];
    wire [2:0]                  m_axi_awprot[0:27];
    wire [3:0]                  m_axi_awqos[0:27];
    wire [3:0]                  m_axi_awregion[0:27];
    wire [0:0]                  m_axi_awuser[0:27];
    wire [0:27]                 m_axi_awvalid;
    wire [0:27]                 m_axi_awready;
    wire [511:0]                m_axi_wdata[0:27];
    wire [63:0]                 m_axi_wstrb[0:27];
    wire [0:27]                 m_axi_wlast;
    wire [0:0]                  m_axi_wuser[0:27];
    wire [0:27]                 m_axi_wvalid;
    wire [0:27]                 m_axi_wready;
    wire [0:0]                  m_axi_bid[0:27];
    wire [1:0]                  m_axi_bresp[0:27];
    wire [0:0]                  m_axi_buser[0:27];
    wire [0:27]                 m_axi_bvalid;
    wire [0:27]                 m_axi_bready;
    wire [0:0]                  m_axi_arid[0:27];
    wire [63:0]                 m_axi_araddr[0:27];
    wire [7:0]                  m_axi_arlen[0:27];
    wire [2:0]                  m_axi_arsize[0:27];
    wire [1:0]                  m_axi_arburst[0:27];
    wire [0:27]                 m_axi_arlock;
    wire [3:0]                  m_axi_arcache[0:27];
    wire [2:0]                  m_axi_arprot[0:27];
    wire [3:0]                  m_axi_arqos[0:27];
    wire [3:0]                  m_axi_arregion[0:27];
    wire [0:0]                  m_axi_aruser[0:27];
    wire [0:27]                 m_axi_arvalid;
    wire [0:27]                 m_axi_arready;
    wire [7:0]                  m_axi_rid[0:27];
    wire [511:0]                m_axi_rdata[0:27];
    wire [1:0]                  m_axi_rresp[0:27];
    wire [0:27]                 m_axi_rlast;
    wire [0:0]                  m_axi_ruser[0:27];
    wire [0:27]                 m_axi_rvalid;
    wire [0:27]                 m_axi_rready;

    // AXI interfaces connected to NoC routers which represent DDR memory
    wire [0:0]                  m_axi_noc_awid[0:1];
    wire [63:0]                 m_axi_noc_awaddr[0:1];
    wire [7:0]                  m_axi_noc_awlen[0:1];
    wire [2:0]                  m_axi_noc_awsize[0:1];
    wire [1:0]                  m_axi_noc_awburst[0:1];
    wire [0:1]                  m_axi_noc_awlock;
    wire [3:0]                  m_axi_noc_awcache[0:1];
    wire [2:0]                  m_axi_noc_awprot[0:1];
    wire [3:0]                  m_axi_noc_awqos[0:1];
    wire [3:0]                  m_axi_noc_awregion[0:1];
    wire [0:0]                  m_axi_noc_awuser[0:1];
    wire [0:1]                  m_axi_noc_awvalid;
    wire [0:1]                  m_axi_noc_awready;
    wire [511:0]                m_axi_noc_wdata[0:1];
    wire [63:0]                 m_axi_noc_wstrb[0:1];
    wire [0:1]                  m_axi_noc_wlast;
    wire [0:0]                  m_axi_noc_wuser[0:1];
    wire [0:1]                  m_axi_noc_wvalid;
    wire [0:1]                  m_axi_noc_wready;
    wire [0:0]                  m_axi_noc_bid[0:1];
    wire [1:0]                  m_axi_noc_bresp[0:1];
    wire [0:0]                  m_axi_noc_buser[0:1];
    wire [0:1]                  m_axi_noc_bvalid;
    wire [0:1]                  m_axi_noc_bready;
    wire [0:0]                  m_axi_noc_arid[0:1];
    wire [63:0]                 m_axi_noc_araddr[0:1];
    wire [7:0]                  m_axi_noc_arlen[0:1];
    wire [2:0]                  m_axi_noc_arsize[0:1];
    wire [1:0]                  m_axi_noc_arburst[0:1];
    wire [0:1]                  m_axi_noc_arlock;
    wire [3:0]                  m_axi_noc_arcache[0:1];
    wire [2:0]                  m_axi_noc_arprot[0:1];
    wire [3:0]                  m_axi_noc_arqos[0:1];
    wire [3:0]                  m_axi_noc_arregion[0:1];
    wire [0:0]                  m_axi_noc_aruser[0:1];
    wire [0:1]                  m_axi_noc_arvalid;
    wire [0:1]                  m_axi_noc_arready;
    wire [7:0]                  m_axi_noc_rid[0:1];
    wire [511:0]                m_axi_noc_rdata[0:1];
    wire [1:0]                  m_axi_noc_rresp[0:1];
    wire [0:1]                  m_axi_noc_rlast;
    wire [0:0]                  m_axi_noc_ruser[0:1];
    wire [0:1]                  m_axi_noc_rvalid;
    wire [0:1]                  m_axi_noc_rready;

    genvar i;

    generate
        for (i = 0; i < 28; i = i + 1) begin : gen_kmeans
            kmeans_512bit kmeans_512bit_inst (
                .clk(clk),
                .rst(rst),

                .m_axi_awid(m_axi_awid[i]),
                .m_axi_awaddr(m_axi_awaddr[i]),
                .m_axi_awlen(m_axi_awlen[i]),
                .m_axi_awsize(m_axi_awsize[i]),
                .m_axi_awburst(m_axi_awburst[i]),
                .m_axi_awlock(m_axi_awlock[i]),
                .m_axi_awcache(m_axi_awcache[i]),
                .m_axi_awprot(m_axi_awprot[i]),
                .m_axi_awqos(m_axi_awqos[i]),
                .m_axi_awregion(m_axi_awregion[i]),
                .m_axi_awuser(m_axi_awuser[i]),
                .m_axi_awvalid(m_axi_awvalid[i]),
                .m_axi_awready(m_axi_awready[i]),
                .m_axi_wdata(m_axi_wdata[i]),
                .m_axi_wstrb(m_axi_wstrb[i]),
                .m_axi_wlast(m_axi_wlast[i]),
                .m_axi_wuser(m_axi_wuser[i]),
                .m_axi_wvalid(m_axi_wvalid[i]),
                .m_axi_wready(m_axi_wready[i]),
                .m_axi_bid(m_axi_bid[i]),
                .m_axi_bresp(m_axi_bresp[i]),
                .m_axi_buser(m_axi_buser[i]),
                .m_axi_bvalid(m_axi_bvalid[i]),
                .m_axi_bready(m_axi_bready[i]),
                .m_axi_arid(m_axi_arid[i]),
                .m_axi_araddr(m_axi_araddr[i]),
                .m_axi_arlen(m_axi_arlen[i]),
                .m_axi_arsize(m_axi_arsize[i]),
                .m_axi_arburst(m_axi_arburst[i]),
                .m_axi_arlock(m_axi_arlock[i]),
                .m_axi_arcache(m_axi_arcache[i]),
                .m_axi_arprot(m_axi_arprot[i]),
                .m_axi_arqos(m_axi_arqos[i]),
                .m_axi_arregion(m_axi_arregion[i]),
                .m_axi_aruser(m_axi_aruser[i]),
                .m_axi_arvalid(m_axi_arvalid[i]),
                .m_axi_arready(m_axi_arready[i]),
                .m_axi_rid(m_axi_rid[i]),
                .m_axi_rdata(m_axi_rdata[i]),
                .m_axi_rresp(m_axi_rresp[i]),
                .m_axi_rlast(m_axi_rlast[i]),
                .m_axi_ruser(m_axi_ruser[i]),
                .m_axi_rvalid(m_axi_rvalid[i]),
                .m_axi_rready(m_axi_rready[i])

            );
        end
    endgenerate


    axi_interconnect_wrap_24x2 #
    (
        .DATA_WIDTH(512),
        .ADDR_WIDTH(64),
        .STRB_WIDTH(64),
        .M00_BASE_ADDR( 64'h000000000 ),
        .M00_ADDR_WIDTH( {1{32'd64}} ),
        .M01_BASE_ADDR( 64'h100000000 ), // 4 GB
        .M01_ADDR_WIDTH( {1{32'd64}} )
    )
    axi_interconnect_wrap_28x2_inst
    (
        .clk(clk),
        .rst(rst),

        .s00_axi_awid(m_axi_awid[0]),
        .s00_axi_awaddr(m_axi_awaddr[0]),
        .s00_axi_awlen(m_axi_awlen[0]),
        .s00_axi_awsize(m_axi_awsize[0]),
        .s00_axi_awburst(m_axi_awburst[0]),
        .s00_axi_awlock(m_axi_awlock[0]),
        .s00_axi_awcache(m_axi_awcache[0]),
        .s00_axi_awprot(m_axi_awprot[0]),
        .s00_axi_awqos(m_axi_awqos[0]),
        .s00_axi_awuser(m_axi_awuser[0]),
        .s00_axi_awvalid(m_axi_awvalid[0]),
        .s00_axi_awready(m_axi_awready[0]),
        .s00_axi_wdata(m_axi_wdata[0]),
        .s00_axi_wstrb(m_axi_wstrb[0]),
        .s00_axi_wlast(m_axi_wlast[0]),
        .s00_axi_wuser(m_axi_wuser[0]),
        .s00_axi_wvalid(m_axi_wvalid[0]),
        .s00_axi_wready(m_axi_wready[0]),
        .s00_axi_bid(m_axi_bid[0]),
        .s00_axi_bresp(m_axi_bresp[0]),
        .s00_axi_buser(m_axi_buser[0]),
        .s00_axi_bvalid(m_axi_bvalid[0]),
        .s00_axi_bready(m_axi_bready[0]),
        .s00_axi_arid(m_axi_arid[0]),
        .s00_axi_araddr(m_axi_araddr[0]),
        .s00_axi_arlen(m_axi_arlen[0]),
        .s00_axi_arsize(m_axi_arsize[0]),
        .s00_axi_arburst(m_axi_arburst[0]),
        .s00_axi_arlock(m_axi_arlock[0]),
        .s00_axi_arcache(m_axi_arcache[0]),
        .s00_axi_arprot(m_axi_arprot[0]),
        .s00_axi_arqos(m_axi_arqos[0]),
        .s00_axi_aruser(m_axi_aruser[0]),
        .s00_axi_arvalid(m_axi_arvalid[0]),
        .s00_axi_arready(m_axi_arready[0]),
        .s00_axi_rid(m_axi_rid[0]),
        .s00_axi_rdata(m_axi_rdata[0]),
        .s00_axi_rresp(m_axi_rresp[0]),
        .s00_axi_rlast(m_axi_rlast[0]),
        .s00_axi_ruser(m_axi_ruser[0]),
        .s00_axi_rvalid(m_axi_rvalid[0]),
        .s00_axi_rready(m_axi_rready[0]),

        .s01_axi_awid(m_axi_awid[1]),
        .s01_axi_awaddr(m_axi_awaddr[1]),
        .s01_axi_awlen(m_axi_awlen[1]),
        .s01_axi_awsize(m_axi_awsize[1]),
        .s01_axi_awburst(m_axi_awburst[1]),
        .s01_axi_awlock(m_axi_awlock[1]),
        .s01_axi_awcache(m_axi_awcache[1]),
        .s01_axi_awprot(m_axi_awprot[1]),
        .s01_axi_awqos(m_axi_awqos[1]),
        .s01_axi_awuser(m_axi_awuser[1]),
        .s01_axi_awvalid(m_axi_awvalid[1]),
        .s01_axi_awready(m_axi_awready[1]),
        .s01_axi_wdata(m_axi_wdata[1]),
        .s01_axi_wstrb(m_axi_wstrb[1]),
        .s01_axi_wlast(m_axi_wlast[1]),
        .s01_axi_wuser(m_axi_wuser[1]),
        .s01_axi_wvalid(m_axi_wvalid[1]),
        .s01_axi_wready(m_axi_wready[1]),
        .s01_axi_bid(m_axi_bid[1]),
        .s01_axi_bresp(m_axi_bresp[1]),
        .s01_axi_buser(m_axi_buser[1]),
        .s01_axi_bvalid(m_axi_bvalid[1]),
        .s01_axi_bready(m_axi_bready[1]),
        .s01_axi_arid(m_axi_arid[1]),
        .s01_axi_araddr(m_axi_araddr[1]),
        .s01_axi_arlen(m_axi_arlen[1]),
        .s01_axi_arsize(m_axi_arsize[1]),
        .s01_axi_arburst(m_axi_arburst[1]),
        .s01_axi_arlock(m_axi_arlock[1]),
        .s01_axi_arcache(m_axi_arcache[1]),
        .s01_axi_arprot(m_axi_arprot[1]),
        .s01_axi_arqos(m_axi_arqos[1]),
        .s01_axi_aruser(m_axi_aruser[1]),
        .s01_axi_arvalid(m_axi_arvalid[1]),
        .s01_axi_arready(m_axi_arready[1]),
        .s01_axi_rid(m_axi_rid[1]),
        .s01_axi_rdata(m_axi_rdata[1]),
        .s01_axi_rresp(m_axi_rresp[1]),
        .s01_axi_rlast(m_axi_rlast[1]),
        .s01_axi_ruser(m_axi_ruser[1]),
        .s01_axi_rvalid(m_axi_rvalid[1]),
        .s01_axi_rready(m_axi_rready[1]),

        .s02_axi_awid(m_axi_awid[2]),
        .s02_axi_awaddr(m_axi_awaddr[2]),
        .s02_axi_awlen(m_axi_awlen[2]),
        .s02_axi_awsize(m_axi_awsize[2]),
        .s02_axi_awburst(m_axi_awburst[2]),
        .s02_axi_awlock(m_axi_awlock[2]),
        .s02_axi_awcache(m_axi_awcache[2]),
        .s02_axi_awprot(m_axi_awprot[2]),
        .s02_axi_awqos(m_axi_awqos[2]),
        .s02_axi_awuser(m_axi_awuser[2]),
        .s02_axi_awvalid(m_axi_awvalid[2]),
        .s02_axi_awready(m_axi_awready[2]),
        .s02_axi_wdata(m_axi_wdata[2]),
        .s02_axi_wstrb(m_axi_wstrb[2]),
        .s02_axi_wlast(m_axi_wlast[2]),
        .s02_axi_wuser(m_axi_wuser[2]),
        .s02_axi_wvalid(m_axi_wvalid[2]),
        .s02_axi_wready(m_axi_wready[2]),
        .s02_axi_bid(m_axi_bid[2]),
        .s02_axi_bresp(m_axi_bresp[2]),
        .s02_axi_buser(m_axi_buser[2]),
        .s02_axi_bvalid(m_axi_bvalid[2]),
        .s02_axi_bready(m_axi_bready[2]),
        .s02_axi_arid(m_axi_arid[2]),
        .s02_axi_araddr(m_axi_araddr[2]),
        .s02_axi_arlen(m_axi_arlen[2]),
        .s02_axi_arsize(m_axi_arsize[2]),
        .s02_axi_arburst(m_axi_arburst[2]),
        .s02_axi_arlock(m_axi_arlock[2]),
        .s02_axi_arcache(m_axi_arcache[2]),
        .s02_axi_arprot(m_axi_arprot[2]),
        .s02_axi_arqos(m_axi_arqos[2]),
        .s02_axi_aruser(m_axi_aruser[2]),
        .s02_axi_arvalid(m_axi_arvalid[2]),
        .s02_axi_arready(m_axi_arready[2]),
        .s02_axi_rid(m_axi_rid[2]),
        .s02_axi_rdata(m_axi_rdata[2]),
        .s02_axi_rresp(m_axi_rresp[2]),
        .s02_axi_rlast(m_axi_rlast[2]),
        .s02_axi_ruser(m_axi_ruser[2]),
        .s02_axi_rvalid(m_axi_rvalid[2]),
        .s02_axi_rready(m_axi_rready[2]),
        
        .s03_axi_awid(m_axi_awid[3]),
        .s03_axi_awaddr(m_axi_awaddr[3]),
        .s03_axi_awlen(m_axi_awlen[3]),
        .s03_axi_awsize(m_axi_awsize[3]),
        .s03_axi_awburst(m_axi_awburst[3]),
        .s03_axi_awlock(m_axi_awlock[3]),
        .s03_axi_awcache(m_axi_awcache[3]),
        .s03_axi_awprot(m_axi_awprot[3]),
        .s03_axi_awqos(m_axi_awqos[3]),
        .s03_axi_awuser(m_axi_awuser[3]),
        .s03_axi_awvalid(m_axi_awvalid[3]),
        .s03_axi_awready(m_axi_awready[3]),
        .s03_axi_wdata(m_axi_wdata[3]),
        .s03_axi_wstrb(m_axi_wstrb[3]),
        .s03_axi_wlast(m_axi_wlast[3]),
        .s03_axi_wuser(m_axi_wuser[3]),
        .s03_axi_wvalid(m_axi_wvalid[3]),
        .s03_axi_wready(m_axi_wready[3]),
        .s03_axi_bid(m_axi_bid[3]),
        .s03_axi_bresp(m_axi_bresp[3]),
        .s03_axi_buser(m_axi_buser[3]),
        .s03_axi_bvalid(m_axi_bvalid[3]),
        .s03_axi_bready(m_axi_bready[3]),
        .s03_axi_arid(m_axi_arid[3]),
        .s03_axi_araddr(m_axi_araddr[3]),
        .s03_axi_arlen(m_axi_arlen[3]),
        .s03_axi_arsize(m_axi_arsize[3]),
        .s03_axi_arburst(m_axi_arburst[3]),
        .s03_axi_arlock(m_axi_arlock[3]),
        .s03_axi_arcache(m_axi_arcache[3]),
        .s03_axi_arprot(m_axi_arprot[3]),
        .s03_axi_arqos(m_axi_arqos[3]),
        .s03_axi_aruser(m_axi_aruser[3]),
        .s03_axi_arvalid(m_axi_arvalid[3]),
        .s03_axi_arready(m_axi_arready[3]),
        .s03_axi_rid(m_axi_rid[3]),
        .s03_axi_rdata(m_axi_rdata[3]),
        .s03_axi_rresp(m_axi_rresp[3]),
        .s03_axi_rlast(m_axi_rlast[3]),
        .s03_axi_ruser(m_axi_ruser[3]),
        .s03_axi_rvalid(m_axi_rvalid[3]),
        .s03_axi_rready(m_axi_rready[3]),
        
        .s04_axi_awid(m_axi_awid[4]),
        .s04_axi_awaddr(m_axi_awaddr[4]),
        .s04_axi_awlen(m_axi_awlen[4]),
        .s04_axi_awsize(m_axi_awsize[4]),
        .s04_axi_awburst(m_axi_awburst[4]),
        .s04_axi_awlock(m_axi_awlock[4]),
        .s04_axi_awcache(m_axi_awcache[4]),
        .s04_axi_awprot(m_axi_awprot[4]),
        .s04_axi_awqos(m_axi_awqos[4]),
        .s04_axi_awuser(m_axi_awuser[4]),
        .s04_axi_awvalid(m_axi_awvalid[4]),
        .s04_axi_awready(m_axi_awready[4]),
        .s04_axi_wdata(m_axi_wdata[4]),
        .s04_axi_wstrb(m_axi_wstrb[4]),
        .s04_axi_wlast(m_axi_wlast[4]),
        .s04_axi_wuser(m_axi_wuser[4]),
        .s04_axi_wvalid(m_axi_wvalid[4]),
        .s04_axi_wready(m_axi_wready[4]),
        .s04_axi_bid(m_axi_bid[4]),
        .s04_axi_bresp(m_axi_bresp[4]),
        .s04_axi_buser(m_axi_buser[4]),
        .s04_axi_bvalid(m_axi_bvalid[4]),
        .s04_axi_bready(m_axi_bready[4]),
        .s04_axi_arid(m_axi_arid[4]),
        .s04_axi_araddr(m_axi_araddr[4]),
        .s04_axi_arlen(m_axi_arlen[4]),
        .s04_axi_arsize(m_axi_arsize[4]),
        .s04_axi_arburst(m_axi_arburst[4]),
        .s04_axi_arlock(m_axi_arlock[4]),
        .s04_axi_arcache(m_axi_arcache[4]),
        .s04_axi_arprot(m_axi_arprot[4]),
        .s04_axi_arqos(m_axi_arqos[4]),
        .s04_axi_aruser(m_axi_aruser[4]),
        .s04_axi_arvalid(m_axi_arvalid[4]),
        .s04_axi_arready(m_axi_arready[4]),
        .s04_axi_rid(m_axi_rid[4]),
        .s04_axi_rdata(m_axi_rdata[4]),
        .s04_axi_rresp(m_axi_rresp[4]),
        .s04_axi_rlast(m_axi_rlast[4]),
        .s04_axi_ruser(m_axi_ruser[4]),
        .s04_axi_rvalid(m_axi_rvalid[4]),
        .s04_axi_rready(m_axi_rready[4]),

        .s05_axi_awid(m_axi_awid[5]),
        .s05_axi_awaddr(m_axi_awaddr[5]),
        .s05_axi_awlen(m_axi_awlen[5]),
        .s05_axi_awsize(m_axi_awsize[5]),
        .s05_axi_awburst(m_axi_awburst[5]),
        .s05_axi_awlock(m_axi_awlock[5]),
        .s05_axi_awcache(m_axi_awcache[5]),
        .s05_axi_awprot(m_axi_awprot[5]),
        .s05_axi_awqos(m_axi_awqos[5]),
        .s05_axi_awuser(m_axi_awuser[5]),
        .s05_axi_awvalid(m_axi_awvalid[5]),
        .s05_axi_awready(m_axi_awready[5]),
        .s05_axi_wdata(m_axi_wdata[5]),
        .s05_axi_wstrb(m_axi_wstrb[5]),
        .s05_axi_wlast(m_axi_wlast[5]),
        .s05_axi_wuser(m_axi_wuser[5]),
        .s05_axi_wvalid(m_axi_wvalid[5]),
        .s05_axi_wready(m_axi_wready[5]),
        .s05_axi_bid(m_axi_bid[5]),
        .s05_axi_bresp(m_axi_bresp[5]),
        .s05_axi_buser(m_axi_buser[5]),
        .s05_axi_bvalid(m_axi_bvalid[5]),
        .s05_axi_bready(m_axi_bready[5]),
        .s05_axi_arid(m_axi_arid[5]),
        .s05_axi_araddr(m_axi_araddr[5]),
        .s05_axi_arlen(m_axi_arlen[5]),
        .s05_axi_arsize(m_axi_arsize[5]),
        .s05_axi_arburst(m_axi_arburst[5]),
        .s05_axi_arlock(m_axi_arlock[5]),
        .s05_axi_arcache(m_axi_arcache[5]),
        .s05_axi_arprot(m_axi_arprot[5]),
        .s05_axi_arqos(m_axi_arqos[5]),
        .s05_axi_aruser(m_axi_aruser[5]),
        .s05_axi_arvalid(m_axi_arvalid[5]),
        .s05_axi_arready(m_axi_arready[5]),
        .s05_axi_rid(m_axi_rid[5]),
        .s05_axi_rdata(m_axi_rdata[5]),
        .s05_axi_rresp(m_axi_rresp[5]),
        .s05_axi_rlast(m_axi_rlast[5]),
        .s05_axi_ruser(m_axi_ruser[5]),
        .s05_axi_rvalid(m_axi_rvalid[5]),
        .s05_axi_rready(m_axi_rready[5]),

        .s06_axi_awid(m_axi_awid[6]),
        .s06_axi_awaddr(m_axi_awaddr[6]),
        .s06_axi_awlen(m_axi_awlen[6]),
        .s06_axi_awsize(m_axi_awsize[6]),
        .s06_axi_awburst(m_axi_awburst[6]),
        .s06_axi_awlock(m_axi_awlock[6]),
        .s06_axi_awcache(m_axi_awcache[6]),
        .s06_axi_awprot(m_axi_awprot[6]),
        .s06_axi_awqos(m_axi_awqos[6]),
        .s06_axi_awuser(m_axi_awuser[6]),
        .s06_axi_awvalid(m_axi_awvalid[6]),
        .s06_axi_awready(m_axi_awready[6]),
        .s06_axi_wdata(m_axi_wdata[6]),
        .s06_axi_wstrb(m_axi_wstrb[6]),
        .s06_axi_wlast(m_axi_wlast[6]),
        .s06_axi_wuser(m_axi_wuser[6]),
        .s06_axi_wvalid(m_axi_wvalid[6]),
        .s06_axi_wready(m_axi_wready[6]),
        .s06_axi_bid(m_axi_bid[6]),
        .s06_axi_bresp(m_axi_bresp[6]),
        .s06_axi_buser(m_axi_buser[6]),
        .s06_axi_bvalid(m_axi_bvalid[6]),
        .s06_axi_bready(m_axi_bready[6]),
        .s06_axi_arid(m_axi_arid[6]),
        .s06_axi_araddr(m_axi_araddr[6]),
        .s06_axi_arlen(m_axi_arlen[6]),
        .s06_axi_arsize(m_axi_arsize[6]),
        .s06_axi_arburst(m_axi_arburst[6]),
        .s06_axi_arlock(m_axi_arlock[6]),
        .s06_axi_arcache(m_axi_arcache[6]),
        .s06_axi_arprot(m_axi_arprot[6]),
        .s06_axi_arqos(m_axi_arqos[6]),
        .s06_axi_aruser(m_axi_aruser[6]),
        .s06_axi_arvalid(m_axi_arvalid[6]),
        .s06_axi_arready(m_axi_arready[6]),
        .s06_axi_rid(m_axi_rid[6]),
        .s06_axi_rdata(m_axi_rdata[6]),
        .s06_axi_rresp(m_axi_rresp[6]),
        .s06_axi_rlast(m_axi_rlast[6]),
        .s06_axi_ruser(m_axi_ruser[6]),
        .s06_axi_rvalid(m_axi_rvalid[6]),
        .s06_axi_rready(m_axi_rready[6]),        
        
        .s07_axi_awid(m_axi_awid[7]),
        .s07_axi_awaddr(m_axi_awaddr[7]),
        .s07_axi_awlen(m_axi_awlen[7]),
        .s07_axi_awsize(m_axi_awsize[7]),
        .s07_axi_awburst(m_axi_awburst[7]),
        .s07_axi_awlock(m_axi_awlock[7]),
        .s07_axi_awcache(m_axi_awcache[7]),
        .s07_axi_awprot(m_axi_awprot[7]),
        .s07_axi_awqos(m_axi_awqos[7]),
        .s07_axi_awuser(m_axi_awuser[7]),
        .s07_axi_awvalid(m_axi_awvalid[7]),
        .s07_axi_awready(m_axi_awready[7]),
        .s07_axi_wdata(m_axi_wdata[7]),
        .s07_axi_wstrb(m_axi_wstrb[7]),
        .s07_axi_wlast(m_axi_wlast[7]),
        .s07_axi_wuser(m_axi_wuser[7]),
        .s07_axi_wvalid(m_axi_wvalid[7]),
        .s07_axi_wready(m_axi_wready[7]),
        .s07_axi_bid(m_axi_bid[7]),
        .s07_axi_bresp(m_axi_bresp[7]),
        .s07_axi_buser(m_axi_buser[7]),
        .s07_axi_bvalid(m_axi_bvalid[7]),
        .s07_axi_bready(m_axi_bready[7]),
        .s07_axi_arid(m_axi_arid[7]),
        .s07_axi_araddr(m_axi_araddr[7]),
        .s07_axi_arlen(m_axi_arlen[7]),
        .s07_axi_arsize(m_axi_arsize[7]),
        .s07_axi_arburst(m_axi_arburst[7]),
        .s07_axi_arlock(m_axi_arlock[7]),
        .s07_axi_arcache(m_axi_arcache[7]),
        .s07_axi_arprot(m_axi_arprot[7]),
        .s07_axi_arqos(m_axi_arqos[7]),
        .s07_axi_aruser(m_axi_aruser[7]),
        .s07_axi_arvalid(m_axi_arvalid[7]),
        .s07_axi_arready(m_axi_arready[7]),
        .s07_axi_rid(m_axi_rid[7]),
        .s07_axi_rdata(m_axi_rdata[7]),
        .s07_axi_rresp(m_axi_rresp[7]),
        .s07_axi_rlast(m_axi_rlast[7]),
        .s07_axi_ruser(m_axi_ruser[7]),
        .s07_axi_rvalid(m_axi_rvalid[7]),
        .s07_axi_rready(m_axi_rready[7]),
        
        .s08_axi_awid(m_axi_awid[8]),
        .s08_axi_awaddr(m_axi_awaddr[8]),
        .s08_axi_awlen(m_axi_awlen[8]),
        .s08_axi_awsize(m_axi_awsize[8]),
        .s08_axi_awburst(m_axi_awburst[8]),
        .s08_axi_awlock(m_axi_awlock[8]),
        .s08_axi_awcache(m_axi_awcache[8]),
        .s08_axi_awprot(m_axi_awprot[8]),
        .s08_axi_awqos(m_axi_awqos[8]),
        .s08_axi_awuser(m_axi_awuser[8]),
        .s08_axi_awvalid(m_axi_awvalid[8]),
        .s08_axi_awready(m_axi_awready[8]),
        .s08_axi_wdata(m_axi_wdata[8]),
        .s08_axi_wstrb(m_axi_wstrb[8]),
        .s08_axi_wlast(m_axi_wlast[8]),
        .s08_axi_wuser(m_axi_wuser[8]),
        .s08_axi_wvalid(m_axi_wvalid[8]),
        .s08_axi_wready(m_axi_wready[8]),
        .s08_axi_bid(m_axi_bid[8]),
        .s08_axi_bresp(m_axi_bresp[8]),
        .s08_axi_buser(m_axi_buser[8]),
        .s08_axi_bvalid(m_axi_bvalid[8]),
        .s08_axi_bready(m_axi_bready[8]),
        .s08_axi_arid(m_axi_arid[8]),
        .s08_axi_araddr(m_axi_araddr[8]),
        .s08_axi_arlen(m_axi_arlen[8]),
        .s08_axi_arsize(m_axi_arsize[8]),
        .s08_axi_arburst(m_axi_arburst[8]),
        .s08_axi_arlock(m_axi_arlock[8]),
        .s08_axi_arcache(m_axi_arcache[8]),
        .s08_axi_arprot(m_axi_arprot[8]),
        .s08_axi_arqos(m_axi_arqos[8]),
        .s08_axi_aruser(m_axi_aruser[8]),
        .s08_axi_arvalid(m_axi_arvalid[8]),
        .s08_axi_arready(m_axi_arready[8]),
        .s08_axi_rid(m_axi_rid[8]),
        .s08_axi_rdata(m_axi_rdata[8]),
        .s08_axi_rresp(m_axi_rresp[8]),
        .s08_axi_rlast(m_axi_rlast[8]),
        .s08_axi_ruser(m_axi_ruser[8]),
        .s08_axi_rvalid(m_axi_rvalid[8]),
        .s08_axi_rready(m_axi_rready[8]),
        
        .s09_axi_awid(m_axi_awid[9]),
        .s09_axi_awaddr(m_axi_awaddr[9]),
        .s09_axi_awlen(m_axi_awlen[9]),
        .s09_axi_awsize(m_axi_awsize[9]),
        .s09_axi_awburst(m_axi_awburst[9]),
        .s09_axi_awlock(m_axi_awlock[9]),
        .s09_axi_awcache(m_axi_awcache[9]),
        .s09_axi_awprot(m_axi_awprot[9]),
        .s09_axi_awqos(m_axi_awqos[9]),
        .s09_axi_awuser(m_axi_awuser[9]),
        .s09_axi_awvalid(m_axi_awvalid[9]),
        .s09_axi_awready(m_axi_awready[9]),
        .s09_axi_wdata(m_axi_wdata[9]),
        .s09_axi_wstrb(m_axi_wstrb[9]),
        .s09_axi_wlast(m_axi_wlast[9]),
        .s09_axi_wuser(m_axi_wuser[9]),
        .s09_axi_wvalid(m_axi_wvalid[9]),
        .s09_axi_wready(m_axi_wready[9]),
        .s09_axi_bid(m_axi_bid[9]),
        .s09_axi_bresp(m_axi_bresp[9]),
        .s09_axi_buser(m_axi_buser[9]),
        .s09_axi_bvalid(m_axi_bvalid[9]),
        .s09_axi_bready(m_axi_bready[9]),
        .s09_axi_arid(m_axi_arid[9]),
        .s09_axi_araddr(m_axi_araddr[9]),
        .s09_axi_arlen(m_axi_arlen[9]),
        .s09_axi_arsize(m_axi_arsize[9]),
        .s09_axi_arburst(m_axi_arburst[9]),
        .s09_axi_arlock(m_axi_arlock[9]),
        .s09_axi_arcache(m_axi_arcache[9]),
        .s09_axi_arprot(m_axi_arprot[9]),
        .s09_axi_arqos(m_axi_arqos[9]),
        .s09_axi_aruser(m_axi_aruser[9]),
        .s09_axi_arvalid(m_axi_arvalid[9]),
        .s09_axi_arready(m_axi_arready[9]),
        .s09_axi_rid(m_axi_rid[9]),
        .s09_axi_rdata(m_axi_rdata[9]),
        .s09_axi_rresp(m_axi_rresp[9]),
        .s09_axi_rlast(m_axi_rlast[9]),
        .s09_axi_ruser(m_axi_ruser[9]),
        .s09_axi_rvalid(m_axi_rvalid[9]),
        .s09_axi_rready(m_axi_rready[9]),

        .s10_axi_awid(m_axi_awid[10]),
        .s10_axi_awaddr(m_axi_awaddr[10]),
        .s10_axi_awlen(m_axi_awlen[10]),
        .s10_axi_awsize(m_axi_awsize[10]),
        .s10_axi_awburst(m_axi_awburst[10]),
        .s10_axi_awlock(m_axi_awlock[10]),
        .s10_axi_awcache(m_axi_awcache[10]),
        .s10_axi_awprot(m_axi_awprot[10]),
        .s10_axi_awqos(m_axi_awqos[10]),
        .s10_axi_awuser(m_axi_awuser[10]),
        .s10_axi_awvalid(m_axi_awvalid[10]),
        .s10_axi_awready(m_axi_awready[10]),
        .s10_axi_wdata(m_axi_wdata[10]),
        .s10_axi_wstrb(m_axi_wstrb[10]),
        .s10_axi_wlast(m_axi_wlast[10]),
        .s10_axi_wuser(m_axi_wuser[10]),
        .s10_axi_wvalid(m_axi_wvalid[10]),
        .s10_axi_wready(m_axi_wready[10]),
        .s10_axi_bid(m_axi_bid[10]),
        .s10_axi_bresp(m_axi_bresp[10]),
        .s10_axi_buser(m_axi_buser[10]),
        .s10_axi_bvalid(m_axi_bvalid[10]),
        .s10_axi_bready(m_axi_bready[10]),
        .s10_axi_arid(m_axi_arid[10]),
        .s10_axi_araddr(m_axi_araddr[10]),
        .s10_axi_arlen(m_axi_arlen[10]),
        .s10_axi_arsize(m_axi_arsize[10]),
        .s10_axi_arburst(m_axi_arburst[10]),
        .s10_axi_arlock(m_axi_arlock[10]),
        .s10_axi_arcache(m_axi_arcache[10]),
        .s10_axi_arprot(m_axi_arprot[10]),
        .s10_axi_arqos(m_axi_arqos[10]),
        .s10_axi_aruser(m_axi_aruser[10]),
        .s10_axi_arvalid(m_axi_arvalid[10]),
        .s10_axi_arready(m_axi_arready[10]),
        .s10_axi_rid(m_axi_rid[10]),
        .s10_axi_rdata(m_axi_rdata[10]),
        .s10_axi_rresp(m_axi_rresp[10]),
        .s10_axi_rlast(m_axi_rlast[10]),
        .s10_axi_ruser(m_axi_ruser[10]),
        .s10_axi_rvalid(m_axi_rvalid[10]),
        .s10_axi_rready(m_axi_rready[10]),
        
        .s11_axi_awid(m_axi_awid[11]),
        .s11_axi_awaddr(m_axi_awaddr[11]),
        .s11_axi_awlen(m_axi_awlen[11]),
        .s11_axi_awsize(m_axi_awsize[11]),
        .s11_axi_awburst(m_axi_awburst[11]),
        .s11_axi_awlock(m_axi_awlock[11]),
        .s11_axi_awcache(m_axi_awcache[11]),
        .s11_axi_awprot(m_axi_awprot[11]),
        .s11_axi_awqos(m_axi_awqos[11]),
        .s11_axi_awuser(m_axi_awuser[11]),
        .s11_axi_awvalid(m_axi_awvalid[11]),
        .s11_axi_awready(m_axi_awready[11]),
        .s11_axi_wdata(m_axi_wdata[11]),
        .s11_axi_wstrb(m_axi_wstrb[11]),
        .s11_axi_wlast(m_axi_wlast[11]),
        .s11_axi_wuser(m_axi_wuser[11]),
        .s11_axi_wvalid(m_axi_wvalid[11]),
        .s11_axi_wready(m_axi_wready[11]),
        .s11_axi_bid(m_axi_bid[11]),
        .s11_axi_bresp(m_axi_bresp[11]),
        .s11_axi_buser(m_axi_buser[11]),
        .s11_axi_bvalid(m_axi_bvalid[11]),
        .s11_axi_bready(m_axi_bready[11]),
        .s11_axi_arid(m_axi_arid[11]),
        .s11_axi_araddr(m_axi_araddr[11]),
        .s11_axi_arlen(m_axi_arlen[11]),
        .s11_axi_arsize(m_axi_arsize[11]),
        .s11_axi_arburst(m_axi_arburst[11]),
        .s11_axi_arlock(m_axi_arlock[11]),
        .s11_axi_arcache(m_axi_arcache[11]),
        .s11_axi_arprot(m_axi_arprot[11]),
        .s11_axi_arqos(m_axi_arqos[11]),
        .s11_axi_aruser(m_axi_aruser[11]),
        .s11_axi_arvalid(m_axi_arvalid[11]),
        .s11_axi_arready(m_axi_arready[11]),
        .s11_axi_rid(m_axi_rid[11]),
        .s11_axi_rdata(m_axi_rdata[11]),
        .s11_axi_rresp(m_axi_rresp[11]),
        .s11_axi_rlast(m_axi_rlast[11]),
        .s11_axi_ruser(m_axi_ruser[11]),
        .s11_axi_rvalid(m_axi_rvalid[11]),
        .s11_axi_rready(m_axi_rready[11]),
        
        .s12_axi_awid(m_axi_awid[12]),
        .s12_axi_awaddr(m_axi_awaddr[12]),
        .s12_axi_awlen(m_axi_awlen[12]),
        .s12_axi_awsize(m_axi_awsize[12]),
        .s12_axi_awburst(m_axi_awburst[12]),
        .s12_axi_awlock(m_axi_awlock[12]),
        .s12_axi_awcache(m_axi_awcache[12]),
        .s12_axi_awprot(m_axi_awprot[12]),
        .s12_axi_awqos(m_axi_awqos[12]),
        .s12_axi_awuser(m_axi_awuser[12]),
        .s12_axi_awvalid(m_axi_awvalid[12]),
        .s12_axi_awready(m_axi_awready[12]),
        .s12_axi_wdata(m_axi_wdata[12]),
        .s12_axi_wstrb(m_axi_wstrb[12]),
        .s12_axi_wlast(m_axi_wlast[12]),
        .s12_axi_wuser(m_axi_wuser[12]),
        .s12_axi_wvalid(m_axi_wvalid[12]),
        .s12_axi_wready(m_axi_wready[12]),
        .s12_axi_bid(m_axi_bid[12]),
        .s12_axi_bresp(m_axi_bresp[12]),
        .s12_axi_buser(m_axi_buser[12]),
        .s12_axi_bvalid(m_axi_bvalid[12]),
        .s12_axi_bready(m_axi_bready[12]),
        .s12_axi_arid(m_axi_arid[12]),
        .s12_axi_araddr(m_axi_araddr[12]),
        .s12_axi_arlen(m_axi_arlen[12]),
        .s12_axi_arsize(m_axi_arsize[12]),
        .s12_axi_arburst(m_axi_arburst[12]),
        .s12_axi_arlock(m_axi_arlock[12]),
        .s12_axi_arcache(m_axi_arcache[12]),
        .s12_axi_arprot(m_axi_arprot[12]),
        .s12_axi_arqos(m_axi_arqos[12]),
        .s12_axi_aruser(m_axi_aruser[12]),
        .s12_axi_arvalid(m_axi_arvalid[12]),
        .s12_axi_arready(m_axi_arready[12]),
        .s12_axi_rid(m_axi_rid[12]),
        .s12_axi_rdata(m_axi_rdata[12]),
        .s12_axi_rresp(m_axi_rresp[12]),
        .s12_axi_rlast(m_axi_rlast[12]),
        .s12_axi_ruser(m_axi_ruser[12]),
        .s12_axi_rvalid(m_axi_rvalid[12]),
        .s12_axi_rready(m_axi_rready[12]),                                                
        
        .s13_axi_awid(m_axi_awid[13]),
        .s13_axi_awaddr(m_axi_awaddr[13]),
        .s13_axi_awlen(m_axi_awlen[13]),
        .s13_axi_awsize(m_axi_awsize[13]),
        .s13_axi_awburst(m_axi_awburst[13]),
        .s13_axi_awlock(m_axi_awlock[13]),
        .s13_axi_awcache(m_axi_awcache[13]),
        .s13_axi_awprot(m_axi_awprot[13]),
        .s13_axi_awqos(m_axi_awqos[13]),
        .s13_axi_awuser(m_axi_awuser[13]),
        .s13_axi_awvalid(m_axi_awvalid[13]),
        .s13_axi_awready(m_axi_awready[13]),
        .s13_axi_wdata(m_axi_wdata[13]),
        .s13_axi_wstrb(m_axi_wstrb[13]),
        .s13_axi_wlast(m_axi_wlast[13]),
        .s13_axi_wuser(m_axi_wuser[13]),
        .s13_axi_wvalid(m_axi_wvalid[13]),
        .s13_axi_wready(m_axi_wready[13]),
        .s13_axi_bid(m_axi_bid[13]),
        .s13_axi_bresp(m_axi_bresp[13]),
        .s13_axi_buser(m_axi_buser[13]),
        .s13_axi_bvalid(m_axi_bvalid[13]),
        .s13_axi_bready(m_axi_bready[13]),
        .s13_axi_arid(m_axi_arid[13]),
        .s13_axi_araddr(m_axi_araddr[13]),
        .s13_axi_arlen(m_axi_arlen[13]),
        .s13_axi_arsize(m_axi_arsize[13]),
        .s13_axi_arburst(m_axi_arburst[13]),
        .s13_axi_arlock(m_axi_arlock[13]),
        .s13_axi_arcache(m_axi_arcache[13]),
        .s13_axi_arprot(m_axi_arprot[13]),
        .s13_axi_arqos(m_axi_arqos[13]),
        .s13_axi_aruser(m_axi_aruser[13]),
        .s13_axi_arvalid(m_axi_arvalid[13]),
        .s13_axi_arready(m_axi_arready[13]),
        .s13_axi_rid(m_axi_rid[13]),
        .s13_axi_rdata(m_axi_rdata[13]),
        .s13_axi_rresp(m_axi_rresp[13]),
        .s13_axi_rlast(m_axi_rlast[13]),
        .s13_axi_ruser(m_axi_ruser[13]),
        .s13_axi_rvalid(m_axi_rvalid[13]),
        .s13_axi_rready(m_axi_rready[13]),
        
        .s14_axi_awid(m_axi_awid[14]),
        .s14_axi_awaddr(m_axi_awaddr[14]),
        .s14_axi_awlen(m_axi_awlen[14]),
        .s14_axi_awsize(m_axi_awsize[14]),
        .s14_axi_awburst(m_axi_awburst[14]),
        .s14_axi_awlock(m_axi_awlock[14]),
        .s14_axi_awcache(m_axi_awcache[14]),
        .s14_axi_awprot(m_axi_awprot[14]),
        .s14_axi_awqos(m_axi_awqos[14]),
        .s14_axi_awuser(m_axi_awuser[14]),
        .s14_axi_awvalid(m_axi_awvalid[14]),
        .s14_axi_awready(m_axi_awready[14]),
        .s14_axi_wdata(m_axi_wdata[14]),
        .s14_axi_wstrb(m_axi_wstrb[14]),
        .s14_axi_wlast(m_axi_wlast[14]),
        .s14_axi_wuser(m_axi_wuser[14]),
        .s14_axi_wvalid(m_axi_wvalid[14]),
        .s14_axi_wready(m_axi_wready[14]),
        .s14_axi_bid(m_axi_bid[14]),
        .s14_axi_bresp(m_axi_bresp[14]),
        .s14_axi_buser(m_axi_buser[14]),
        .s14_axi_bvalid(m_axi_bvalid[14]),
        .s14_axi_bready(m_axi_bready[14]),
        .s14_axi_arid(m_axi_arid[14]),
        .s14_axi_araddr(m_axi_araddr[14]),
        .s14_axi_arlen(m_axi_arlen[14]),
        .s14_axi_arsize(m_axi_arsize[14]),
        .s14_axi_arburst(m_axi_arburst[14]),
        .s14_axi_arlock(m_axi_arlock[14]),
        .s14_axi_arcache(m_axi_arcache[14]),
        .s14_axi_arprot(m_axi_arprot[14]),
        .s14_axi_arqos(m_axi_arqos[14]),
        .s14_axi_aruser(m_axi_aruser[14]),
        .s14_axi_arvalid(m_axi_arvalid[14]),
        .s14_axi_arready(m_axi_arready[14]),
        .s14_axi_rid(m_axi_rid[14]),
        .s14_axi_rdata(m_axi_rdata[14]),
        .s14_axi_rresp(m_axi_rresp[14]),
        .s14_axi_rlast(m_axi_rlast[14]),
        .s14_axi_ruser(m_axi_ruser[14]),
        .s14_axi_rvalid(m_axi_rvalid[14]),
        .s14_axi_rready(m_axi_rready[14]),
        
        .s15_axi_awid(m_axi_awid[15]),
        .s15_axi_awaddr(m_axi_awaddr[15]),
        .s15_axi_awlen(m_axi_awlen[15]),
        .s15_axi_awsize(m_axi_awsize[15]),
        .s15_axi_awburst(m_axi_awburst[15]),
        .s15_axi_awlock(m_axi_awlock[15]),
        .s15_axi_awcache(m_axi_awcache[15]),
        .s15_axi_awprot(m_axi_awprot[15]),
        .s15_axi_awqos(m_axi_awqos[15]),
        .s15_axi_awuser(m_axi_awuser[15]),
        .s15_axi_awvalid(m_axi_awvalid[15]),
        .s15_axi_awready(m_axi_awready[15]),
        .s15_axi_wdata(m_axi_wdata[15]),
        .s15_axi_wstrb(m_axi_wstrb[15]),
        .s15_axi_wlast(m_axi_wlast[15]),
        .s15_axi_wuser(m_axi_wuser[15]),
        .s15_axi_wvalid(m_axi_wvalid[15]),
        .s15_axi_wready(m_axi_wready[15]),
        .s15_axi_bid(m_axi_bid[15]),
        .s15_axi_bresp(m_axi_bresp[15]),
        .s15_axi_buser(m_axi_buser[15]),
        .s15_axi_bvalid(m_axi_bvalid[15]),
        .s15_axi_bready(m_axi_bready[15]),
        .s15_axi_arid(m_axi_arid[15]),
        .s15_axi_araddr(m_axi_araddr[15]),
        .s15_axi_arlen(m_axi_arlen[15]),
        .s15_axi_arsize(m_axi_arsize[15]),
        .s15_axi_arburst(m_axi_arburst[15]),
        .s15_axi_arlock(m_axi_arlock[15]),
        .s15_axi_arcache(m_axi_arcache[15]),
        .s15_axi_arprot(m_axi_arprot[15]),
        .s15_axi_arqos(m_axi_arqos[15]),
        .s15_axi_aruser(m_axi_aruser[15]),
        .s15_axi_arvalid(m_axi_arvalid[15]),
        .s15_axi_arready(m_axi_arready[15]),
        .s15_axi_rid(m_axi_rid[15]),
        .s15_axi_rdata(m_axi_rdata[15]),
        .s15_axi_rresp(m_axi_rresp[15]),
        .s15_axi_rlast(m_axi_rlast[15]),
        .s15_axi_ruser(m_axi_ruser[15]),
        .s15_axi_rvalid(m_axi_rvalid[15]),
        .s15_axi_rready(m_axi_rready[15]),
        
        .s16_axi_awid(m_axi_awid[16]),
        .s16_axi_awaddr(m_axi_awaddr[16]),
        .s16_axi_awlen(m_axi_awlen[16]),
        .s16_axi_awsize(m_axi_awsize[16]),
        .s16_axi_awburst(m_axi_awburst[16]),
        .s16_axi_awlock(m_axi_awlock[16]),
        .s16_axi_awcache(m_axi_awcache[16]),
        .s16_axi_awprot(m_axi_awprot[16]),
        .s16_axi_awqos(m_axi_awqos[16]),
        .s16_axi_awuser(m_axi_awuser[16]),
        .s16_axi_awvalid(m_axi_awvalid[16]),
        .s16_axi_awready(m_axi_awready[16]),
        .s16_axi_wdata(m_axi_wdata[16]),
        .s16_axi_wstrb(m_axi_wstrb[16]),
        .s16_axi_wlast(m_axi_wlast[16]),
        .s16_axi_wuser(m_axi_wuser[16]),
        .s16_axi_wvalid(m_axi_wvalid[16]),
        .s16_axi_wready(m_axi_wready[16]),
        .s16_axi_bid(m_axi_bid[16]),
        .s16_axi_bresp(m_axi_bresp[16]),
        .s16_axi_buser(m_axi_buser[16]),
        .s16_axi_bvalid(m_axi_bvalid[16]),
        .s16_axi_bready(m_axi_bready[16]),
        .s16_axi_arid(m_axi_arid[16]),
        .s16_axi_araddr(m_axi_araddr[16]),
        .s16_axi_arlen(m_axi_arlen[16]),
        .s16_axi_arsize(m_axi_arsize[16]),
        .s16_axi_arburst(m_axi_arburst[16]),
        .s16_axi_arlock(m_axi_arlock[16]),
        .s16_axi_arcache(m_axi_arcache[16]),
        .s16_axi_arprot(m_axi_arprot[16]),
        .s16_axi_arqos(m_axi_arqos[16]),
        .s16_axi_aruser(m_axi_aruser[16]),
        .s16_axi_arvalid(m_axi_arvalid[16]),
        .s16_axi_arready(m_axi_arready[16]),
        .s16_axi_rid(m_axi_rid[16]),
        .s16_axi_rdata(m_axi_rdata[16]),
        .s16_axi_rresp(m_axi_rresp[16]),
        .s16_axi_rlast(m_axi_rlast[16]),
        .s16_axi_ruser(m_axi_ruser[16]),
        .s16_axi_rvalid(m_axi_rvalid[16]),
        .s16_axi_rready(m_axi_rready[16]),
        
        .s17_axi_awid(m_axi_awid[17]),
        .s17_axi_awaddr(m_axi_awaddr[17]),
        .s17_axi_awlen(m_axi_awlen[17]),
        .s17_axi_awsize(m_axi_awsize[17]),
        .s17_axi_awburst(m_axi_awburst[17]),
        .s17_axi_awlock(m_axi_awlock[17]),
        .s17_axi_awcache(m_axi_awcache[17]),
        .s17_axi_awprot(m_axi_awprot[17]),
        .s17_axi_awqos(m_axi_awqos[17]),
        .s17_axi_awuser(m_axi_awuser[17]),
        .s17_axi_awvalid(m_axi_awvalid[17]),
        .s17_axi_awready(m_axi_awready[17]),
        .s17_axi_wdata(m_axi_wdata[17]),
        .s17_axi_wstrb(m_axi_wstrb[17]),
        .s17_axi_wlast(m_axi_wlast[17]),
        .s17_axi_wuser(m_axi_wuser[17]),
        .s17_axi_wvalid(m_axi_wvalid[17]),
        .s17_axi_wready(m_axi_wready[17]),
        .s17_axi_bid(m_axi_bid[17]),
        .s17_axi_bresp(m_axi_bresp[17]),
        .s17_axi_buser(m_axi_buser[17]),
        .s17_axi_bvalid(m_axi_bvalid[17]),
        .s17_axi_bready(m_axi_bready[17]),
        .s17_axi_arid(m_axi_arid[17]),
        .s17_axi_araddr(m_axi_araddr[17]),
        .s17_axi_arlen(m_axi_arlen[17]),
        .s17_axi_arsize(m_axi_arsize[17]),
        .s17_axi_arburst(m_axi_arburst[17]),
        .s17_axi_arlock(m_axi_arlock[17]),
        .s17_axi_arcache(m_axi_arcache[17]),
        .s17_axi_arprot(m_axi_arprot[17]),
        .s17_axi_arqos(m_axi_arqos[17]),
        .s17_axi_aruser(m_axi_aruser[17]),
        .s17_axi_arvalid(m_axi_arvalid[17]),
        .s17_axi_arready(m_axi_arready[17]),
        .s17_axi_rid(m_axi_rid[17]),
        .s17_axi_rdata(m_axi_rdata[17]),
        .s17_axi_rresp(m_axi_rresp[17]),
        .s17_axi_rlast(m_axi_rlast[17]),
        .s17_axi_ruser(m_axi_ruser[17]),
        .s17_axi_rvalid(m_axi_rvalid[17]),
        .s17_axi_rready(m_axi_rready[17]),
        
        .s18_axi_awid(m_axi_awid[18]),
        .s18_axi_awaddr(m_axi_awaddr[18]),
        .s18_axi_awlen(m_axi_awlen[18]),
        .s18_axi_awsize(m_axi_awsize[18]),
        .s18_axi_awburst(m_axi_awburst[18]),
        .s18_axi_awlock(m_axi_awlock[18]),
        .s18_axi_awcache(m_axi_awcache[18]),
        .s18_axi_awprot(m_axi_awprot[18]),
        .s18_axi_awqos(m_axi_awqos[18]),
        .s18_axi_awuser(m_axi_awuser[18]),
        .s18_axi_awvalid(m_axi_awvalid[18]),
        .s18_axi_awready(m_axi_awready[18]),
        .s18_axi_wdata(m_axi_wdata[18]),
        .s18_axi_wstrb(m_axi_wstrb[18]),
        .s18_axi_wlast(m_axi_wlast[18]),
        .s18_axi_wuser(m_axi_wuser[18]),
        .s18_axi_wvalid(m_axi_wvalid[18]),
        .s18_axi_wready(m_axi_wready[18]),
        .s18_axi_bid(m_axi_bid[18]),
        .s18_axi_bresp(m_axi_bresp[18]),
        .s18_axi_buser(m_axi_buser[18]),
        .s18_axi_bvalid(m_axi_bvalid[18]),
        .s18_axi_bready(m_axi_bready[18]),
        .s18_axi_arid(m_axi_arid[18]),
        .s18_axi_araddr(m_axi_araddr[18]),
        .s18_axi_arlen(m_axi_arlen[18]),
        .s18_axi_arsize(m_axi_arsize[18]),
        .s18_axi_arburst(m_axi_arburst[18]),
        .s18_axi_arlock(m_axi_arlock[18]),
        .s18_axi_arcache(m_axi_arcache[18]),
        .s18_axi_arprot(m_axi_arprot[18]),
        .s18_axi_arqos(m_axi_arqos[18]),
        .s18_axi_aruser(m_axi_aruser[18]),
        .s18_axi_arvalid(m_axi_arvalid[18]),
        .s18_axi_arready(m_axi_arready[18]),
        .s18_axi_rid(m_axi_rid[18]),
        .s18_axi_rdata(m_axi_rdata[18]),
        .s18_axi_rresp(m_axi_rresp[18]),
        .s18_axi_rlast(m_axi_rlast[18]),
        .s18_axi_ruser(m_axi_ruser[18]),
        .s18_axi_rvalid(m_axi_rvalid[18]),
        .s18_axi_rready(m_axi_rready[18]),
        
        .s19_axi_awid(m_axi_awid[19]),
        .s19_axi_awaddr(m_axi_awaddr[19]),
        .s19_axi_awlen(m_axi_awlen[19]),
        .s19_axi_awsize(m_axi_awsize[19]),
        .s19_axi_awburst(m_axi_awburst[19]),
        .s19_axi_awlock(m_axi_awlock[19]),
        .s19_axi_awcache(m_axi_awcache[19]),
        .s19_axi_awprot(m_axi_awprot[19]),
        .s19_axi_awqos(m_axi_awqos[19]),
        .s19_axi_awuser(m_axi_awuser[19]),
        .s19_axi_awvalid(m_axi_awvalid[19]),
        .s19_axi_awready(m_axi_awready[19]),
        .s19_axi_wdata(m_axi_wdata[19]),
        .s19_axi_wstrb(m_axi_wstrb[19]),
        .s19_axi_wlast(m_axi_wlast[19]),
        .s19_axi_wuser(m_axi_wuser[19]),
        .s19_axi_wvalid(m_axi_wvalid[19]),
        .s19_axi_wready(m_axi_wready[19]),
        .s19_axi_bid(m_axi_bid[19]),
        .s19_axi_bresp(m_axi_bresp[19]),
        .s19_axi_buser(m_axi_buser[19]),
        .s19_axi_bvalid(m_axi_bvalid[19]),
        .s19_axi_bready(m_axi_bready[19]),
        .s19_axi_arid(m_axi_arid[19]),
        .s19_axi_araddr(m_axi_araddr[19]),
        .s19_axi_arlen(m_axi_arlen[19]),
        .s19_axi_arsize(m_axi_arsize[19]),
        .s19_axi_arburst(m_axi_arburst[19]),
        .s19_axi_arlock(m_axi_arlock[19]),
        .s19_axi_arcache(m_axi_arcache[19]),
        .s19_axi_arprot(m_axi_arprot[19]),
        .s19_axi_arqos(m_axi_arqos[19]),
        .s19_axi_aruser(m_axi_aruser[19]),
        .s19_axi_arvalid(m_axi_arvalid[19]),
        .s19_axi_arready(m_axi_arready[19]),
        .s19_axi_rid(m_axi_rid[19]),
        .s19_axi_rdata(m_axi_rdata[19]),
        .s19_axi_rresp(m_axi_rresp[19]),
        .s19_axi_rlast(m_axi_rlast[19]),
        .s19_axi_ruser(m_axi_ruser[19]),
        .s19_axi_rvalid(m_axi_rvalid[19]),
        .s19_axi_rready(m_axi_rready[19]),
        
        .s20_axi_awid(m_axi_awid[20]),
        .s20_axi_awaddr(m_axi_awaddr[20]),
        .s20_axi_awlen(m_axi_awlen[20]),
        .s20_axi_awsize(m_axi_awsize[20]),
        .s20_axi_awburst(m_axi_awburst[20]),
        .s20_axi_awlock(m_axi_awlock[20]),
        .s20_axi_awcache(m_axi_awcache[20]),
        .s20_axi_awprot(m_axi_awprot[20]),
        .s20_axi_awqos(m_axi_awqos[20]),
        .s20_axi_awuser(m_axi_awuser[20]),
        .s20_axi_awvalid(m_axi_awvalid[20]),
        .s20_axi_awready(m_axi_awready[20]),
        .s20_axi_wdata(m_axi_wdata[20]),
        .s20_axi_wstrb(m_axi_wstrb[20]),
        .s20_axi_wlast(m_axi_wlast[20]),
        .s20_axi_wuser(m_axi_wuser[20]),
        .s20_axi_wvalid(m_axi_wvalid[20]),
        .s20_axi_wready(m_axi_wready[20]),
        .s20_axi_bid(m_axi_bid[20]),
        .s20_axi_bresp(m_axi_bresp[20]),
        .s20_axi_buser(m_axi_buser[20]),
        .s20_axi_bvalid(m_axi_bvalid[20]),
        .s20_axi_bready(m_axi_bready[20]),
        .s20_axi_arid(m_axi_arid[20]),
        .s20_axi_araddr(m_axi_araddr[20]),
        .s20_axi_arlen(m_axi_arlen[20]),
        .s20_axi_arsize(m_axi_arsize[20]),
        .s20_axi_arburst(m_axi_arburst[20]),
        .s20_axi_arlock(m_axi_arlock[20]),
        .s20_axi_arcache(m_axi_arcache[20]),
        .s20_axi_arprot(m_axi_arprot[20]),
        .s20_axi_arqos(m_axi_arqos[20]),
        .s20_axi_aruser(m_axi_aruser[20]),
        .s20_axi_arvalid(m_axi_arvalid[20]),
        .s20_axi_arready(m_axi_arready[20]),
        .s20_axi_rid(m_axi_rid[20]),
        .s20_axi_rdata(m_axi_rdata[20]),
        .s20_axi_rresp(m_axi_rresp[20]),
        .s20_axi_rlast(m_axi_rlast[20]),
        .s20_axi_ruser(m_axi_ruser[20]),
        .s20_axi_rvalid(m_axi_rvalid[20]),
        .s20_axi_rready(m_axi_rready[20]),
        
        .s21_axi_awid(m_axi_awid[21]),
        .s21_axi_awaddr(m_axi_awaddr[21]),
        .s21_axi_awlen(m_axi_awlen[21]),
        .s21_axi_awsize(m_axi_awsize[21]),
        .s21_axi_awburst(m_axi_awburst[21]),
        .s21_axi_awlock(m_axi_awlock[21]),
        .s21_axi_awcache(m_axi_awcache[21]),
        .s21_axi_awprot(m_axi_awprot[21]),
        .s21_axi_awqos(m_axi_awqos[21]),
        .s21_axi_awuser(m_axi_awuser[21]),
        .s21_axi_awvalid(m_axi_awvalid[21]),
        .s21_axi_awready(m_axi_awready[21]),
        .s21_axi_wdata(m_axi_wdata[21]),
        .s21_axi_wstrb(m_axi_wstrb[21]),
        .s21_axi_wlast(m_axi_wlast[21]),
        .s21_axi_wuser(m_axi_wuser[21]),
        .s21_axi_wvalid(m_axi_wvalid[21]),
        .s21_axi_wready(m_axi_wready[21]),
        .s21_axi_bid(m_axi_bid[21]),
        .s21_axi_bresp(m_axi_bresp[21]),
        .s21_axi_buser(m_axi_buser[21]),
        .s21_axi_bvalid(m_axi_bvalid[21]),
        .s21_axi_bready(m_axi_bready[21]),
        .s21_axi_arid(m_axi_arid[21]),
        .s21_axi_araddr(m_axi_araddr[21]),
        .s21_axi_arlen(m_axi_arlen[21]),
        .s21_axi_arsize(m_axi_arsize[21]),
        .s21_axi_arburst(m_axi_arburst[21]),
        .s21_axi_arlock(m_axi_arlock[21]),
        .s21_axi_arcache(m_axi_arcache[21]),
        .s21_axi_arprot(m_axi_arprot[21]),
        .s21_axi_arqos(m_axi_arqos[21]),
        .s21_axi_aruser(m_axi_aruser[21]),
        .s21_axi_arvalid(m_axi_arvalid[21]),
        .s21_axi_arready(m_axi_arready[21]),
        .s21_axi_rid(m_axi_rid[21]),
        .s21_axi_rdata(m_axi_rdata[21]),
        .s21_axi_rresp(m_axi_rresp[21]),
        .s21_axi_rlast(m_axi_rlast[21]),
        .s21_axi_ruser(m_axi_ruser[21]),
        .s21_axi_rvalid(m_axi_rvalid[21]),
        .s21_axi_rready(m_axi_rready[21]),
        
        .s22_axi_awid(m_axi_awid[22]),
        .s22_axi_awaddr(m_axi_awaddr[22]),
        .s22_axi_awlen(m_axi_awlen[22]),
        .s22_axi_awsize(m_axi_awsize[22]),
        .s22_axi_awburst(m_axi_awburst[22]),
        .s22_axi_awlock(m_axi_awlock[22]),
        .s22_axi_awcache(m_axi_awcache[22]),
        .s22_axi_awprot(m_axi_awprot[22]),
        .s22_axi_awqos(m_axi_awqos[22]),
        .s22_axi_awuser(m_axi_awuser[22]),
        .s22_axi_awvalid(m_axi_awvalid[22]),
        .s22_axi_awready(m_axi_awready[22]),
        .s22_axi_wdata(m_axi_wdata[22]),
        .s22_axi_wstrb(m_axi_wstrb[22]),
        .s22_axi_wlast(m_axi_wlast[22]),
        .s22_axi_wuser(m_axi_wuser[22]),
        .s22_axi_wvalid(m_axi_wvalid[22]),
        .s22_axi_wready(m_axi_wready[22]),
        .s22_axi_bid(m_axi_bid[22]),
        .s22_axi_bresp(m_axi_bresp[22]),
        .s22_axi_buser(m_axi_buser[22]),
        .s22_axi_bvalid(m_axi_bvalid[22]),
        .s22_axi_bready(m_axi_bready[22]),
        .s22_axi_arid(m_axi_arid[22]),
        .s22_axi_araddr(m_axi_araddr[22]),
        .s22_axi_arlen(m_axi_arlen[22]),
        .s22_axi_arsize(m_axi_arsize[22]),
        .s22_axi_arburst(m_axi_arburst[22]),
        .s22_axi_arlock(m_axi_arlock[22]),
        .s22_axi_arcache(m_axi_arcache[22]),
        .s22_axi_arprot(m_axi_arprot[22]),
        .s22_axi_arqos(m_axi_arqos[22]),
        .s22_axi_aruser(m_axi_aruser[22]),
        .s22_axi_arvalid(m_axi_arvalid[22]),
        .s22_axi_arready(m_axi_arready[22]),
        .s22_axi_rid(m_axi_rid[22]),
        .s22_axi_rdata(m_axi_rdata[22]),
        .s22_axi_rresp(m_axi_rresp[22]),
        .s22_axi_rlast(m_axi_rlast[22]),
        .s22_axi_ruser(m_axi_ruser[22]),
        .s22_axi_rvalid(m_axi_rvalid[22]),
        .s22_axi_rready(m_axi_rready[22]),
        
        .s23_axi_awid(m_axi_awid[23]),
        .s23_axi_awaddr(m_axi_awaddr[23]),
        .s23_axi_awlen(m_axi_awlen[23]),
        .s23_axi_awsize(m_axi_awsize[23]),
        .s23_axi_awburst(m_axi_awburst[23]),
        .s23_axi_awlock(m_axi_awlock[23]),
        .s23_axi_awcache(m_axi_awcache[23]),
        .s23_axi_awprot(m_axi_awprot[23]),
        .s23_axi_awqos(m_axi_awqos[23]),
        .s23_axi_awuser(m_axi_awuser[23]),
        .s23_axi_awvalid(m_axi_awvalid[23]),
        .s23_axi_awready(m_axi_awready[23]),
        .s23_axi_wdata(m_axi_wdata[23]),
        .s23_axi_wstrb(m_axi_wstrb[23]),
        .s23_axi_wlast(m_axi_wlast[23]),
        .s23_axi_wuser(m_axi_wuser[23]),
        .s23_axi_wvalid(m_axi_wvalid[23]),
        .s23_axi_wready(m_axi_wready[23]),
        .s23_axi_bid(m_axi_bid[23]),
        .s23_axi_bresp(m_axi_bresp[23]),
        .s23_axi_buser(m_axi_buser[23]),
        .s23_axi_bvalid(m_axi_bvalid[23]),
        .s23_axi_bready(m_axi_bready[23]),
        .s23_axi_arid(m_axi_arid[23]),
        .s23_axi_araddr(m_axi_araddr[23]),
        .s23_axi_arlen(m_axi_arlen[23]),
        .s23_axi_arsize(m_axi_arsize[23]),
        .s23_axi_arburst(m_axi_arburst[23]),
        .s23_axi_arlock(m_axi_arlock[23]),
        .s23_axi_arcache(m_axi_arcache[23]),
        .s23_axi_arprot(m_axi_arprot[23]),
        .s23_axi_arqos(m_axi_arqos[23]),
        .s23_axi_aruser(m_axi_aruser[23]),
        .s23_axi_arvalid(m_axi_arvalid[23]),
        .s23_axi_arready(m_axi_arready[23]),
        .s23_axi_rid(m_axi_rid[23]),
        .s23_axi_rdata(m_axi_rdata[23]),
        .s23_axi_rresp(m_axi_rresp[23]),
        .s23_axi_rlast(m_axi_rlast[23]),
        .s23_axi_ruser(m_axi_ruser[23]),
        .s23_axi_rvalid(m_axi_rvalid[23]),
        .s23_axi_rready(m_axi_rready[23]),
        
        .s24_axi_awid(m_axi_awid[24]),
        .s24_axi_awaddr(m_axi_awaddr[24]),
        .s24_axi_awlen(m_axi_awlen[24]),
        .s24_axi_awsize(m_axi_awsize[24]),
        .s24_axi_awburst(m_axi_awburst[24]),
        .s24_axi_awlock(m_axi_awlock[24]),
        .s24_axi_awcache(m_axi_awcache[24]),
        .s24_axi_awprot(m_axi_awprot[24]),
        .s24_axi_awqos(m_axi_awqos[24]),
        .s24_axi_awuser(m_axi_awuser[24]),
        .s24_axi_awvalid(m_axi_awvalid[24]),
        .s24_axi_awready(m_axi_awready[24]),
        .s24_axi_wdata(m_axi_wdata[24]),
        .s24_axi_wstrb(m_axi_wstrb[24]),
        .s24_axi_wlast(m_axi_wlast[24]),
        .s24_axi_wuser(m_axi_wuser[24]),
        .s24_axi_wvalid(m_axi_wvalid[24]),
        .s24_axi_wready(m_axi_wready[24]),
        .s24_axi_bid(m_axi_bid[24]),
        .s24_axi_bresp(m_axi_bresp[24]),
        .s24_axi_buser(m_axi_buser[24]),
        .s24_axi_bvalid(m_axi_bvalid[24]),
        .s24_axi_bready(m_axi_bready[24]),
        .s24_axi_arid(m_axi_arid[24]),
        .s24_axi_araddr(m_axi_araddr[24]),
        .s24_axi_arlen(m_axi_arlen[24]),
        .s24_axi_arsize(m_axi_arsize[24]),
        .s24_axi_arburst(m_axi_arburst[24]),
        .s24_axi_arlock(m_axi_arlock[24]),
        .s24_axi_arcache(m_axi_arcache[24]),
        .s24_axi_arprot(m_axi_arprot[24]),
        .s24_axi_arqos(m_axi_arqos[24]),
        .s24_axi_aruser(m_axi_aruser[24]),
        .s24_axi_arvalid(m_axi_arvalid[24]),
        .s24_axi_arready(m_axi_arready[24]),
        .s24_axi_rid(m_axi_rid[24]),
        .s24_axi_rdata(m_axi_rdata[24]),
        .s24_axi_rresp(m_axi_rresp[24]),
        .s24_axi_rlast(m_axi_rlast[24]),
        .s24_axi_ruser(m_axi_ruser[24]),
        .s24_axi_rvalid(m_axi_rvalid[24]),
        .s24_axi_rready(m_axi_rready[24]),

        .s25_axi_awid(m_axi_awid[25]),
        .s25_axi_awaddr(m_axi_awaddr[25]),
        .s25_axi_awlen(m_axi_awlen[25]),
        .s25_axi_awsize(m_axi_awsize[25]),
        .s25_axi_awburst(m_axi_awburst[25]),
        .s25_axi_awlock(m_axi_awlock[25]),
        .s25_axi_awcache(m_axi_awcache[25]),
        .s25_axi_awprot(m_axi_awprot[25]),
        .s25_axi_awqos(m_axi_awqos[25]),
        .s25_axi_awuser(m_axi_awuser[25]),
        .s25_axi_awvalid(m_axi_awvalid[25]),
        .s25_axi_awready(m_axi_awready[25]),
        .s25_axi_wdata(m_axi_wdata[25]),
        .s25_axi_wstrb(m_axi_wstrb[25]),
        .s25_axi_wlast(m_axi_wlast[25]),
        .s25_axi_wuser(m_axi_wuser[25]),
        .s25_axi_wvalid(m_axi_wvalid[25]),
        .s25_axi_wready(m_axi_wready[25]),
        .s25_axi_bid(m_axi_bid[25]),
        .s25_axi_bresp(m_axi_bresp[25]),
        .s25_axi_buser(m_axi_buser[25]),
        .s25_axi_bvalid(m_axi_bvalid[25]),
        .s25_axi_bready(m_axi_bready[25]),
        .s25_axi_arid(m_axi_arid[25]),
        .s25_axi_araddr(m_axi_araddr[25]),
        .s25_axi_arlen(m_axi_arlen[25]),
        .s25_axi_arsize(m_axi_arsize[25]),
        .s25_axi_arburst(m_axi_arburst[25]),
        .s25_axi_arlock(m_axi_arlock[25]),
        .s25_axi_arcache(m_axi_arcache[25]),
        .s25_axi_arprot(m_axi_arprot[25]),
        .s25_axi_arqos(m_axi_arqos[25]),
        .s25_axi_aruser(m_axi_aruser[25]),
        .s25_axi_arvalid(m_axi_arvalid[25]),
        .s25_axi_arready(m_axi_arready[25]),
        .s25_axi_rid(m_axi_rid[25]),
        .s25_axi_rdata(m_axi_rdata[25]),
        .s25_axi_rresp(m_axi_rresp[25]),
        .s25_axi_rlast(m_axi_rlast[25]),
        .s25_axi_ruser(m_axi_ruser[25]),
        .s25_axi_rvalid(m_axi_rvalid[25]),
        .s25_axi_rready(m_axi_rready[25]),
        
        .s26_axi_awid(m_axi_awid[26]),
        .s26_axi_awaddr(m_axi_awaddr[26]),
        .s26_axi_awlen(m_axi_awlen[26]),
        .s26_axi_awsize(m_axi_awsize[26]),
        .s26_axi_awburst(m_axi_awburst[26]),
        .s26_axi_awlock(m_axi_awlock[26]),
        .s26_axi_awcache(m_axi_awcache[26]),
        .s26_axi_awprot(m_axi_awprot[26]),
        .s26_axi_awqos(m_axi_awqos[26]),
        .s26_axi_awuser(m_axi_awuser[26]),
        .s26_axi_awvalid(m_axi_awvalid[26]),
        .s26_axi_awready(m_axi_awready[26]),
        .s26_axi_wdata(m_axi_wdata[26]),
        .s26_axi_wstrb(m_axi_wstrb[26]),
        .s26_axi_wlast(m_axi_wlast[26]),
        .s26_axi_wuser(m_axi_wuser[26]),
        .s26_axi_wvalid(m_axi_wvalid[26]),
        .s26_axi_wready(m_axi_wready[26]),
        .s26_axi_bid(m_axi_bid[26]),
        .s26_axi_bresp(m_axi_bresp[26]),
        .s26_axi_buser(m_axi_buser[26]),
        .s26_axi_bvalid(m_axi_bvalid[26]),
        .s26_axi_bready(m_axi_bready[26]),
        .s26_axi_arid(m_axi_arid[26]),
        .s26_axi_araddr(m_axi_araddr[26]),
        .s26_axi_arlen(m_axi_arlen[26]),
        .s26_axi_arsize(m_axi_arsize[26]),
        .s26_axi_arburst(m_axi_arburst[26]),
        .s26_axi_arlock(m_axi_arlock[26]),
        .s26_axi_arcache(m_axi_arcache[26]),
        .s26_axi_arprot(m_axi_arprot[26]),
        .s26_axi_arqos(m_axi_arqos[26]),
        .s26_axi_aruser(m_axi_aruser[26]),
        .s26_axi_arvalid(m_axi_arvalid[26]),
        .s26_axi_arready(m_axi_arready[26]),
        .s26_axi_rid(m_axi_rid[26]),
        .s26_axi_rdata(m_axi_rdata[26]),
        .s26_axi_rresp(m_axi_rresp[26]),
        .s26_axi_rlast(m_axi_rlast[26]),
        .s26_axi_ruser(m_axi_ruser[26]),
        .s26_axi_rvalid(m_axi_rvalid[26]),
        .s26_axi_rready(m_axi_rready[26]),
        
        .s27_axi_awid(m_axi_awid[27]),
        .s27_axi_awaddr(m_axi_awaddr[27]),
        .s27_axi_awlen(m_axi_awlen[27]),
        .s27_axi_awsize(m_axi_awsize[27]),
        .s27_axi_awburst(m_axi_awburst[27]),
        .s27_axi_awlock(m_axi_awlock[27]),
        .s27_axi_awcache(m_axi_awcache[27]),
        .s27_axi_awprot(m_axi_awprot[27]),
        .s27_axi_awqos(m_axi_awqos[27]),
        .s27_axi_awuser(m_axi_awuser[27]),
        .s27_axi_awvalid(m_axi_awvalid[27]),
        .s27_axi_awready(m_axi_awready[27]),
        .s27_axi_wdata(m_axi_wdata[27]),
        .s27_axi_wstrb(m_axi_wstrb[27]),
        .s27_axi_wlast(m_axi_wlast[27]),
        .s27_axi_wuser(m_axi_wuser[27]),
        .s27_axi_wvalid(m_axi_wvalid[27]),
        .s27_axi_wready(m_axi_wready[27]),
        .s27_axi_bid(m_axi_bid[27]),
        .s27_axi_bresp(m_axi_bresp[27]),
        .s27_axi_buser(m_axi_buser[27]),
        .s27_axi_bvalid(m_axi_bvalid[27]),
        .s27_axi_bready(m_axi_bready[27]),
        .s27_axi_arid(m_axi_arid[27]),
        .s27_axi_araddr(m_axi_araddr[27]),
        .s27_axi_arlen(m_axi_arlen[27]),
        .s27_axi_arsize(m_axi_arsize[27]),
        .s27_axi_arburst(m_axi_arburst[27]),
        .s27_axi_arlock(m_axi_arlock[27]),
        .s27_axi_arcache(m_axi_arcache[27]),
        .s27_axi_arprot(m_axi_arprot[27]),
        .s27_axi_arqos(m_axi_arqos[27]),
        .s27_axi_aruser(m_axi_aruser[27]),
        .s27_axi_arvalid(m_axi_arvalid[27]),
        .s27_axi_arready(m_axi_arready[27]),
        .s27_axi_rid(m_axi_rid[27]),
        .s27_axi_rdata(m_axi_rdata[27]),
        .s27_axi_rresp(m_axi_rresp[27]),
        .s27_axi_rlast(m_axi_rlast[27]),
        .s27_axi_ruser(m_axi_ruser[27]),
        .s27_axi_rvalid(m_axi_rvalid[27]),
        .s27_axi_rready(m_axi_rready[27]),
      
        /*
         * AXI master interface
         */
        .m00_axi_awid(m_axi_noc_awid[0]),
        .m00_axi_awaddr(m_axi_noc_awaddr[0]),
        .m00_axi_awlen(m_axi_noc_awlen[0]),
        .m00_axi_awsize(m_axi_noc_awsize[0]),
        .m00_axi_awburst(m_axi_noc_awburst[0]),
        .m00_axi_awlock(m_axi_noc_awlock[0]),
        .m00_axi_awcache(m_axi_noc_awcache[0]),
        .m00_axi_awprot(m_axi_noc_awprot[0]),
        .m00_axi_awqos(m_axi_noc_awqos[0]),
        .m00_axi_awregion(m_axi_noc_awregion[0]),
        .m00_axi_awuser(m_axi_noc_awuser[0]),
        .m00_axi_awvalid(m_axi_noc_awvalid[0]),
        .m00_axi_awready(m_axi_noc_awready[0]),
        .m00_axi_wdata(m_axi_noc_wdata[0]),
        .m00_axi_wstrb(m_axi_noc_wstrb[0]),
        .m00_axi_wlast(m_axi_noc_wlast[0]),
        .m00_axi_wuser(m_axi_noc_wuser[0]),
        .m00_axi_wvalid(m_axi_noc_wvalid[0]),
        .m00_axi_wready(m_axi_noc_wready[0]),
        .m00_axi_bid(m_axi_noc_bid[0]),
        .m00_axi_bresp(m_axi_noc_bresp[0]),
        .m00_axi_buser(m_axi_noc_buser[0]),
        .m00_axi_bvalid(m_axi_noc_bvalid[0]),
        .m00_axi_bready(m_axi_noc_bready[0]),
        .m00_axi_arid(m_axi_noc_arid[0]),
        .m00_axi_araddr(m_axi_noc_araddr[0]),
        .m00_axi_arlen(m_axi_noc_arlen[0]),
        .m00_axi_arsize(m_axi_noc_arsize[0]),
        .m00_axi_arburst(m_axi_noc_arburst[0]),
        .m00_axi_arlock(m_axi_noc_arlock[0]),
        .m00_axi_arcache(m_axi_noc_arcache[0]),
        .m00_axi_arprot(m_axi_noc_arprot[0]),
        .m00_axi_arqos(m_axi_noc_arqos[0]),
        .m00_axi_arregion(m_axi_noc_arregion[0]),
        .m00_axi_aruser(m_axi_noc_aruser[0]),
        .m00_axi_arvalid(m_axi_noc_arvalid[0]),
        .m00_axi_arready(m_axi_noc_arready[0]),
        .m00_axi_rid(m_axi_noc_rid[0]),
        .m00_axi_rdata(m_axi_noc_rdata[0]),
        .m00_axi_rresp(m_axi_noc_rresp[0]),
        .m00_axi_rlast(m_axi_noc_rlast[0]),
        .m00_axi_ruser(m_axi_noc_ruser[0]),
        .m00_axi_rvalid(m_axi_noc_rvalid[0]),
        .m00_axi_rready(m_axi_noc_rready[0]),

        .m01_axi_awid(m_axi_noc_awid[1]),
        .m01_axi_awaddr(m_axi_noc_awaddr[1]),
        .m01_axi_awlen(m_axi_noc_awlen[1]),
        .m01_axi_awsize(m_axi_noc_awsize[1]),
        .m01_axi_awburst(m_axi_noc_awburst[1]),
        .m01_axi_awlock(m_axi_noc_awlock[1]),
        .m01_axi_awcache(m_axi_noc_awcache[1]),
        .m01_axi_awprot(m_axi_noc_awprot[1]),
        .m01_axi_awqos(m_axi_noc_awqos[1]),
        .m01_axi_awregion(m_axi_noc_awregion[1]),
        .m01_axi_awuser(m_axi_noc_awuser[1]),
        .m01_axi_awvalid(m_axi_noc_awvalid[1]),
        .m01_axi_awready(m_axi_noc_awready[1]),
        .m01_axi_wdata(m_axi_noc_wdata[1]),
        .m01_axi_wstrb(m_axi_noc_wstrb[1]),
        .m01_axi_wlast(m_axi_noc_wlast[1]),
        .m01_axi_wuser(m_axi_noc_wuser[1]),
        .m01_axi_wvalid(m_axi_noc_wvalid[1]),
        .m01_axi_wready(m_axi_noc_wready[1]),
        .m01_axi_bid(m_axi_noc_bid[1]),
        .m01_axi_bresp(m_axi_noc_bresp[1]),
        .m01_axi_buser(m_axi_noc_buser[1]),
        .m01_axi_bvalid(m_axi_noc_bvalid[1]),
        .m01_axi_bready(m_axi_noc_bready[1]),
        .m01_axi_arid(m_axi_noc_arid[1]),
        .m01_axi_araddr(m_axi_noc_araddr[1]),
        .m01_axi_arlen(m_axi_noc_arlen[1]),
        .m01_axi_arsize(m_axi_noc_arsize[1]),
        .m01_axi_arburst(m_axi_noc_arburst[1]),
        .m01_axi_arlock(m_axi_noc_arlock[1]),
        .m01_axi_arcache(m_axi_noc_arcache[1]),
        .m01_axi_arprot(m_axi_noc_arprot[1]),
        .m01_axi_arqos(m_axi_noc_arqos[1]),
        .m01_axi_arregion(m_axi_noc_arregion[1]),
        .m01_axi_aruser(m_axi_noc_aruser[1]),
        .m01_axi_arvalid(m_axi_noc_arvalid[1]),
        .m01_axi_arready(m_axi_noc_arready[1]),
        .m01_axi_rid(m_axi_noc_rid[1]),
        .m01_axi_rdata(m_axi_noc_rdata[1]),
        .m01_axi_rresp(m_axi_noc_rresp[1]),
        .m01_axi_rlast(m_axi_noc_rlast[1]),
        .m01_axi_ruser(m_axi_noc_ruser[1]),
        .m01_axi_rvalid(m_axi_noc_rvalid[1]),
        .m01_axi_rready(m_axi_noc_rready[1])
    );
    
    
    generate
        for (i = 0; i < 2; i = i + 1) begin : gen_noc_routers
            noc_router_module noc_router_module_inst (
                .clk(clk),
                .resetn(~rst),
        
                .s_axi_awaddr(m_axi_noc_awaddr[i]),
                .s_axi_awlen(m_axi_noc_awlen[i]),
                .s_axi_awsize(m_axi_noc_awsize[i]),
                .s_axi_awburst(m_axi_noc_awburst[i]),
                .s_axi_awvalid(m_axi_noc_awvalid[i]),
                .s_axi_awready(m_axi_noc_awready[i]),
                .s_axi_wdata(m_axi_noc_wdata[i]),
                .s_axi_wstrb(m_axi_noc_wstrb[i]),
                .s_axi_wlast(m_axi_noc_wlast[i]),
                .s_axi_wvalid(m_axi_noc_wvalid[i]),
                .s_axi_wready(m_axi_noc_wready[i]),
                .s_axi_bresp(m_axi_noc_bresp[i]),
                .s_axi_bvalid(m_axi_noc_bvalid[i]),
                .s_axi_bready(m_axi_noc_bready[i]),
                .s_axi_araddr(m_axi_noc_araddr[i]),
                .s_axi_arlen(m_axi_noc_arlen[i]),
                .s_axi_arsize(m_axi_noc_arsize[i]),
                .s_axi_arburst(m_axi_noc_arburst[i]),
                .s_axi_arvalid(m_axi_noc_arvalid[i]),
                .s_axi_arready(m_axi_noc_arready[i]),
                .s_axi_rdata(m_axi_noc_rdata[i]),
                .s_axi_rresp(m_axi_noc_rresp[i]),
                .s_axi_rlast(m_axi_noc_rlast[i]),
                .s_axi_rvalid(m_axi_noc_rvalid[i]),
                .s_axi_rready(m_axi_noc_rready[i])
            );

        end
    endgenerate

endmodule