`default_nettype wire 
`default_nettype tri

module simple_op(in,out);

    input in;
    output out;

    assign out = in;
	 
endmodule 