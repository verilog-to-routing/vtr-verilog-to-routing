module simple_op ( input signed in,
                                output out );

    assign out = in << 1;

endmodule
