
 module ex2BT16_fir(clk, In_X, Out_Y); 

 input clk;
 input [11:0] In_X; 
 output [28 :0] Out_Y; 

 reg [11:0] x0 ;

 wire [14:0] x1 ;
 wire [20:0] x5 ;
 wire [24:0] x23 ;
 wire [25:0] y27 ;
 wire [25:0] y43 ;
 wire [28:0] x28 ;
 wire [28:0] y32 ;
 wire [28:0] y38 ;
 wire [20:0] x6 ;
 wire [23:0] x16 ;
 wire [23:0] y25 ;
 wire [23:0] y45 ;
 wire [26:0] x17 ;
 wire [28:0] y31 ;
 wire [28:0] y39 ;
 wire [19:0] x10 ;
 wire [19:0] x10_0_1 ;
 wire [19:0] y20 ;
 wire [19:0] x10_1_1 ;
 wire [19:0] y50 ;
 wire [19:0] x11 ;
 wire [19:0] x11_0_1 ;
 wire [20:0] y22 ;
 wire [19:0] x11_1_1 ;
 wire [20:0] y48 ;
 wire [21:0] x12 ;
 wire [25:0] x22 ;
 wire [25:0] y26 ;
 wire [25:0] y44 ;
 wire [25:0] x13 ;
 wire [26:0] x24 ;
 wire [27:0] y30 ;
 wire [27:0] y40 ;
 wire [23:0] x18 ;
 wire [28:0] x26 ;
 wire [28:0] y29 ;
 wire [28:0] y41 ;
 wire [23:0] x19 ;
 wire [28:0] x27 ;
 wire [28:0] y33 ;
 wire [28:0] y37 ;
 wire [22:0] x20 ;
 wire [22:0] x20_0_1 ;
 wire [22:0] y23 ;
 wire [22:0] x20_1_1 ;
 wire [22:0] y47 ;
 wire [26:0] x21 ;
 wire [26:0] x21_0_1 ;
 wire [26:0] y28 ;
 wire [26:0] x21_1_1 ;
 wire [26:0] y42 ;
 wire [14:0] x1_13_1 ;
 wire [14:0] x1_13_2 ;
 wire [15:0] y18 ;
 wire [14:0] x1_14_1 ;
 wire [14:0] x1_14_2 ;
 wire [15:0] y52 ;
 wire [14:0] x2 ;
 wire [21:0] x4 ;
 wire [19:0] x14 ;
 wire [15:0] x3 ;
 wire [26:0] x15 ;
 wire [27:0] x25 ;
 wire [28:0] y34 ;
 wire [28:0] y36 ;
 wire [15:0] x3_4_1 ;
 wire [15:0] x3_4_2 ;
 wire [19:0] y21 ;
 wire [15:0] x3_5_1 ;
 wire [15:0] x3_5_2 ;
 wire [19:0] y49 ;
 wire [15:0] x7 ;
 wire [15:0] x7_0_1 ;
 wire [15:0] x7_0_2 ;
 wire [16:0] y19 ;
 wire [15:0] x7_1_1 ;
 wire [15:0] x7_1_2 ;
 wire [16:0] y51 ;
 wire [21:0] x8 ;
 wire [25:0] x9 ;
 wire [11:0] x0_21_1 ;
 wire [11:0] x0_21_2 ;
 wire [11:0] x0_21_3 ;
 wire [12:0] y17 ;
 wire [11:0] x0_22_1 ;
 wire [11:0] x0_22_2 ;
 wire [11:0] x0_22_3 ;
 wire [21:0] y24 ;
 wire [11:0] x0_23_1 ;
 wire [11:0] x0_23_2 ;
 wire [11:0] x0_23_3 ;
 wire [26:0] y35 ;
 wire [11:0] x0_24_1 ;
 wire [11:0] x0_24_2 ;
 wire [11:0] x0_24_3 ;
 wire [21:0] y46 ;
 wire [11:0] x0_25_1 ;
 wire [11:0] x0_25_2 ;
 wire [11:0] x0_25_3 ;
 wire [12:0] y53 ;
 wire [11:0] x29 ;
 wire [12:0] x30 ;
 wire [12:0] x30_1 ;
 wire [13:0] x31 ;
 wire [13:0] x31_1 ;
 wire [14:0] x32 ;
 wire [14:0] x32_1 ;
 wire [15:0] x33 ;
 wire [15:0] x33_1 ;
 wire [16:0] x34 ;
 wire [16:0] x34_1 ;
 wire [17:0] x35 ;
 wire [17:0] x35_1 ;
 wire [18:0] x36 ;
 wire [18:0] x36_1 ;
 wire [19:0] x37 ;
 wire [19:0] x37_1 ;
 wire [20:0] x38 ;
 wire [20:0] x38_1 ;
 wire [21:0] x39 ;
 wire [21:0] x39_1 ;
 wire [22:0] x40 ;
 wire [22:0] x40_1 ;
 wire [23:0] x41 ;
 wire [23:0] x41_1 ;
 wire [24:0] x42 ;
 wire [24:0] x42_1 ;
 wire [25:0] x43 ;
 wire [25:0] x43_1 ;
 wire [26:0] x44 ;
 wire [26:0] x44_1 ;
 wire [27:0] x45 ;
 wire [27:0] x45_1 ;
 wire [28:0] x46 ;
 wire [28:0] x46_1 ;
 wire [28:0] x47 ;
 wire [28:0] x47_1 ;
 wire [28:0] x48 ;
 wire [28:0] x48_1 ;
 wire [28:0] x49 ;
 wire [28:0] x49_1 ;
 wire [28:0] x50 ;
 wire [28:0] x50_1 ;
 wire [28:0] x51 ;
 wire [28:0] x51_1 ;
 wire [28:0] x52 ;
 wire [28:0] x52_1 ;
 wire [28:0] x53 ;
 wire [28:0] x53_1 ;
 wire [28:0] x54 ;
 wire [28:0] x54_1 ;
 wire [28:0] x55 ;
 wire [28:0] x55_1 ;
 wire [28:0] x56 ;
 wire [28:0] x56_1 ;
 wire [28:0] x57 ;
 wire [28:0] x57_1 ;
 wire [28:0] x58 ;
 wire [28:0] x58_1 ;
 wire [28:0] x59 ;
 wire [28:0] x59_1 ;
 wire [28:0] x60 ;
 wire [28:0] x60_1 ;
 wire [28:0] x61 ;
 wire [28:0] x61_1 ;
 wire [28:0] x62 ;
 wire [28:0] x62_1 ;
 wire [28:0] x63 ;
 wire [28:0] x63_1 ;
 wire [28:0] x64 ;
 wire [28:0] x64_1 ;
 wire [28:0] x65 ;
 wire [28:0] x65_1 ;
 wire [28:0] x66 ;
 wire [28:0] x66_1 ;
 wire [28:0] x67 ;
 wire [28:0] x67_1 ;
 wire [28:0] x68 ;
 wire [28:0] x68_1 ;
 wire [28:0] x69 ;
 wire [28:0] x69_1 ;
 wire [28:0] x70 ;
 wire [28:0] x70_1 ;
 wire [28:0] x71 ;
 wire [28:0] x71_1 ;
 wire [28:0] x72 ;
 wire [28:0] x72_1 ;
 wire [28:0] x73 ;
 wire [28:0] x73_1 ;
 wire [28:0] x74 ;
 wire [28:0] x74_1 ;
 wire [28:0] x75 ;
 wire [28:0] x75_1 ;
 wire [28:0] x76 ;
 wire [28:0] x76_1 ;
 wire [28:0] x77 ;
 wire [28:0] x77_1 ;
 wire [28:0] x78 ;
 wire [28:0] x78_1 ;
 wire [28:0] x79 ;
 wire [28:0] x79_1 ;
 wire [28:0] x80 ;
 wire [28:0] x80_1 ;
 wire [28:0] x81 ;
 wire [28:0] x81_1 ;
 wire [28:0] x82 ;
 wire [28:0] x82_1 ;
 wire [28:0] x83 ;
 wire [28:0] x83_1 ;
 wire [28:0] x84 ;
 wire [28:0] x84_1 ;
 wire [28:0] x85 ;
 wire [28:0] x85_1 ;
 wire [28:0] x86 ;
 wire [28:0] x86_1 ;
 wire [28:0] x87 ;
 wire [28:0] x87_1 ;
 wire [28:0] x88 ;
 wire [28:0] x88_1 ;
 wire [28:0] x89 ;
 wire [28:0] x89_1 ;
 wire [28:0] x90 ;
 wire [28:0] x90_1 ;
 wire [28:0] x91 ;
 wire [28:0] x91_1 ;
 wire [28:0] x92 ;
 wire [28:0] x92_1 ;
 wire [28:0] x93 ;
 wire [28:0] x93_1 ;
 wire [28:0] x94 ;
 wire [28:0] x94_1 ;
 wire [28:0] x95 ;
 wire [28:0] x95_1 ;
 wire [28:0] x96 ;
 wire [28:0] x96_1 ;
 wire [28:0] x97 ;
 wire [28:0] x97_1 ;
 wire [28:0] x98 ;
 wire [28:0] x98_1 ;
 wire [28:0] Out_Y_wire ;
 wire [11:0] y0 ;
 wire [11:0] y1 ;
 wire [11:0] y2 ;
 wire [11:0] y3 ;
 wire [11:0] y4 ;
 wire [11:0] y5 ;
 wire [11:0] y6 ;
 wire [11:0] y7 ;
 wire [11:0] y8 ;
 wire [11:0] y9 ;
 wire [11:0] y10 ;
 wire [11:0] y11 ;
 wire [11:0] y12 ;
 wire [11:0] y13 ;
 wire [11:0] y14 ;
 wire [11:0] y15 ;
 wire [11:0] y16 ;
 wire [11:0] y54 ;
 wire [11:0] y55 ;
 wire [11:0] y56 ;
 wire [11:0] y57 ;
 wire [11:0] y58 ;
 wire [11:0] y59 ;
 wire [11:0] y60 ;
 wire [11:0] y61 ;
 wire [11:0] y62 ;
 wire [11:0] y63 ;
 wire [11:0] y64 ;
 wire [11:0] y65 ;
 wire [11:0] y66 ;
 wire [11:0] y67 ;
 wire [11:0] y68 ;
 wire [11:0] y69 ;
 wire [11:0] y70 ;
 reg [11:0] Out_Y;

 reg [11:0] ZeroReg; 

 always @(posedge clk) 
 begin
 x0 <= In_X; 
 ZeroReg <= 12'b0 ;
 end 


 always @(posedge clk) 
 begin
 Out_Y = Out_Y_wire;
 end

 assign y0 = ZeroReg; 
 assign y1 = ZeroReg; 
 assign y2 = ZeroReg; 
 assign y3 = ZeroReg; 
 assign y4 = ZeroReg; 
 assign y5 = ZeroReg; 
 assign y6 = ZeroReg; 
 assign y7 = ZeroReg; 
 assign y8 = ZeroReg; 
 assign y9 = ZeroReg; 
 assign y10 = ZeroReg; 
 assign y11 = ZeroReg; 
 assign y12 = ZeroReg; 
 assign y13 = ZeroReg; 
 assign y14 = ZeroReg; 
 assign y15 = ZeroReg; 
 assign y16 = ZeroReg; 
 assign y54 = ZeroReg; 
 assign y55 = ZeroReg; 
 assign y56 = ZeroReg; 
 assign y57 = ZeroReg; 
 assign y58 = ZeroReg; 
 assign y59 = ZeroReg; 
 assign y60 = ZeroReg; 
 assign y61 = ZeroReg; 
 assign y62 = ZeroReg; 
 assign y63 = ZeroReg; 
 assign y64 = ZeroReg; 
 assign y65 = ZeroReg; 
 assign y66 = ZeroReg; 
 assign y67 = ZeroReg; 
 assign y68 = ZeroReg; 
 assign y69 = ZeroReg; 
 assign y70 = ZeroReg; 

 Subtractor14Bit Sub0(clk, { x0[11: 0], 2'b0 }, {x0[11],x0[11], x0[11: 0] }, x1); 


 Adder20Bit Adder0(clk,  {x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0] },  { x1[14: 0], 5'b0 },x5); 


 Subtractor19Bit Sub1(clk, { x1[14: 0], 4'b0 }, {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] }, x10); 

 Register20Bit Reg0 (clk,x10, x10_0_1 );
 Register20Bit Reg1 (clk,x10_0_1, y20 );
 Register20Bit Reg2 (clk,x10, x10_1_1 );
 Register20Bit Reg3 (clk,x10_1_1, y50 );

 Subtractor19Bit Sub2(clk, { x0[11: 0], 7'b0 }, {x1[14],x1[14],x1[14],x1[14], x1[14: 0] }, x11); 

 Register20Bit Reg4 (clk,x11, x11_0_1 );
 Register21Bit Reg5 (clk, {x11_0_1, 1'b0}, y22 );
 Register20Bit Reg6 (clk,x11, x11_1_1 );
 Register21Bit Reg7 (clk, {x11_1_1, 1'b0}, y48 );

 Subtractor21Bit Sub3(clk, { x1[14: 0], 6'b0 }, {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] }, x12); 


 Adder25Bit Adder1(clk,  { x1[14: 0], 10'b0 }, {x12[21],x12[21],x12[21], x12[21: 0]  }, x22); 

 Register26Bit Reg8 (clk,x22, y26 );
 Register26Bit Reg9 (clk,x22, y44 );

 Adder25Bit Adder2(clk,  { x0[11: 0], 13'b0 }, {x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0]  }, x13); 


 Adder23Bit Adder3(clk,  {x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0] },  { x1[14: 0], 8'b0 },x18); 

 Register15Bit Reg10 (clk,x1, x1_13_1 );
 Register15Bit Reg11 (clk,x1_13_1, x1_13_2 );
 Register16Bit Reg12 (clk, {x1_13_2, 1'b0}, y18 );
 Register15Bit Reg13 (clk,x1, x1_14_1 );
 Register15Bit Reg14 (clk,x1_14_1, x1_14_2 );
 Register16Bit Reg15 (clk, {x1_14_2, 1'b0}, y52 );

 Adder14Bit Adder4(clk,  {x0[11],x0[11], x0[11: 0] },  { x0[11: 0], 2'b0 },x2); 


 Subtractor21Bit Sub4(clk, {x2[14],x2[14],x2[14],x2[14],x2[14],x2[14], x2[14: 0] },  { x0[11: 0], 9'b0 },x4); 


 Adder28Bit Adder5(clk,  {x4[21],x4[21],x4[21],x4[21],x4[21],x4[21], x4[21: 0] },  { x18[23: 0], 4'b0 },x26); 

 Register29Bit Reg16 (clk,x26, y29 );
 Register29Bit Reg17 (clk,x26, y41 );

 Adder20Bit Adder6(clk,  {x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0] },  { x2[14: 0], 5'b0 },x6); 


 Subtractor23Bit Sub5(clk, { x0[11: 0], 11'b0 }, {x6[20],x6[20], x6[20: 0] }, x16); 

 Register24Bit Reg18 (clk,x16, y25 );
 Register24Bit Reg19 (clk,x16, y45 );

 Subtractor26Bit Sub6(clk, { x6[20: 0], 5'b0 }, {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] }, x17); 

 Register29Bit Reg20 (clk, {x17, 2'b0}, y31 );
 Register29Bit Reg21 (clk, {x17, 2'b0}, y39 );

 Subtractor19Bit Sub7(clk, { x2[14: 0], 4'b0 }, {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] }, x14); 


 Adder29Bit Adder7(clk,  { x5[20: 0], 8'b0 }, {x14[19],x14[19],x14[19],x14[19],x14[19],x14[19],x14[19],x14[19],x14[19], x14[19: 0]  }, x28); 

 Register29Bit Reg22 (clk,x28, y32 );
 Register29Bit Reg23 (clk,x28, y38 );

 Adder24Bit Adder8(clk,  { x2[14: 0], 9'b0 }, {x5[20],x5[20],x5[20], x5[20: 0]  }, x23); 

 Register26Bit Reg24 (clk, {x23, 1'b0}, y27 );
 Register26Bit Reg25 (clk, {x23, 1'b0}, y43 );

 Subtractor15Bit Sub8(clk, { x0[11: 0], 3'b0 }, {x0[11],x0[11],x0[11], x0[11: 0] }, x3); 


 Subtractor26Bit Sub9(clk, { x0[11: 0], 14'b0 }, {x3[15],x3[15],x3[15],x3[15],x3[15],x3[15],x3[15],x3[15],x3[15],x3[15], x3[15: 0] }, x15); 


 Subtractor27Bit Sub10(clk, { x15[26: 0] },  {x3[15],x3[15],x3[15],x3[15],x3[15], x3[15: 0], 6'b0 },x25); 

 Register29Bit Reg26 (clk, {x25, 1'b0}, y34 );
 Register29Bit Reg27 (clk, {x25, 1'b0}, y36 );

 Adder23Bit Adder9(clk,  {x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0] },  { x3[15: 0], 7'b0 },x19); 


 Subtractor29Bit Sub11(clk, { x19[23: 0], 5'b0 }, {x4[21],x4[21],x4[21],x4[21],x4[21],x4[21],x4[21], x4[21: 0] }, x27); 

 Register29Bit Reg28 (clk,x27, y33 );
 Register29Bit Reg29 (clk,x27, y37 );

 Subtractor26Bit Sub12(clk, { x13[25: 0] },  {x3[15],x3[15],x3[15],x3[15],x3[15],x3[15], x3[15: 0], 4'b0 },x24); 

 Register28Bit Reg30 (clk, {x24, 1'b0}, y30 );
 Register28Bit Reg31 (clk, {x24, 1'b0}, y40 );
 Register16Bit Reg32 (clk,x3, x3_4_1 );
 Register16Bit Reg33 (clk,x3_4_1, x3_4_2 );
 Register20Bit Reg34 (clk, {x3_4_2, 4'b0}, y21 );
 Register16Bit Reg35 (clk,x3, x3_5_1 );
 Register16Bit Reg36 (clk,x3_5_1, x3_5_2 );
 Register20Bit Reg37 (clk, {x3_5_2, 4'b0}, y49 );

 Adder15Bit Adder10(clk,  {x0[11],x0[11],x0[11], x0[11: 0] },  { x0[11: 0], 3'b0 },x7); 

 Register16Bit Reg38 (clk,x7, x7_0_1 );
 Register16Bit Reg39 (clk,x7_0_1, x7_0_2 );
 Register17Bit Reg40 (clk, {x7_0_2, 1'b0}, y19 );
 Register16Bit Reg41 (clk,x7, x7_1_1 );
 Register16Bit Reg42 (clk,x7_1_1, x7_1_2 );
 Register17Bit Reg43 (clk, {x7_1_2, 1'b0}, y51 );

 Subtractor21Bit Sub13(clk, { x0[11: 0], 9'b0 }, {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] }, x8); 


 Adder22Bit Adder11(clk,  {x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0], 2'b0 }, { x8[21: 0]  }, x20); 

 Register23Bit Reg44 (clk,x20, x20_0_1 );
 Register23Bit Reg45 (clk,x20_0_1, y23 );
 Register23Bit Reg46 (clk,x20, x20_1_1 );
 Register23Bit Reg47 (clk,x20_1_1, y47 );

 Subtractor25Bit Sub14(clk, { x0[11: 0], 13'b0 }, {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] }, x9); 


 Subtractor26Bit Sub15(clk, { x9[25: 0] },  {x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0], 3'b0 },x21); 

 Register27Bit Reg48 (clk,x21, x21_0_1 );
 Register27Bit Reg49 (clk,x21_0_1, y28 );
 Register27Bit Reg50 (clk,x21, x21_1_1 );
 Register27Bit Reg51 (clk,x21_1_1, y42 );
 Register12Bit Reg52 (clk,x0, x0_21_1 );
 Register12Bit Reg53 (clk,x0_21_1, x0_21_2 );
 Register12Bit Reg54 (clk,x0_21_2, x0_21_3 );
 Register13Bit Reg55 (clk, {x0_21_3, 1'b0}, y17 );
 Register12Bit Reg56 (clk,x0, x0_22_1 );
 Register12Bit Reg57 (clk,x0_22_1, x0_22_2 );
 Register12Bit Reg58 (clk,x0_22_2, x0_22_3 );
 Register22Bit Reg59 (clk, {x0_22_3, 10'b0}, y24 );
 Register12Bit Reg60 (clk,x0, x0_23_1 );
 Register12Bit Reg61 (clk,x0_23_1, x0_23_2 );
 Register12Bit Reg62 (clk,x0_23_2, x0_23_3 );
 Register27Bit Reg63 (clk, {x0_23_3, 15'b0}, y35 );
 Register12Bit Reg64 (clk,x0, x0_24_1 );
 Register12Bit Reg65 (clk,x0_24_1, x0_24_2 );
 Register12Bit Reg66 (clk,x0_24_2, x0_24_3 );
 Register22Bit Reg67 (clk, {x0_24_3, 10'b0}, y46 );
 Register12Bit Reg68 (clk,x0, x0_25_1 );
 Register12Bit Reg69 (clk,x0_25_1, x0_25_2 );
 Register12Bit Reg70 (clk,x0_25_2, x0_25_3 );
 Register13Bit Reg71 (clk, {x0_25_3, 1'b0}, y53 );
 Register12Bit Reg72 (clk,y0, x29 );

 Adder12Bit Adder12(clk,  { x29[11: 0] },  { y1[11: 0]  }, x30); 

 Register13Bit Reg73 (clk,x30, x30_1 );

 Adder13Bit Adder13(clk,  { x30_1[12: 0] },  {y2[11], y2[11: 0]  }, x31); 

 Register14Bit Reg74 (clk,x31, x31_1 );

 Adder14Bit Adder14(clk,  { x31_1[13: 0] },  {y3[11],y3[11], y3[11: 0]  }, x32); 

 Register15Bit Reg75 (clk,x32, x32_1 );

 Adder15Bit Adder15(clk,  { x32_1[14: 0] },  {y4[11],y4[11],y4[11], y4[11: 0]  }, x33); 

 Register16Bit Reg76 (clk,x33, x33_1 );

 Adder16Bit Adder16(clk,  { x33_1[15: 0] },  {y5[11],y5[11],y5[11],y5[11], y5[11: 0]  }, x34); 

 Register17Bit Reg77 (clk,x34, x34_1 );

 Adder17Bit Adder17(clk,  { x34_1[16: 0] },  {y6[11],y6[11],y6[11],y6[11],y6[11], y6[11: 0]  }, x35); 

 Register18Bit Reg78 (clk,x35, x35_1 );

 Adder18Bit Adder18(clk,  { x35_1[17: 0] },  {y7[11],y7[11],y7[11],y7[11],y7[11],y7[11], y7[11: 0]  }, x36); 

 Register19Bit Reg79 (clk,x36, x36_1 );

 Adder19Bit Adder19(clk,  { x36_1[18: 0] },  {y8[11],y8[11],y8[11],y8[11],y8[11],y8[11],y8[11], y8[11: 0]  }, x37); 

 Register20Bit Reg80 (clk,x37, x37_1 );

 Adder20Bit Adder20(clk,  { x37_1[19: 0] },  {y9[11],y9[11],y9[11],y9[11],y9[11],y9[11],y9[11],y9[11], y9[11: 0]  }, x38); 

 Register21Bit Reg81 (clk,x38, x38_1 );

 Adder21Bit Adder21(clk,  { x38_1[20: 0] },  {y10[11],y10[11],y10[11],y10[11],y10[11],y10[11],y10[11],y10[11],y10[11], y10[11: 0]  }, x39); 

 Register22Bit Reg82 (clk,x39, x39_1 );

 Adder22Bit Adder22(clk,  { x39_1[21: 0] },  {y11[11],y11[11],y11[11],y11[11],y11[11],y11[11],y11[11],y11[11],y11[11],y11[11], y11[11: 0]  }, x40); 

 Register23Bit Reg83 (clk,x40, x40_1 );

 Adder23Bit Adder23(clk,  { x40_1[22: 0] },  {y12[11],y12[11],y12[11],y12[11],y12[11],y12[11],y12[11],y12[11],y12[11],y12[11],y12[11], y12[11: 0]  }, x41); 

 Register24Bit Reg84 (clk,x41, x41_1 );

 Adder24Bit Adder24(clk,  { x41_1[23: 0] },  {y13[11],y13[11],y13[11],y13[11],y13[11],y13[11],y13[11],y13[11],y13[11],y13[11],y13[11],y13[11], y13[11: 0]  }, x42); 

 Register25Bit Reg85 (clk,x42, x42_1 );

 Adder25Bit Adder25(clk,  { x42_1[24: 0] },  {y14[11],y14[11],y14[11],y14[11],y14[11],y14[11],y14[11],y14[11],y14[11],y14[11],y14[11],y14[11],y14[11], y14[11: 0]  }, x43); 

 Register26Bit Reg86 (clk,x43, x43_1 );

 Adder26Bit Adder26(clk,  { x43_1[25: 0] },  {y15[11],y15[11],y15[11],y15[11],y15[11],y15[11],y15[11],y15[11],y15[11],y15[11],y15[11],y15[11],y15[11],y15[11], y15[11: 0]  }, x44); 

 Register27Bit Reg87 (clk,x44, x44_1 );

 Adder27Bit Adder27(clk,  { x44_1[26: 0] },  {y16[11],y16[11],y16[11],y16[11],y16[11],y16[11],y16[11],y16[11],y16[11],y16[11],y16[11],y16[11],y16[11],y16[11],y16[11], y16[11: 0]  }, x45); 

 Register28Bit Reg88 (clk,x45, x45_1 );

 Adder28Bit Adder28(clk,  { x45_1[27: 0] },  {y17[12],y17[12],y17[12],y17[12],y17[12],y17[12],y17[12],y17[12],y17[12],y17[12],y17[12],y17[12],y17[12],y17[12],y17[12], y17[12: 0]  }, x46); 

 Register29Bit Reg89 (clk,x46, x46_1 );

 Adder29Bit Adder29(clk,  { x46_1[28: 0] },  {y18[15],y18[15],y18[15],y18[15],y18[15],y18[15],y18[15],y18[15],y18[15],y18[15],y18[15],y18[15],y18[15], y18[15: 0]  }, x47); 

 Register29Bit Reg90 (clk,x47, x47_1 );

 Adder29Bit Adder30(clk,  { x47_1[28: 0] },  {y19[16],y19[16],y19[16],y19[16],y19[16],y19[16],y19[16],y19[16],y19[16],y19[16],y19[16],y19[16], y19[16: 0]  }, x48); 

 Register29Bit Reg91 (clk,x48, x48_1 );

 Adder29Bit Adder31(clk,  { x48_1[28: 0] },  {y20[19],y20[19],y20[19],y20[19],y20[19],y20[19],y20[19],y20[19],y20[19], y20[19: 0]  }, x49); 

 Register29Bit Reg92 (clk,x49, x49_1 );

 Adder29Bit Adder32(clk,  { x49_1[28: 0] },  {y21[19],y21[19],y21[19],y21[19],y21[19],y21[19],y21[19],y21[19],y21[19], y21[19: 0]  }, x50); 

 Register29Bit Reg93 (clk,x50, x50_1 );

 Adder29Bit Adder33(clk,  { x50_1[28: 0] },  {y22[20],y22[20],y22[20],y22[20],y22[20],y22[20],y22[20],y22[20], y22[20: 0]  }, x51); 

 Register29Bit Reg94 (clk,x51, x51_1 );

 Adder29Bit Adder34(clk,  { x51_1[28: 0] },  {y23[22],y23[22],y23[22],y23[22],y23[22],y23[22], y23[22: 0]  }, x52); 

 Register29Bit Reg95 (clk,x52, x52_1 );

 Adder29Bit Adder35(clk,  { x52_1[28: 0] },  {y24[21],y24[21],y24[21],y24[21],y24[21],y24[21],y24[21], y24[21: 0]  }, x53); 

 Register29Bit Reg96 (clk,x53, x53_1 );

 Adder29Bit Adder36(clk,  { x53_1[28: 0] },  {y25[23],y25[23],y25[23],y25[23],y25[23], y25[23: 0]  }, x54); 

 Register29Bit Reg97 (clk,x54, x54_1 );

 Adder29Bit Adder37(clk,  { x54_1[28: 0] },  {y26[25],y26[25],y26[25], y26[25: 0]  }, x55); 

 Register29Bit Reg98 (clk,x55, x55_1 );

 Adder29Bit Adder38(clk,  { x55_1[28: 0] },  {y27[25],y27[25],y27[25], y27[25: 0]  }, x56); 

 Register29Bit Reg99 (clk,x56, x56_1 );

 Adder29Bit Adder39(clk,  { x56_1[28: 0] },  {y28[26],y28[26], y28[26: 0]  }, x57); 

 Register29Bit Reg100 (clk,x57, x57_1 );

 Adder29Bit Adder40(clk,  { x57_1[28: 0] },  { y29[28: 0]  }, x58); 

 Register29Bit Reg101 (clk,x58, x58_1 );

 Adder29Bit Adder41(clk,  { x58_1[28: 0] },  {y30[27], y30[27: 0]  }, x59); 

 Register29Bit Reg102 (clk,x59, x59_1 );

 Adder29Bit Adder42(clk,  { x59_1[28: 0] },  { y31[28: 0]  }, x60); 

 Register29Bit Reg103 (clk,x60, x60_1 );

 Adder29Bit Adder43(clk,  { x60_1[28: 0] },  { y32[28: 0]  }, x61); 

 Register29Bit Reg104 (clk,x61, x61_1 );

 Adder29Bit Adder44(clk,  { x61_1[28: 0] },  { y33[28: 0]  }, x62); 

 Register29Bit Reg105 (clk,x62, x62_1 );

 Adder29Bit Adder45(clk,  { x62_1[28: 0] },  { y34[28: 0]  }, x63); 

 Register29Bit Reg106 (clk,x63, x63_1 );

 Adder29Bit Adder46(clk,  { x63_1[28: 0] },  {y35[26],y35[26], y35[26: 0]  }, x64); 

 Register29Bit Reg107 (clk,x64, x64_1 );

 Adder29Bit Adder47(clk,  { x64_1[28: 0] },  { y36[28: 0]  }, x65); 

 Register29Bit Reg108 (clk,x65, x65_1 );

 Adder29Bit Adder48(clk,  { x65_1[28: 0] },  { y37[28: 0]  }, x66); 

 Register29Bit Reg109 (clk,x66, x66_1 );

 Adder29Bit Adder49(clk,  { x66_1[28: 0] },  { y38[28: 0]  }, x67); 

 Register29Bit Reg110 (clk,x67, x67_1 );

 Adder29Bit Adder50(clk,  { x67_1[28: 0] },  { y39[28: 0]  }, x68); 

 Register29Bit Reg111 (clk,x68, x68_1 );

 Adder29Bit Adder51(clk,  { x68_1[28: 0] },  {y40[27], y40[27: 0]  }, x69); 

 Register29Bit Reg112 (clk,x69, x69_1 );

 Adder29Bit Adder52(clk,  { x69_1[28: 0] },  { y41[28: 0]  }, x70); 

 Register29Bit Reg113 (clk,x70, x70_1 );

 Adder29Bit Adder53(clk,  { x70_1[28: 0] },  {y42[26],y42[26], y42[26: 0]  }, x71); 

 Register29Bit Reg114 (clk,x71, x71_1 );

 Adder29Bit Adder54(clk,  { x71_1[28: 0] },  {y43[25],y43[25],y43[25], y43[25: 0]  }, x72); 

 Register29Bit Reg115 (clk,x72, x72_1 );

 Adder29Bit Adder55(clk,  { x72_1[28: 0] },  {y44[25],y44[25],y44[25], y44[25: 0]  }, x73); 

 Register29Bit Reg116 (clk,x73, x73_1 );

 Adder29Bit Adder56(clk,  { x73_1[28: 0] },  {y45[23],y45[23],y45[23],y45[23],y45[23], y45[23: 0]  }, x74); 

 Register29Bit Reg117 (clk,x74, x74_1 );

 Adder29Bit Adder57(clk,  { x74_1[28: 0] },  {y46[21],y46[21],y46[21],y46[21],y46[21],y46[21],y46[21], y46[21: 0]  }, x75); 

 Register29Bit Reg118 (clk,x75, x75_1 );

 Adder29Bit Adder58(clk,  { x75_1[28: 0] },  {y47[22],y47[22],y47[22],y47[22],y47[22],y47[22], y47[22: 0]  }, x76); 

 Register29Bit Reg119 (clk,x76, x76_1 );

 Adder29Bit Adder59(clk,  { x76_1[28: 0] },  {y48[20],y48[20],y48[20],y48[20],y48[20],y48[20],y48[20],y48[20], y48[20: 0]  }, x77); 

 Register29Bit Reg120 (clk,x77, x77_1 );

 Adder29Bit Adder60(clk,  { x77_1[28: 0] },  {y49[19],y49[19],y49[19],y49[19],y49[19],y49[19],y49[19],y49[19],y49[19], y49[19: 0]  }, x78); 

 Register29Bit Reg121 (clk,x78, x78_1 );

 Adder29Bit Adder61(clk,  { x78_1[28: 0] },  {y50[19],y50[19],y50[19],y50[19],y50[19],y50[19],y50[19],y50[19],y50[19], y50[19: 0]  }, x79); 

 Register29Bit Reg122 (clk,x79, x79_1 );

 Adder29Bit Adder62(clk,  { x79_1[28: 0] },  {y51[16],y51[16],y51[16],y51[16],y51[16],y51[16],y51[16],y51[16],y51[16],y51[16],y51[16],y51[16], y51[16: 0]  }, x80); 

 Register29Bit Reg123 (clk,x80, x80_1 );

 Adder29Bit Adder63(clk,  { x80_1[28: 0] },  {y52[15],y52[15],y52[15],y52[15],y52[15],y52[15],y52[15],y52[15],y52[15],y52[15],y52[15],y52[15],y52[15], y52[15: 0]  }, x81); 

 Register29Bit Reg124 (clk,x81, x81_1 );

 Adder29Bit Adder64(clk,  { x81_1[28: 0] },  {y53[12],y53[12],y53[12],y53[12],y53[12],y53[12],y53[12],y53[12],y53[12],y53[12],y53[12],y53[12],y53[12],y53[12],y53[12],y53[12], y53[12: 0]  }, x82); 

 Register29Bit Reg125 (clk,x82, x82_1 );

 Adder29Bit Adder65(clk,  { x82_1[28: 0] },  {y54[11],y54[11],y54[11],y54[11],y54[11],y54[11],y54[11],y54[11],y54[11],y54[11],y54[11],y54[11],y54[11],y54[11],y54[11],y54[11],y54[11], y54[11: 0]  }, x83); 

 Register29Bit Reg126 (clk,x83, x83_1 );

 Adder29Bit Adder66(clk,  { x83_1[28: 0] },  {y55[11],y55[11],y55[11],y55[11],y55[11],y55[11],y55[11],y55[11],y55[11],y55[11],y55[11],y55[11],y55[11],y55[11],y55[11],y55[11],y55[11], y55[11: 0]  }, x84); 

 Register29Bit Reg127 (clk,x84, x84_1 );

 Adder29Bit Adder67(clk,  { x84_1[28: 0] },  {y56[11],y56[11],y56[11],y56[11],y56[11],y56[11],y56[11],y56[11],y56[11],y56[11],y56[11],y56[11],y56[11],y56[11],y56[11],y56[11],y56[11], y56[11: 0]  }, x85); 

 Register29Bit Reg128 (clk,x85, x85_1 );

 Adder29Bit Adder68(clk,  { x85_1[28: 0] },  {y57[11],y57[11],y57[11],y57[11],y57[11],y57[11],y57[11],y57[11],y57[11],y57[11],y57[11],y57[11],y57[11],y57[11],y57[11],y57[11],y57[11], y57[11: 0]  }, x86); 

 Register29Bit Reg129 (clk,x86, x86_1 );

 Adder29Bit Adder69(clk,  { x86_1[28: 0] },  {y58[11],y58[11],y58[11],y58[11],y58[11],y58[11],y58[11],y58[11],y58[11],y58[11],y58[11],y58[11],y58[11],y58[11],y58[11],y58[11],y58[11], y58[11: 0]  }, x87); 

 Register29Bit Reg130 (clk,x87, x87_1 );

 Adder29Bit Adder70(clk,  { x87_1[28: 0] },  {y59[11],y59[11],y59[11],y59[11],y59[11],y59[11],y59[11],y59[11],y59[11],y59[11],y59[11],y59[11],y59[11],y59[11],y59[11],y59[11],y59[11], y59[11: 0]  }, x88); 

 Register29Bit Reg131 (clk,x88, x88_1 );

 Adder29Bit Adder71(clk,  { x88_1[28: 0] },  {y60[11],y60[11],y60[11],y60[11],y60[11],y60[11],y60[11],y60[11],y60[11],y60[11],y60[11],y60[11],y60[11],y60[11],y60[11],y60[11],y60[11], y60[11: 0]  }, x89); 

 Register29Bit Reg132 (clk,x89, x89_1 );

 Adder29Bit Adder72(clk,  { x89_1[28: 0] },  {y61[11],y61[11],y61[11],y61[11],y61[11],y61[11],y61[11],y61[11],y61[11],y61[11],y61[11],y61[11],y61[11],y61[11],y61[11],y61[11],y61[11], y61[11: 0]  }, x90); 

 Register29Bit Reg133 (clk,x90, x90_1 );

 Adder29Bit Adder73(clk,  { x90_1[28: 0] },  {y62[11],y62[11],y62[11],y62[11],y62[11],y62[11],y62[11],y62[11],y62[11],y62[11],y62[11],y62[11],y62[11],y62[11],y62[11],y62[11],y62[11], y62[11: 0]  }, x91); 

 Register29Bit Reg134 (clk,x91, x91_1 );

 Adder29Bit Adder74(clk,  { x91_1[28: 0] },  {y63[11],y63[11],y63[11],y63[11],y63[11],y63[11],y63[11],y63[11],y63[11],y63[11],y63[11],y63[11],y63[11],y63[11],y63[11],y63[11],y63[11], y63[11: 0]  }, x92); 

 Register29Bit Reg135 (clk,x92, x92_1 );

 Adder29Bit Adder75(clk,  { x92_1[28: 0] },  {y64[11],y64[11],y64[11],y64[11],y64[11],y64[11],y64[11],y64[11],y64[11],y64[11],y64[11],y64[11],y64[11],y64[11],y64[11],y64[11],y64[11], y64[11: 0]  }, x93); 

 Register29Bit Reg136 (clk,x93, x93_1 );

 Adder29Bit Adder76(clk,  { x93_1[28: 0] },  {y65[11],y65[11],y65[11],y65[11],y65[11],y65[11],y65[11],y65[11],y65[11],y65[11],y65[11],y65[11],y65[11],y65[11],y65[11],y65[11],y65[11], y65[11: 0]  }, x94); 

 Register29Bit Reg137 (clk,x94, x94_1 );

 Adder29Bit Adder77(clk,  { x94_1[28: 0] },  {y66[11],y66[11],y66[11],y66[11],y66[11],y66[11],y66[11],y66[11],y66[11],y66[11],y66[11],y66[11],y66[11],y66[11],y66[11],y66[11],y66[11], y66[11: 0]  }, x95); 

 Register29Bit Reg138 (clk,x95, x95_1 );

 Adder29Bit Adder78(clk,  { x95_1[28: 0] },  {y67[11],y67[11],y67[11],y67[11],y67[11],y67[11],y67[11],y67[11],y67[11],y67[11],y67[11],y67[11],y67[11],y67[11],y67[11],y67[11],y67[11], y67[11: 0]  }, x96); 

 Register29Bit Reg139 (clk,x96, x96_1 );

 Adder29Bit Adder79(clk,  { x96_1[28: 0] },  {y68[11],y68[11],y68[11],y68[11],y68[11],y68[11],y68[11],y68[11],y68[11],y68[11],y68[11],y68[11],y68[11],y68[11],y68[11],y68[11],y68[11], y68[11: 0]  }, x97); 

 Register29Bit Reg140 (clk,x97, x97_1 );

 Adder29Bit Adder80(clk,  { x97_1[28: 0] },  {y69[11],y69[11],y69[11],y69[11],y69[11],y69[11],y69[11],y69[11],y69[11],y69[11],y69[11],y69[11],y69[11],y69[11],y69[11],y69[11],y69[11], y69[11: 0]  }, x98); 

 Register29Bit Reg141 (clk,x98, x98_1 );

 Adder29Bit Adder81(clk,  { x98_1[28: 0] },  {y70[11],y70[11],y70[11],y70[11],y70[11],y70[11],y70[11],y70[11],y70[11],y70[11],y70[11],y70[11],y70[11],y70[11],y70[11],y70[11],y70[11], y70[11: 0]  }, Out_Y_wire); 

 endmodule 



module Adder20Bit (clk, In1, In2, AddOut);
 input clk;
 input [19:0] In1, In2; 

 output [20:0] AddOut;

 reg [20 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder24Bit (clk, In1, In2, AddOut);
 input clk;
 input [23:0] In1, In2; 

 output [24:0] AddOut;

 reg [24 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder29Bit (clk, In1, In2, AddOut);
 input clk;
 input [28:0] In1, In2; 

 output [28:0] AddOut;

 reg [28 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder25Bit (clk, In1, In2, AddOut);
 input clk;
 input [24:0] In1, In2; 

 output [25:0] AddOut;

 reg [25 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder23Bit (clk, In1, In2, AddOut);
 input clk;
 input [22:0] In1, In2; 

 output [23:0] AddOut;

 reg [23 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder28Bit (clk, In1, In2, AddOut);
 input clk;
 input [27:0] In1, In2; 

 output [28:0] AddOut;

 reg [28 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder22Bit (clk, In1, In2, AddOut);
 input clk;
 input [21:0] In1, In2; 

 output [22:0] AddOut;

 reg [22 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder14Bit (clk, In1, In2, AddOut);
 input clk;
 input [13:0] In1, In2; 

 output [14:0] AddOut;

 reg [14 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder15Bit (clk, In1, In2, AddOut);
 input clk;
 input [14:0] In1, In2; 

 output [15:0] AddOut;

 reg [15 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder12Bit (clk, In1, In2, AddOut);
 input clk;
 input [11:0] In1, In2; 

 output [12:0] AddOut;

 reg [12 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder13Bit (clk, In1, In2, AddOut);
 input clk;
 input [12:0] In1, In2; 

 output [13:0] AddOut;

 reg [13 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder16Bit (clk, In1, In2, AddOut);
 input clk;
 input [15:0] In1, In2; 

 output [16:0] AddOut;

 reg [16 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder17Bit (clk, In1, In2, AddOut);
 input clk;
 input [16:0] In1, In2; 

 output [17:0] AddOut;

 reg [17 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder18Bit (clk, In1, In2, AddOut);
 input clk;
 input [17:0] In1, In2; 

 output [18:0] AddOut;

 reg [18 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder19Bit (clk, In1, In2, AddOut);
 input clk;
 input [18:0] In1, In2; 

 output [19:0] AddOut;

 reg [19 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder21Bit (clk, In1, In2, AddOut);
 input clk;
 input [20:0] In1, In2; 

 output [21:0] AddOut;

 reg [21 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder26Bit (clk, In1, In2, AddOut);
 input clk;
 input [25:0] In1, In2; 

 output [26:0] AddOut;

 reg [26 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder27Bit (clk, In1, In2, AddOut);
 input clk;
 input [26:0] In1, In2; 

 output [27:0] AddOut;

 reg [27 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule



module Subtractor14Bit (clk, In1, In2, SubOut);
 input clk;
 input [13:0] In1, In2;
 output [14 :0] SubOut;

 reg [14 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule

module Subtractor23Bit (clk, In1, In2, SubOut);
 input clk;
 input [22:0] In1, In2;
 output [23 :0] SubOut;

 reg [23 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule

module Subtractor26Bit (clk, In1, In2, SubOut);
 input clk;
 input [25:0] In1, In2;
 output [26 :0] SubOut;

 reg [26 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule

module Subtractor19Bit (clk, In1, In2, SubOut);
 input clk;
 input [18:0] In1, In2;
 output [19 :0] SubOut;

 reg [19 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule

module Subtractor21Bit (clk, In1, In2, SubOut);
 input clk;
 input [20:0] In1, In2;
 output [21 :0] SubOut;

 reg [21 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule

module Subtractor29Bit (clk, In1, In2, SubOut);
 input clk;
 input [28:0] In1, In2;
 output [29 :0] SubOut;

 reg [29 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule

module Subtractor15Bit (clk, In1, In2, SubOut);
 input clk;
 input [14:0] In1, In2;
 output [15 :0] SubOut;

 reg [15 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule

module Subtractor27Bit (clk, In1, In2, SubOut);
 input clk;
 input [26:0] In1, In2;
 output [27 :0] SubOut;

 reg [27 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule

module Subtractor25Bit (clk, In1, In2, SubOut);
 input clk;
 input [24:0] In1, In2;
 output [25 :0] SubOut;

 reg [25 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule



module Register26Bit (clk, In1, RegOut);
 input clk;
 input [25:0] In1;
 output [25 :0] RegOut;

 reg [25 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register29Bit (clk, In1, RegOut);
 input clk;
 input [28:0] In1;
 output [28 :0] RegOut;

 reg [28 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register24Bit (clk, In1, RegOut);
 input clk;
 input [23:0] In1;
 output [23 :0] RegOut;

 reg [23 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register20Bit (clk, In1, RegOut);
 input clk;
 input [19:0] In1;
 output [19 :0] RegOut;

 reg [19 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register21Bit (clk, In1, RegOut);
 input clk;
 input [20:0] In1;
 output [20 :0] RegOut;

 reg [20 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register28Bit (clk, In1, RegOut);
 input clk;
 input [27:0] In1;
 output [27 :0] RegOut;

 reg [27 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register23Bit (clk, In1, RegOut);
 input clk;
 input [22:0] In1;
 output [22 :0] RegOut;

 reg [22 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register27Bit (clk, In1, RegOut);
 input clk;
 input [26:0] In1;
 output [26 :0] RegOut;

 reg [26 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register15Bit (clk, In1, RegOut);
 input clk;
 input [14:0] In1;
 output [14 :0] RegOut;

 reg [14 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register16Bit (clk, In1, RegOut);
 input clk;
 input [15:0] In1;
 output [15 :0] RegOut;

 reg [15 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register17Bit (clk, In1, RegOut);
 input clk;
 input [16:0] In1;
 output [16 :0] RegOut;

 reg [16 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register12Bit (clk, In1, RegOut);
 input clk;
 input [11:0] In1;
 output [11 :0] RegOut;

 reg [11 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register13Bit (clk, In1, RegOut);
 input clk;
 input [12:0] In1;
 output [12 :0] RegOut;

 reg [12 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register22Bit (clk, In1, RegOut);
 input clk;
 input [21:0] In1;
 output [21 :0] RegOut;

 reg [21 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register14Bit (clk, In1, RegOut);
 input clk;
 input [13:0] In1;
 output [13 :0] RegOut;

 reg [13 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register18Bit (clk, In1, RegOut);
 input clk;
 input [17:0] In1;
 output [17 :0] RegOut;

 reg [17 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register19Bit (clk, In1, RegOut);
 input clk;
 input [18:0] In1;
 output [18 :0] RegOut;

 reg [18 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register25Bit (clk, In1, RegOut);
 input clk;
 input [24:0] In1;
 output [24 :0] RegOut;

 reg [24 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule


