module and_primitive(
	out
);
	/*  input declaration	*/
	wire   a;
	wire   b;

	/*	output declaration	*/
	output	out;

    assign out = a&b; 

endmodule