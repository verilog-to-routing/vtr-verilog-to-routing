module simple_op(a,b);
input unsigned [3:0] a;
output signed [5:0] b;

assign b = a;

endmodule