/*
 * This header file provides definitions for ch_intrinsic_modified.v
 * located at: 
 *      vtr_flow/benchmarks/hdl_include/ch_intrinsic_modified.v
*/
`define MEMORY_CONTROLLER_TAGS 1
`define MEMORY_CONTROLLER_TAG_SIZE 1
`define TAG__str 1'b0