/*

Copyright (c) 2020 Alex Forencich

Permission is hereby granted, free of charge, to any person obtaining a copy
of this software and associated documentation files (the "Software"), to deal
in the Software without restriction, including without limitation the rights
to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
copies of the Software, and to permit persons to whom the Software is
furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in
all copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY
FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
THE SOFTWARE.

*/

// Language: Verilog 2001

`resetall
`timescale 1ns / 1ps
`default_nettype none

/*
 * AXI4 28x2 interconnect (wrapper)
 */
module axi_interconnect_wrap_28x2 #
(
    parameter DATA_WIDTH = 32,
    parameter ADDR_WIDTH = 32,
    parameter STRB_WIDTH = (DATA_WIDTH/8),
    parameter ID_WIDTH = 8,
    parameter AWUSER_ENABLE = 0,
    parameter AWUSER_WIDTH = 1,
    parameter WUSER_ENABLE = 0,
    parameter WUSER_WIDTH = 1,
    parameter BUSER_ENABLE = 0,
    parameter BUSER_WIDTH = 1,
    parameter ARUSER_ENABLE = 0,
    parameter ARUSER_WIDTH = 1,
    parameter RUSER_ENABLE = 0,
    parameter RUSER_WIDTH = 1,
    parameter FORWARD_ID = 0,
    parameter M_REGIONS = 1,
    parameter M00_BASE_ADDR = 0,
    parameter M00_ADDR_WIDTH = {M_REGIONS{32'd24}},
    parameter M00_CONNECT_READ = 28'b1111111111111111111111111111,
    parameter M00_CONNECT_WRITE = 28'b1111111111111111111111111111,
    parameter M00_SECURE = 1'b0,
    parameter M01_BASE_ADDR = 0,
    parameter M01_ADDR_WIDTH = {M_REGIONS{32'd24}},
    parameter M01_CONNECT_READ = 28'b1111111111111111111111111111,
    parameter M01_CONNECT_WRITE = 28'b1111111111111111111111111111,
    parameter M01_SECURE = 1'b0
)
(
    input  wire                     clk,
    input  wire                     rst,

    /*
     * AXI slave interface
     */
    input  wire [ID_WIDTH-1:0]      s00_axi_awid,
    input  wire [ADDR_WIDTH-1:0]    s00_axi_awaddr,
    input  wire [7:0]               s00_axi_awlen,
    input  wire [2:0]               s00_axi_awsize,
    input  wire [1:0]               s00_axi_awburst,
    input  wire                     s00_axi_awlock,
    input  wire [3:0]               s00_axi_awcache,
    input  wire [2:0]               s00_axi_awprot,
    input  wire [3:0]               s00_axi_awqos,
    input  wire [AWUSER_WIDTH-1:0]  s00_axi_awuser,
    input  wire                     s00_axi_awvalid,
    output wire                     s00_axi_awready,
    input  wire [DATA_WIDTH-1:0]    s00_axi_wdata,
    input  wire [STRB_WIDTH-1:0]    s00_axi_wstrb,
    input  wire                     s00_axi_wlast,
    input  wire [WUSER_WIDTH-1:0]   s00_axi_wuser,
    input  wire                     s00_axi_wvalid,
    output wire                     s00_axi_wready,
    output wire [ID_WIDTH-1:0]      s00_axi_bid,
    output wire [1:0]               s00_axi_bresp,
    output wire [BUSER_WIDTH-1:0]   s00_axi_buser,
    output wire                     s00_axi_bvalid,
    input  wire                     s00_axi_bready,
    input  wire [ID_WIDTH-1:0]      s00_axi_arid,
    input  wire [ADDR_WIDTH-1:0]    s00_axi_araddr,
    input  wire [7:0]               s00_axi_arlen,
    input  wire [2:0]               s00_axi_arsize,
    input  wire [1:0]               s00_axi_arburst,
    input  wire                     s00_axi_arlock,
    input  wire [3:0]               s00_axi_arcache,
    input  wire [2:0]               s00_axi_arprot,
    input  wire [3:0]               s00_axi_arqos,
    input  wire [ARUSER_WIDTH-1:0]  s00_axi_aruser,
    input  wire                     s00_axi_arvalid,
    output wire                     s00_axi_arready,
    output wire [ID_WIDTH-1:0]      s00_axi_rid,
    output wire [DATA_WIDTH-1:0]    s00_axi_rdata,
    output wire [1:0]               s00_axi_rresp,
    output wire                     s00_axi_rlast,
    output wire [RUSER_WIDTH-1:0]   s00_axi_ruser,
    output wire                     s00_axi_rvalid,
    input  wire                     s00_axi_rready,

    input  wire [ID_WIDTH-1:0]      s01_axi_awid,
    input  wire [ADDR_WIDTH-1:0]    s01_axi_awaddr,
    input  wire [7:0]               s01_axi_awlen,
    input  wire [2:0]               s01_axi_awsize,
    input  wire [1:0]               s01_axi_awburst,
    input  wire                     s01_axi_awlock,
    input  wire [3:0]               s01_axi_awcache,
    input  wire [2:0]               s01_axi_awprot,
    input  wire [3:0]               s01_axi_awqos,
    input  wire [AWUSER_WIDTH-1:0]  s01_axi_awuser,
    input  wire                     s01_axi_awvalid,
    output wire                     s01_axi_awready,
    input  wire [DATA_WIDTH-1:0]    s01_axi_wdata,
    input  wire [STRB_WIDTH-1:0]    s01_axi_wstrb,
    input  wire                     s01_axi_wlast,
    input  wire [WUSER_WIDTH-1:0]   s01_axi_wuser,
    input  wire                     s01_axi_wvalid,
    output wire                     s01_axi_wready,
    output wire [ID_WIDTH-1:0]      s01_axi_bid,
    output wire [1:0]               s01_axi_bresp,
    output wire [BUSER_WIDTH-1:0]   s01_axi_buser,
    output wire                     s01_axi_bvalid,
    input  wire                     s01_axi_bready,
    input  wire [ID_WIDTH-1:0]      s01_axi_arid,
    input  wire [ADDR_WIDTH-1:0]    s01_axi_araddr,
    input  wire [7:0]               s01_axi_arlen,
    input  wire [2:0]               s01_axi_arsize,
    input  wire [1:0]               s01_axi_arburst,
    input  wire                     s01_axi_arlock,
    input  wire [3:0]               s01_axi_arcache,
    input  wire [2:0]               s01_axi_arprot,
    input  wire [3:0]               s01_axi_arqos,
    input  wire [ARUSER_WIDTH-1:0]  s01_axi_aruser,
    input  wire                     s01_axi_arvalid,
    output wire                     s01_axi_arready,
    output wire [ID_WIDTH-1:0]      s01_axi_rid,
    output wire [DATA_WIDTH-1:0]    s01_axi_rdata,
    output wire [1:0]               s01_axi_rresp,
    output wire                     s01_axi_rlast,
    output wire [RUSER_WIDTH-1:0]   s01_axi_ruser,
    output wire                     s01_axi_rvalid,
    input  wire                     s01_axi_rready,

    input  wire [ID_WIDTH-1:0]      s02_axi_awid,
    input  wire [ADDR_WIDTH-1:0]    s02_axi_awaddr,
    input  wire [7:0]               s02_axi_awlen,
    input  wire [2:0]               s02_axi_awsize,
    input  wire [1:0]               s02_axi_awburst,
    input  wire                     s02_axi_awlock,
    input  wire [3:0]               s02_axi_awcache,
    input  wire [2:0]               s02_axi_awprot,
    input  wire [3:0]               s02_axi_awqos,
    input  wire [AWUSER_WIDTH-1:0]  s02_axi_awuser,
    input  wire                     s02_axi_awvalid,
    output wire                     s02_axi_awready,
    input  wire [DATA_WIDTH-1:0]    s02_axi_wdata,
    input  wire [STRB_WIDTH-1:0]    s02_axi_wstrb,
    input  wire                     s02_axi_wlast,
    input  wire [WUSER_WIDTH-1:0]   s02_axi_wuser,
    input  wire                     s02_axi_wvalid,
    output wire                     s02_axi_wready,
    output wire [ID_WIDTH-1:0]      s02_axi_bid,
    output wire [1:0]               s02_axi_bresp,
    output wire [BUSER_WIDTH-1:0]   s02_axi_buser,
    output wire                     s02_axi_bvalid,
    input  wire                     s02_axi_bready,
    input  wire [ID_WIDTH-1:0]      s02_axi_arid,
    input  wire [ADDR_WIDTH-1:0]    s02_axi_araddr,
    input  wire [7:0]               s02_axi_arlen,
    input  wire [2:0]               s02_axi_arsize,
    input  wire [1:0]               s02_axi_arburst,
    input  wire                     s02_axi_arlock,
    input  wire [3:0]               s02_axi_arcache,
    input  wire [2:0]               s02_axi_arprot,
    input  wire [3:0]               s02_axi_arqos,
    input  wire [ARUSER_WIDTH-1:0]  s02_axi_aruser,
    input  wire                     s02_axi_arvalid,
    output wire                     s02_axi_arready,
    output wire [ID_WIDTH-1:0]      s02_axi_rid,
    output wire [DATA_WIDTH-1:0]    s02_axi_rdata,
    output wire [1:0]               s02_axi_rresp,
    output wire                     s02_axi_rlast,
    output wire [RUSER_WIDTH-1:0]   s02_axi_ruser,
    output wire                     s02_axi_rvalid,
    input  wire                     s02_axi_rready,

    input  wire [ID_WIDTH-1:0]      s03_axi_awid,
    input  wire [ADDR_WIDTH-1:0]    s03_axi_awaddr,
    input  wire [7:0]               s03_axi_awlen,
    input  wire [2:0]               s03_axi_awsize,
    input  wire [1:0]               s03_axi_awburst,
    input  wire                     s03_axi_awlock,
    input  wire [3:0]               s03_axi_awcache,
    input  wire [2:0]               s03_axi_awprot,
    input  wire [3:0]               s03_axi_awqos,
    input  wire [AWUSER_WIDTH-1:0]  s03_axi_awuser,
    input  wire                     s03_axi_awvalid,
    output wire                     s03_axi_awready,
    input  wire [DATA_WIDTH-1:0]    s03_axi_wdata,
    input  wire [STRB_WIDTH-1:0]    s03_axi_wstrb,
    input  wire                     s03_axi_wlast,
    input  wire [WUSER_WIDTH-1:0]   s03_axi_wuser,
    input  wire                     s03_axi_wvalid,
    output wire                     s03_axi_wready,
    output wire [ID_WIDTH-1:0]      s03_axi_bid,
    output wire [1:0]               s03_axi_bresp,
    output wire [BUSER_WIDTH-1:0]   s03_axi_buser,
    output wire                     s03_axi_bvalid,
    input  wire                     s03_axi_bready,
    input  wire [ID_WIDTH-1:0]      s03_axi_arid,
    input  wire [ADDR_WIDTH-1:0]    s03_axi_araddr,
    input  wire [7:0]               s03_axi_arlen,
    input  wire [2:0]               s03_axi_arsize,
    input  wire [1:0]               s03_axi_arburst,
    input  wire                     s03_axi_arlock,
    input  wire [3:0]               s03_axi_arcache,
    input  wire [2:0]               s03_axi_arprot,
    input  wire [3:0]               s03_axi_arqos,
    input  wire [ARUSER_WIDTH-1:0]  s03_axi_aruser,
    input  wire                     s03_axi_arvalid,
    output wire                     s03_axi_arready,
    output wire [ID_WIDTH-1:0]      s03_axi_rid,
    output wire [DATA_WIDTH-1:0]    s03_axi_rdata,
    output wire [1:0]               s03_axi_rresp,
    output wire                     s03_axi_rlast,
    output wire [RUSER_WIDTH-1:0]   s03_axi_ruser,
    output wire                     s03_axi_rvalid,
    input  wire                     s03_axi_rready,

    input  wire [ID_WIDTH-1:0]      s04_axi_awid,
    input  wire [ADDR_WIDTH-1:0]    s04_axi_awaddr,
    input  wire [7:0]               s04_axi_awlen,
    input  wire [2:0]               s04_axi_awsize,
    input  wire [1:0]               s04_axi_awburst,
    input  wire                     s04_axi_awlock,
    input  wire [3:0]               s04_axi_awcache,
    input  wire [2:0]               s04_axi_awprot,
    input  wire [3:0]               s04_axi_awqos,
    input  wire [AWUSER_WIDTH-1:0]  s04_axi_awuser,
    input  wire                     s04_axi_awvalid,
    output wire                     s04_axi_awready,
    input  wire [DATA_WIDTH-1:0]    s04_axi_wdata,
    input  wire [STRB_WIDTH-1:0]    s04_axi_wstrb,
    input  wire                     s04_axi_wlast,
    input  wire [WUSER_WIDTH-1:0]   s04_axi_wuser,
    input  wire                     s04_axi_wvalid,
    output wire                     s04_axi_wready,
    output wire [ID_WIDTH-1:0]      s04_axi_bid,
    output wire [1:0]               s04_axi_bresp,
    output wire [BUSER_WIDTH-1:0]   s04_axi_buser,
    output wire                     s04_axi_bvalid,
    input  wire                     s04_axi_bready,
    input  wire [ID_WIDTH-1:0]      s04_axi_arid,
    input  wire [ADDR_WIDTH-1:0]    s04_axi_araddr,
    input  wire [7:0]               s04_axi_arlen,
    input  wire [2:0]               s04_axi_arsize,
    input  wire [1:0]               s04_axi_arburst,
    input  wire                     s04_axi_arlock,
    input  wire [3:0]               s04_axi_arcache,
    input  wire [2:0]               s04_axi_arprot,
    input  wire [3:0]               s04_axi_arqos,
    input  wire [ARUSER_WIDTH-1:0]  s04_axi_aruser,
    input  wire                     s04_axi_arvalid,
    output wire                     s04_axi_arready,
    output wire [ID_WIDTH-1:0]      s04_axi_rid,
    output wire [DATA_WIDTH-1:0]    s04_axi_rdata,
    output wire [1:0]               s04_axi_rresp,
    output wire                     s04_axi_rlast,
    output wire [RUSER_WIDTH-1:0]   s04_axi_ruser,
    output wire                     s04_axi_rvalid,
    input  wire                     s04_axi_rready,

    input  wire [ID_WIDTH-1:0]      s05_axi_awid,
    input  wire [ADDR_WIDTH-1:0]    s05_axi_awaddr,
    input  wire [7:0]               s05_axi_awlen,
    input  wire [2:0]               s05_axi_awsize,
    input  wire [1:0]               s05_axi_awburst,
    input  wire                     s05_axi_awlock,
    input  wire [3:0]               s05_axi_awcache,
    input  wire [2:0]               s05_axi_awprot,
    input  wire [3:0]               s05_axi_awqos,
    input  wire [AWUSER_WIDTH-1:0]  s05_axi_awuser,
    input  wire                     s05_axi_awvalid,
    output wire                     s05_axi_awready,
    input  wire [DATA_WIDTH-1:0]    s05_axi_wdata,
    input  wire [STRB_WIDTH-1:0]    s05_axi_wstrb,
    input  wire                     s05_axi_wlast,
    input  wire [WUSER_WIDTH-1:0]   s05_axi_wuser,
    input  wire                     s05_axi_wvalid,
    output wire                     s05_axi_wready,
    output wire [ID_WIDTH-1:0]      s05_axi_bid,
    output wire [1:0]               s05_axi_bresp,
    output wire [BUSER_WIDTH-1:0]   s05_axi_buser,
    output wire                     s05_axi_bvalid,
    input  wire                     s05_axi_bready,
    input  wire [ID_WIDTH-1:0]      s05_axi_arid,
    input  wire [ADDR_WIDTH-1:0]    s05_axi_araddr,
    input  wire [7:0]               s05_axi_arlen,
    input  wire [2:0]               s05_axi_arsize,
    input  wire [1:0]               s05_axi_arburst,
    input  wire                     s05_axi_arlock,
    input  wire [3:0]               s05_axi_arcache,
    input  wire [2:0]               s05_axi_arprot,
    input  wire [3:0]               s05_axi_arqos,
    input  wire [ARUSER_WIDTH-1:0]  s05_axi_aruser,
    input  wire                     s05_axi_arvalid,
    output wire                     s05_axi_arready,
    output wire [ID_WIDTH-1:0]      s05_axi_rid,
    output wire [DATA_WIDTH-1:0]    s05_axi_rdata,
    output wire [1:0]               s05_axi_rresp,
    output wire                     s05_axi_rlast,
    output wire [RUSER_WIDTH-1:0]   s05_axi_ruser,
    output wire                     s05_axi_rvalid,
    input  wire                     s05_axi_rready,

    input  wire [ID_WIDTH-1:0]      s06_axi_awid,
    input  wire [ADDR_WIDTH-1:0]    s06_axi_awaddr,
    input  wire [7:0]               s06_axi_awlen,
    input  wire [2:0]               s06_axi_awsize,
    input  wire [1:0]               s06_axi_awburst,
    input  wire                     s06_axi_awlock,
    input  wire [3:0]               s06_axi_awcache,
    input  wire [2:0]               s06_axi_awprot,
    input  wire [3:0]               s06_axi_awqos,
    input  wire [AWUSER_WIDTH-1:0]  s06_axi_awuser,
    input  wire                     s06_axi_awvalid,
    output wire                     s06_axi_awready,
    input  wire [DATA_WIDTH-1:0]    s06_axi_wdata,
    input  wire [STRB_WIDTH-1:0]    s06_axi_wstrb,
    input  wire                     s06_axi_wlast,
    input  wire [WUSER_WIDTH-1:0]   s06_axi_wuser,
    input  wire                     s06_axi_wvalid,
    output wire                     s06_axi_wready,
    output wire [ID_WIDTH-1:0]      s06_axi_bid,
    output wire [1:0]               s06_axi_bresp,
    output wire [BUSER_WIDTH-1:0]   s06_axi_buser,
    output wire                     s06_axi_bvalid,
    input  wire                     s06_axi_bready,
    input  wire [ID_WIDTH-1:0]      s06_axi_arid,
    input  wire [ADDR_WIDTH-1:0]    s06_axi_araddr,
    input  wire [7:0]               s06_axi_arlen,
    input  wire [2:0]               s06_axi_arsize,
    input  wire [1:0]               s06_axi_arburst,
    input  wire                     s06_axi_arlock,
    input  wire [3:0]               s06_axi_arcache,
    input  wire [2:0]               s06_axi_arprot,
    input  wire [3:0]               s06_axi_arqos,
    input  wire [ARUSER_WIDTH-1:0]  s06_axi_aruser,
    input  wire                     s06_axi_arvalid,
    output wire                     s06_axi_arready,
    output wire [ID_WIDTH-1:0]      s06_axi_rid,
    output wire [DATA_WIDTH-1:0]    s06_axi_rdata,
    output wire [1:0]               s06_axi_rresp,
    output wire                     s06_axi_rlast,
    output wire [RUSER_WIDTH-1:0]   s06_axi_ruser,
    output wire                     s06_axi_rvalid,
    input  wire                     s06_axi_rready,

    input  wire [ID_WIDTH-1:0]      s07_axi_awid,
    input  wire [ADDR_WIDTH-1:0]    s07_axi_awaddr,
    input  wire [7:0]               s07_axi_awlen,
    input  wire [2:0]               s07_axi_awsize,
    input  wire [1:0]               s07_axi_awburst,
    input  wire                     s07_axi_awlock,
    input  wire [3:0]               s07_axi_awcache,
    input  wire [2:0]               s07_axi_awprot,
    input  wire [3:0]               s07_axi_awqos,
    input  wire [AWUSER_WIDTH-1:0]  s07_axi_awuser,
    input  wire                     s07_axi_awvalid,
    output wire                     s07_axi_awready,
    input  wire [DATA_WIDTH-1:0]    s07_axi_wdata,
    input  wire [STRB_WIDTH-1:0]    s07_axi_wstrb,
    input  wire                     s07_axi_wlast,
    input  wire [WUSER_WIDTH-1:0]   s07_axi_wuser,
    input  wire                     s07_axi_wvalid,
    output wire                     s07_axi_wready,
    output wire [ID_WIDTH-1:0]      s07_axi_bid,
    output wire [1:0]               s07_axi_bresp,
    output wire [BUSER_WIDTH-1:0]   s07_axi_buser,
    output wire                     s07_axi_bvalid,
    input  wire                     s07_axi_bready,
    input  wire [ID_WIDTH-1:0]      s07_axi_arid,
    input  wire [ADDR_WIDTH-1:0]    s07_axi_araddr,
    input  wire [7:0]               s07_axi_arlen,
    input  wire [2:0]               s07_axi_arsize,
    input  wire [1:0]               s07_axi_arburst,
    input  wire                     s07_axi_arlock,
    input  wire [3:0]               s07_axi_arcache,
    input  wire [2:0]               s07_axi_arprot,
    input  wire [3:0]               s07_axi_arqos,
    input  wire [ARUSER_WIDTH-1:0]  s07_axi_aruser,
    input  wire                     s07_axi_arvalid,
    output wire                     s07_axi_arready,
    output wire [ID_WIDTH-1:0]      s07_axi_rid,
    output wire [DATA_WIDTH-1:0]    s07_axi_rdata,
    output wire [1:0]               s07_axi_rresp,
    output wire                     s07_axi_rlast,
    output wire [RUSER_WIDTH-1:0]   s07_axi_ruser,
    output wire                     s07_axi_rvalid,
    input  wire                     s07_axi_rready,

    input  wire [ID_WIDTH-1:0]      s08_axi_awid,
    input  wire [ADDR_WIDTH-1:0]    s08_axi_awaddr,
    input  wire [7:0]               s08_axi_awlen,
    input  wire [2:0]               s08_axi_awsize,
    input  wire [1:0]               s08_axi_awburst,
    input  wire                     s08_axi_awlock,
    input  wire [3:0]               s08_axi_awcache,
    input  wire [2:0]               s08_axi_awprot,
    input  wire [3:0]               s08_axi_awqos,
    input  wire [AWUSER_WIDTH-1:0]  s08_axi_awuser,
    input  wire                     s08_axi_awvalid,
    output wire                     s08_axi_awready,
    input  wire [DATA_WIDTH-1:0]    s08_axi_wdata,
    input  wire [STRB_WIDTH-1:0]    s08_axi_wstrb,
    input  wire                     s08_axi_wlast,
    input  wire [WUSER_WIDTH-1:0]   s08_axi_wuser,
    input  wire                     s08_axi_wvalid,
    output wire                     s08_axi_wready,
    output wire [ID_WIDTH-1:0]      s08_axi_bid,
    output wire [1:0]               s08_axi_bresp,
    output wire [BUSER_WIDTH-1:0]   s08_axi_buser,
    output wire                     s08_axi_bvalid,
    input  wire                     s08_axi_bready,
    input  wire [ID_WIDTH-1:0]      s08_axi_arid,
    input  wire [ADDR_WIDTH-1:0]    s08_axi_araddr,
    input  wire [7:0]               s08_axi_arlen,
    input  wire [2:0]               s08_axi_arsize,
    input  wire [1:0]               s08_axi_arburst,
    input  wire                     s08_axi_arlock,
    input  wire [3:0]               s08_axi_arcache,
    input  wire [2:0]               s08_axi_arprot,
    input  wire [3:0]               s08_axi_arqos,
    input  wire [ARUSER_WIDTH-1:0]  s08_axi_aruser,
    input  wire                     s08_axi_arvalid,
    output wire                     s08_axi_arready,
    output wire [ID_WIDTH-1:0]      s08_axi_rid,
    output wire [DATA_WIDTH-1:0]    s08_axi_rdata,
    output wire [1:0]               s08_axi_rresp,
    output wire                     s08_axi_rlast,
    output wire [RUSER_WIDTH-1:0]   s08_axi_ruser,
    output wire                     s08_axi_rvalid,
    input  wire                     s08_axi_rready,

    input  wire [ID_WIDTH-1:0]      s09_axi_awid,
    input  wire [ADDR_WIDTH-1:0]    s09_axi_awaddr,
    input  wire [7:0]               s09_axi_awlen,
    input  wire [2:0]               s09_axi_awsize,
    input  wire [1:0]               s09_axi_awburst,
    input  wire                     s09_axi_awlock,
    input  wire [3:0]               s09_axi_awcache,
    input  wire [2:0]               s09_axi_awprot,
    input  wire [3:0]               s09_axi_awqos,
    input  wire [AWUSER_WIDTH-1:0]  s09_axi_awuser,
    input  wire                     s09_axi_awvalid,
    output wire                     s09_axi_awready,
    input  wire [DATA_WIDTH-1:0]    s09_axi_wdata,
    input  wire [STRB_WIDTH-1:0]    s09_axi_wstrb,
    input  wire                     s09_axi_wlast,
    input  wire [WUSER_WIDTH-1:0]   s09_axi_wuser,
    input  wire                     s09_axi_wvalid,
    output wire                     s09_axi_wready,
    output wire [ID_WIDTH-1:0]      s09_axi_bid,
    output wire [1:0]               s09_axi_bresp,
    output wire [BUSER_WIDTH-1:0]   s09_axi_buser,
    output wire                     s09_axi_bvalid,
    input  wire                     s09_axi_bready,
    input  wire [ID_WIDTH-1:0]      s09_axi_arid,
    input  wire [ADDR_WIDTH-1:0]    s09_axi_araddr,
    input  wire [7:0]               s09_axi_arlen,
    input  wire [2:0]               s09_axi_arsize,
    input  wire [1:0]               s09_axi_arburst,
    input  wire                     s09_axi_arlock,
    input  wire [3:0]               s09_axi_arcache,
    input  wire [2:0]               s09_axi_arprot,
    input  wire [3:0]               s09_axi_arqos,
    input  wire [ARUSER_WIDTH-1:0]  s09_axi_aruser,
    input  wire                     s09_axi_arvalid,
    output wire                     s09_axi_arready,
    output wire [ID_WIDTH-1:0]      s09_axi_rid,
    output wire [DATA_WIDTH-1:0]    s09_axi_rdata,
    output wire [1:0]               s09_axi_rresp,
    output wire                     s09_axi_rlast,
    output wire [RUSER_WIDTH-1:0]   s09_axi_ruser,
    output wire                     s09_axi_rvalid,
    input  wire                     s09_axi_rready,

    input  wire [ID_WIDTH-1:0]      s10_axi_awid,
    input  wire [ADDR_WIDTH-1:0]    s10_axi_awaddr,
    input  wire [7:0]               s10_axi_awlen,
    input  wire [2:0]               s10_axi_awsize,
    input  wire [1:0]               s10_axi_awburst,
    input  wire                     s10_axi_awlock,
    input  wire [3:0]               s10_axi_awcache,
    input  wire [2:0]               s10_axi_awprot,
    input  wire [3:0]               s10_axi_awqos,
    input  wire [AWUSER_WIDTH-1:0]  s10_axi_awuser,
    input  wire                     s10_axi_awvalid,
    output wire                     s10_axi_awready,
    input  wire [DATA_WIDTH-1:0]    s10_axi_wdata,
    input  wire [STRB_WIDTH-1:0]    s10_axi_wstrb,
    input  wire                     s10_axi_wlast,
    input  wire [WUSER_WIDTH-1:0]   s10_axi_wuser,
    input  wire                     s10_axi_wvalid,
    output wire                     s10_axi_wready,
    output wire [ID_WIDTH-1:0]      s10_axi_bid,
    output wire [1:0]               s10_axi_bresp,
    output wire [BUSER_WIDTH-1:0]   s10_axi_buser,
    output wire                     s10_axi_bvalid,
    input  wire                     s10_axi_bready,
    input  wire [ID_WIDTH-1:0]      s10_axi_arid,
    input  wire [ADDR_WIDTH-1:0]    s10_axi_araddr,
    input  wire [7:0]               s10_axi_arlen,
    input  wire [2:0]               s10_axi_arsize,
    input  wire [1:0]               s10_axi_arburst,
    input  wire                     s10_axi_arlock,
    input  wire [3:0]               s10_axi_arcache,
    input  wire [2:0]               s10_axi_arprot,
    input  wire [3:0]               s10_axi_arqos,
    input  wire [ARUSER_WIDTH-1:0]  s10_axi_aruser,
    input  wire                     s10_axi_arvalid,
    output wire                     s10_axi_arready,
    output wire [ID_WIDTH-1:0]      s10_axi_rid,
    output wire [DATA_WIDTH-1:0]    s10_axi_rdata,
    output wire [1:0]               s10_axi_rresp,
    output wire                     s10_axi_rlast,
    output wire [RUSER_WIDTH-1:0]   s10_axi_ruser,
    output wire                     s10_axi_rvalid,
    input  wire                     s10_axi_rready,

    input  wire [ID_WIDTH-1:0]      s11_axi_awid,
    input  wire [ADDR_WIDTH-1:0]    s11_axi_awaddr,
    input  wire [7:0]               s11_axi_awlen,
    input  wire [2:0]               s11_axi_awsize,
    input  wire [1:0]               s11_axi_awburst,
    input  wire                     s11_axi_awlock,
    input  wire [3:0]               s11_axi_awcache,
    input  wire [2:0]               s11_axi_awprot,
    input  wire [3:0]               s11_axi_awqos,
    input  wire [AWUSER_WIDTH-1:0]  s11_axi_awuser,
    input  wire                     s11_axi_awvalid,
    output wire                     s11_axi_awready,
    input  wire [DATA_WIDTH-1:0]    s11_axi_wdata,
    input  wire [STRB_WIDTH-1:0]    s11_axi_wstrb,
    input  wire                     s11_axi_wlast,
    input  wire [WUSER_WIDTH-1:0]   s11_axi_wuser,
    input  wire                     s11_axi_wvalid,
    output wire                     s11_axi_wready,
    output wire [ID_WIDTH-1:0]      s11_axi_bid,
    output wire [1:0]               s11_axi_bresp,
    output wire [BUSER_WIDTH-1:0]   s11_axi_buser,
    output wire                     s11_axi_bvalid,
    input  wire                     s11_axi_bready,
    input  wire [ID_WIDTH-1:0]      s11_axi_arid,
    input  wire [ADDR_WIDTH-1:0]    s11_axi_araddr,
    input  wire [7:0]               s11_axi_arlen,
    input  wire [2:0]               s11_axi_arsize,
    input  wire [1:0]               s11_axi_arburst,
    input  wire                     s11_axi_arlock,
    input  wire [3:0]               s11_axi_arcache,
    input  wire [2:0]               s11_axi_arprot,
    input  wire [3:0]               s11_axi_arqos,
    input  wire [ARUSER_WIDTH-1:0]  s11_axi_aruser,
    input  wire                     s11_axi_arvalid,
    output wire                     s11_axi_arready,
    output wire [ID_WIDTH-1:0]      s11_axi_rid,
    output wire [DATA_WIDTH-1:0]    s11_axi_rdata,
    output wire [1:0]               s11_axi_rresp,
    output wire                     s11_axi_rlast,
    output wire [RUSER_WIDTH-1:0]   s11_axi_ruser,
    output wire                     s11_axi_rvalid,
    input  wire                     s11_axi_rready,

    input  wire [ID_WIDTH-1:0]      s12_axi_awid,
    input  wire [ADDR_WIDTH-1:0]    s12_axi_awaddr,
    input  wire [7:0]               s12_axi_awlen,
    input  wire [2:0]               s12_axi_awsize,
    input  wire [1:0]               s12_axi_awburst,
    input  wire                     s12_axi_awlock,
    input  wire [3:0]               s12_axi_awcache,
    input  wire [2:0]               s12_axi_awprot,
    input  wire [3:0]               s12_axi_awqos,
    input  wire [AWUSER_WIDTH-1:0]  s12_axi_awuser,
    input  wire                     s12_axi_awvalid,
    output wire                     s12_axi_awready,
    input  wire [DATA_WIDTH-1:0]    s12_axi_wdata,
    input  wire [STRB_WIDTH-1:0]    s12_axi_wstrb,
    input  wire                     s12_axi_wlast,
    input  wire [WUSER_WIDTH-1:0]   s12_axi_wuser,
    input  wire                     s12_axi_wvalid,
    output wire                     s12_axi_wready,
    output wire [ID_WIDTH-1:0]      s12_axi_bid,
    output wire [1:0]               s12_axi_bresp,
    output wire [BUSER_WIDTH-1:0]   s12_axi_buser,
    output wire                     s12_axi_bvalid,
    input  wire                     s12_axi_bready,
    input  wire [ID_WIDTH-1:0]      s12_axi_arid,
    input  wire [ADDR_WIDTH-1:0]    s12_axi_araddr,
    input  wire [7:0]               s12_axi_arlen,
    input  wire [2:0]               s12_axi_arsize,
    input  wire [1:0]               s12_axi_arburst,
    input  wire                     s12_axi_arlock,
    input  wire [3:0]               s12_axi_arcache,
    input  wire [2:0]               s12_axi_arprot,
    input  wire [3:0]               s12_axi_arqos,
    input  wire [ARUSER_WIDTH-1:0]  s12_axi_aruser,
    input  wire                     s12_axi_arvalid,
    output wire                     s12_axi_arready,
    output wire [ID_WIDTH-1:0]      s12_axi_rid,
    output wire [DATA_WIDTH-1:0]    s12_axi_rdata,
    output wire [1:0]               s12_axi_rresp,
    output wire                     s12_axi_rlast,
    output wire [RUSER_WIDTH-1:0]   s12_axi_ruser,
    output wire                     s12_axi_rvalid,
    input  wire                     s12_axi_rready,

    input  wire [ID_WIDTH-1:0]      s13_axi_awid,
    input  wire [ADDR_WIDTH-1:0]    s13_axi_awaddr,
    input  wire [7:0]               s13_axi_awlen,
    input  wire [2:0]               s13_axi_awsize,
    input  wire [1:0]               s13_axi_awburst,
    input  wire                     s13_axi_awlock,
    input  wire [3:0]               s13_axi_awcache,
    input  wire [2:0]               s13_axi_awprot,
    input  wire [3:0]               s13_axi_awqos,
    input  wire [AWUSER_WIDTH-1:0]  s13_axi_awuser,
    input  wire                     s13_axi_awvalid,
    output wire                     s13_axi_awready,
    input  wire [DATA_WIDTH-1:0]    s13_axi_wdata,
    input  wire [STRB_WIDTH-1:0]    s13_axi_wstrb,
    input  wire                     s13_axi_wlast,
    input  wire [WUSER_WIDTH-1:0]   s13_axi_wuser,
    input  wire                     s13_axi_wvalid,
    output wire                     s13_axi_wready,
    output wire [ID_WIDTH-1:0]      s13_axi_bid,
    output wire [1:0]               s13_axi_bresp,
    output wire [BUSER_WIDTH-1:0]   s13_axi_buser,
    output wire                     s13_axi_bvalid,
    input  wire                     s13_axi_bready,
    input  wire [ID_WIDTH-1:0]      s13_axi_arid,
    input  wire [ADDR_WIDTH-1:0]    s13_axi_araddr,
    input  wire [7:0]               s13_axi_arlen,
    input  wire [2:0]               s13_axi_arsize,
    input  wire [1:0]               s13_axi_arburst,
    input  wire                     s13_axi_arlock,
    input  wire [3:0]               s13_axi_arcache,
    input  wire [2:0]               s13_axi_arprot,
    input  wire [3:0]               s13_axi_arqos,
    input  wire [ARUSER_WIDTH-1:0]  s13_axi_aruser,
    input  wire                     s13_axi_arvalid,
    output wire                     s13_axi_arready,
    output wire [ID_WIDTH-1:0]      s13_axi_rid,
    output wire [DATA_WIDTH-1:0]    s13_axi_rdata,
    output wire [1:0]               s13_axi_rresp,
    output wire                     s13_axi_rlast,
    output wire [RUSER_WIDTH-1:0]   s13_axi_ruser,
    output wire                     s13_axi_rvalid,
    input  wire                     s13_axi_rready,

    input  wire [ID_WIDTH-1:0]      s14_axi_awid,
    input  wire [ADDR_WIDTH-1:0]    s14_axi_awaddr,
    input  wire [7:0]               s14_axi_awlen,
    input  wire [2:0]               s14_axi_awsize,
    input  wire [1:0]               s14_axi_awburst,
    input  wire                     s14_axi_awlock,
    input  wire [3:0]               s14_axi_awcache,
    input  wire [2:0]               s14_axi_awprot,
    input  wire [3:0]               s14_axi_awqos,
    input  wire [AWUSER_WIDTH-1:0]  s14_axi_awuser,
    input  wire                     s14_axi_awvalid,
    output wire                     s14_axi_awready,
    input  wire [DATA_WIDTH-1:0]    s14_axi_wdata,
    input  wire [STRB_WIDTH-1:0]    s14_axi_wstrb,
    input  wire                     s14_axi_wlast,
    input  wire [WUSER_WIDTH-1:0]   s14_axi_wuser,
    input  wire                     s14_axi_wvalid,
    output wire                     s14_axi_wready,
    output wire [ID_WIDTH-1:0]      s14_axi_bid,
    output wire [1:0]               s14_axi_bresp,
    output wire [BUSER_WIDTH-1:0]   s14_axi_buser,
    output wire                     s14_axi_bvalid,
    input  wire                     s14_axi_bready,
    input  wire [ID_WIDTH-1:0]      s14_axi_arid,
    input  wire [ADDR_WIDTH-1:0]    s14_axi_araddr,
    input  wire [7:0]               s14_axi_arlen,
    input  wire [2:0]               s14_axi_arsize,
    input  wire [1:0]               s14_axi_arburst,
    input  wire                     s14_axi_arlock,
    input  wire [3:0]               s14_axi_arcache,
    input  wire [2:0]               s14_axi_arprot,
    input  wire [3:0]               s14_axi_arqos,
    input  wire [ARUSER_WIDTH-1:0]  s14_axi_aruser,
    input  wire                     s14_axi_arvalid,
    output wire                     s14_axi_arready,
    output wire [ID_WIDTH-1:0]      s14_axi_rid,
    output wire [DATA_WIDTH-1:0]    s14_axi_rdata,
    output wire [1:0]               s14_axi_rresp,
    output wire                     s14_axi_rlast,
    output wire [RUSER_WIDTH-1:0]   s14_axi_ruser,
    output wire                     s14_axi_rvalid,
    input  wire                     s14_axi_rready,

    input  wire [ID_WIDTH-1:0]      s15_axi_awid,
    input  wire [ADDR_WIDTH-1:0]    s15_axi_awaddr,
    input  wire [7:0]               s15_axi_awlen,
    input  wire [2:0]               s15_axi_awsize,
    input  wire [1:0]               s15_axi_awburst,
    input  wire                     s15_axi_awlock,
    input  wire [3:0]               s15_axi_awcache,
    input  wire [2:0]               s15_axi_awprot,
    input  wire [3:0]               s15_axi_awqos,
    input  wire [AWUSER_WIDTH-1:0]  s15_axi_awuser,
    input  wire                     s15_axi_awvalid,
    output wire                     s15_axi_awready,
    input  wire [DATA_WIDTH-1:0]    s15_axi_wdata,
    input  wire [STRB_WIDTH-1:0]    s15_axi_wstrb,
    input  wire                     s15_axi_wlast,
    input  wire [WUSER_WIDTH-1:0]   s15_axi_wuser,
    input  wire                     s15_axi_wvalid,
    output wire                     s15_axi_wready,
    output wire [ID_WIDTH-1:0]      s15_axi_bid,
    output wire [1:0]               s15_axi_bresp,
    output wire [BUSER_WIDTH-1:0]   s15_axi_buser,
    output wire                     s15_axi_bvalid,
    input  wire                     s15_axi_bready,
    input  wire [ID_WIDTH-1:0]      s15_axi_arid,
    input  wire [ADDR_WIDTH-1:0]    s15_axi_araddr,
    input  wire [7:0]               s15_axi_arlen,
    input  wire [2:0]               s15_axi_arsize,
    input  wire [1:0]               s15_axi_arburst,
    input  wire                     s15_axi_arlock,
    input  wire [3:0]               s15_axi_arcache,
    input  wire [2:0]               s15_axi_arprot,
    input  wire [3:0]               s15_axi_arqos,
    input  wire [ARUSER_WIDTH-1:0]  s15_axi_aruser,
    input  wire                     s15_axi_arvalid,
    output wire                     s15_axi_arready,
    output wire [ID_WIDTH-1:0]      s15_axi_rid,
    output wire [DATA_WIDTH-1:0]    s15_axi_rdata,
    output wire [1:0]               s15_axi_rresp,
    output wire                     s15_axi_rlast,
    output wire [RUSER_WIDTH-1:0]   s15_axi_ruser,
    output wire                     s15_axi_rvalid,
    input  wire                     s15_axi_rready,

    input  wire [ID_WIDTH-1:0]      s16_axi_awid,
    input  wire [ADDR_WIDTH-1:0]    s16_axi_awaddr,
    input  wire [7:0]               s16_axi_awlen,
    input  wire [2:0]               s16_axi_awsize,
    input  wire [1:0]               s16_axi_awburst,
    input  wire                     s16_axi_awlock,
    input  wire [3:0]               s16_axi_awcache,
    input  wire [2:0]               s16_axi_awprot,
    input  wire [3:0]               s16_axi_awqos,
    input  wire [AWUSER_WIDTH-1:0]  s16_axi_awuser,
    input  wire                     s16_axi_awvalid,
    output wire                     s16_axi_awready,
    input  wire [DATA_WIDTH-1:0]    s16_axi_wdata,
    input  wire [STRB_WIDTH-1:0]    s16_axi_wstrb,
    input  wire                     s16_axi_wlast,
    input  wire [WUSER_WIDTH-1:0]   s16_axi_wuser,
    input  wire                     s16_axi_wvalid,
    output wire                     s16_axi_wready,
    output wire [ID_WIDTH-1:0]      s16_axi_bid,
    output wire [1:0]               s16_axi_bresp,
    output wire [BUSER_WIDTH-1:0]   s16_axi_buser,
    output wire                     s16_axi_bvalid,
    input  wire                     s16_axi_bready,
    input  wire [ID_WIDTH-1:0]      s16_axi_arid,
    input  wire [ADDR_WIDTH-1:0]    s16_axi_araddr,
    input  wire [7:0]               s16_axi_arlen,
    input  wire [2:0]               s16_axi_arsize,
    input  wire [1:0]               s16_axi_arburst,
    input  wire                     s16_axi_arlock,
    input  wire [3:0]               s16_axi_arcache,
    input  wire [2:0]               s16_axi_arprot,
    input  wire [3:0]               s16_axi_arqos,
    input  wire [ARUSER_WIDTH-1:0]  s16_axi_aruser,
    input  wire                     s16_axi_arvalid,
    output wire                     s16_axi_arready,
    output wire [ID_WIDTH-1:0]      s16_axi_rid,
    output wire [DATA_WIDTH-1:0]    s16_axi_rdata,
    output wire [1:0]               s16_axi_rresp,
    output wire                     s16_axi_rlast,
    output wire [RUSER_WIDTH-1:0]   s16_axi_ruser,
    output wire                     s16_axi_rvalid,
    input  wire                     s16_axi_rready,

    input  wire [ID_WIDTH-1:0]      s17_axi_awid,
    input  wire [ADDR_WIDTH-1:0]    s17_axi_awaddr,
    input  wire [7:0]               s17_axi_awlen,
    input  wire [2:0]               s17_axi_awsize,
    input  wire [1:0]               s17_axi_awburst,
    input  wire                     s17_axi_awlock,
    input  wire [3:0]               s17_axi_awcache,
    input  wire [2:0]               s17_axi_awprot,
    input  wire [3:0]               s17_axi_awqos,
    input  wire [AWUSER_WIDTH-1:0]  s17_axi_awuser,
    input  wire                     s17_axi_awvalid,
    output wire                     s17_axi_awready,
    input  wire [DATA_WIDTH-1:0]    s17_axi_wdata,
    input  wire [STRB_WIDTH-1:0]    s17_axi_wstrb,
    input  wire                     s17_axi_wlast,
    input  wire [WUSER_WIDTH-1:0]   s17_axi_wuser,
    input  wire                     s17_axi_wvalid,
    output wire                     s17_axi_wready,
    output wire [ID_WIDTH-1:0]      s17_axi_bid,
    output wire [1:0]               s17_axi_bresp,
    output wire [BUSER_WIDTH-1:0]   s17_axi_buser,
    output wire                     s17_axi_bvalid,
    input  wire                     s17_axi_bready,
    input  wire [ID_WIDTH-1:0]      s17_axi_arid,
    input  wire [ADDR_WIDTH-1:0]    s17_axi_araddr,
    input  wire [7:0]               s17_axi_arlen,
    input  wire [2:0]               s17_axi_arsize,
    input  wire [1:0]               s17_axi_arburst,
    input  wire                     s17_axi_arlock,
    input  wire [3:0]               s17_axi_arcache,
    input  wire [2:0]               s17_axi_arprot,
    input  wire [3:0]               s17_axi_arqos,
    input  wire [ARUSER_WIDTH-1:0]  s17_axi_aruser,
    input  wire                     s17_axi_arvalid,
    output wire                     s17_axi_arready,
    output wire [ID_WIDTH-1:0]      s17_axi_rid,
    output wire [DATA_WIDTH-1:0]    s17_axi_rdata,
    output wire [1:0]               s17_axi_rresp,
    output wire                     s17_axi_rlast,
    output wire [RUSER_WIDTH-1:0]   s17_axi_ruser,
    output wire                     s17_axi_rvalid,
    input  wire                     s17_axi_rready,

    input  wire [ID_WIDTH-1:0]      s18_axi_awid,
    input  wire [ADDR_WIDTH-1:0]    s18_axi_awaddr,
    input  wire [7:0]               s18_axi_awlen,
    input  wire [2:0]               s18_axi_awsize,
    input  wire [1:0]               s18_axi_awburst,
    input  wire                     s18_axi_awlock,
    input  wire [3:0]               s18_axi_awcache,
    input  wire [2:0]               s18_axi_awprot,
    input  wire [3:0]               s18_axi_awqos,
    input  wire [AWUSER_WIDTH-1:0]  s18_axi_awuser,
    input  wire                     s18_axi_awvalid,
    output wire                     s18_axi_awready,
    input  wire [DATA_WIDTH-1:0]    s18_axi_wdata,
    input  wire [STRB_WIDTH-1:0]    s18_axi_wstrb,
    input  wire                     s18_axi_wlast,
    input  wire [WUSER_WIDTH-1:0]   s18_axi_wuser,
    input  wire                     s18_axi_wvalid,
    output wire                     s18_axi_wready,
    output wire [ID_WIDTH-1:0]      s18_axi_bid,
    output wire [1:0]               s18_axi_bresp,
    output wire [BUSER_WIDTH-1:0]   s18_axi_buser,
    output wire                     s18_axi_bvalid,
    input  wire                     s18_axi_bready,
    input  wire [ID_WIDTH-1:0]      s18_axi_arid,
    input  wire [ADDR_WIDTH-1:0]    s18_axi_araddr,
    input  wire [7:0]               s18_axi_arlen,
    input  wire [2:0]               s18_axi_arsize,
    input  wire [1:0]               s18_axi_arburst,
    input  wire                     s18_axi_arlock,
    input  wire [3:0]               s18_axi_arcache,
    input  wire [2:0]               s18_axi_arprot,
    input  wire [3:0]               s18_axi_arqos,
    input  wire [ARUSER_WIDTH-1:0]  s18_axi_aruser,
    input  wire                     s18_axi_arvalid,
    output wire                     s18_axi_arready,
    output wire [ID_WIDTH-1:0]      s18_axi_rid,
    output wire [DATA_WIDTH-1:0]    s18_axi_rdata,
    output wire [1:0]               s18_axi_rresp,
    output wire                     s18_axi_rlast,
    output wire [RUSER_WIDTH-1:0]   s18_axi_ruser,
    output wire                     s18_axi_rvalid,
    input  wire                     s18_axi_rready,

    input  wire [ID_WIDTH-1:0]      s19_axi_awid,
    input  wire [ADDR_WIDTH-1:0]    s19_axi_awaddr,
    input  wire [7:0]               s19_axi_awlen,
    input  wire [2:0]               s19_axi_awsize,
    input  wire [1:0]               s19_axi_awburst,
    input  wire                     s19_axi_awlock,
    input  wire [3:0]               s19_axi_awcache,
    input  wire [2:0]               s19_axi_awprot,
    input  wire [3:0]               s19_axi_awqos,
    input  wire [AWUSER_WIDTH-1:0]  s19_axi_awuser,
    input  wire                     s19_axi_awvalid,
    output wire                     s19_axi_awready,
    input  wire [DATA_WIDTH-1:0]    s19_axi_wdata,
    input  wire [STRB_WIDTH-1:0]    s19_axi_wstrb,
    input  wire                     s19_axi_wlast,
    input  wire [WUSER_WIDTH-1:0]   s19_axi_wuser,
    input  wire                     s19_axi_wvalid,
    output wire                     s19_axi_wready,
    output wire [ID_WIDTH-1:0]      s19_axi_bid,
    output wire [1:0]               s19_axi_bresp,
    output wire [BUSER_WIDTH-1:0]   s19_axi_buser,
    output wire                     s19_axi_bvalid,
    input  wire                     s19_axi_bready,
    input  wire [ID_WIDTH-1:0]      s19_axi_arid,
    input  wire [ADDR_WIDTH-1:0]    s19_axi_araddr,
    input  wire [7:0]               s19_axi_arlen,
    input  wire [2:0]               s19_axi_arsize,
    input  wire [1:0]               s19_axi_arburst,
    input  wire                     s19_axi_arlock,
    input  wire [3:0]               s19_axi_arcache,
    input  wire [2:0]               s19_axi_arprot,
    input  wire [3:0]               s19_axi_arqos,
    input  wire [ARUSER_WIDTH-1:0]  s19_axi_aruser,
    input  wire                     s19_axi_arvalid,
    output wire                     s19_axi_arready,
    output wire [ID_WIDTH-1:0]      s19_axi_rid,
    output wire [DATA_WIDTH-1:0]    s19_axi_rdata,
    output wire [1:0]               s19_axi_rresp,
    output wire                     s19_axi_rlast,
    output wire [RUSER_WIDTH-1:0]   s19_axi_ruser,
    output wire                     s19_axi_rvalid,
    input  wire                     s19_axi_rready,

    input  wire [ID_WIDTH-1:0]      s20_axi_awid,
    input  wire [ADDR_WIDTH-1:0]    s20_axi_awaddr,
    input  wire [7:0]               s20_axi_awlen,
    input  wire [2:0]               s20_axi_awsize,
    input  wire [1:0]               s20_axi_awburst,
    input  wire                     s20_axi_awlock,
    input  wire [3:0]               s20_axi_awcache,
    input  wire [2:0]               s20_axi_awprot,
    input  wire [3:0]               s20_axi_awqos,
    input  wire [AWUSER_WIDTH-1:0]  s20_axi_awuser,
    input  wire                     s20_axi_awvalid,
    output wire                     s20_axi_awready,
    input  wire [DATA_WIDTH-1:0]    s20_axi_wdata,
    input  wire [STRB_WIDTH-1:0]    s20_axi_wstrb,
    input  wire                     s20_axi_wlast,
    input  wire [WUSER_WIDTH-1:0]   s20_axi_wuser,
    input  wire                     s20_axi_wvalid,
    output wire                     s20_axi_wready,
    output wire [ID_WIDTH-1:0]      s20_axi_bid,
    output wire [1:0]               s20_axi_bresp,
    output wire [BUSER_WIDTH-1:0]   s20_axi_buser,
    output wire                     s20_axi_bvalid,
    input  wire                     s20_axi_bready,
    input  wire [ID_WIDTH-1:0]      s20_axi_arid,
    input  wire [ADDR_WIDTH-1:0]    s20_axi_araddr,
    input  wire [7:0]               s20_axi_arlen,
    input  wire [2:0]               s20_axi_arsize,
    input  wire [1:0]               s20_axi_arburst,
    input  wire                     s20_axi_arlock,
    input  wire [3:0]               s20_axi_arcache,
    input  wire [2:0]               s20_axi_arprot,
    input  wire [3:0]               s20_axi_arqos,
    input  wire [ARUSER_WIDTH-1:0]  s20_axi_aruser,
    input  wire                     s20_axi_arvalid,
    output wire                     s20_axi_arready,
    output wire [ID_WIDTH-1:0]      s20_axi_rid,
    output wire [DATA_WIDTH-1:0]    s20_axi_rdata,
    output wire [1:0]               s20_axi_rresp,
    output wire                     s20_axi_rlast,
    output wire [RUSER_WIDTH-1:0]   s20_axi_ruser,
    output wire                     s20_axi_rvalid,
    input  wire                     s20_axi_rready,

    input  wire [ID_WIDTH-1:0]      s21_axi_awid,
    input  wire [ADDR_WIDTH-1:0]    s21_axi_awaddr,
    input  wire [7:0]               s21_axi_awlen,
    input  wire [2:0]               s21_axi_awsize,
    input  wire [1:0]               s21_axi_awburst,
    input  wire                     s21_axi_awlock,
    input  wire [3:0]               s21_axi_awcache,
    input  wire [2:0]               s21_axi_awprot,
    input  wire [3:0]               s21_axi_awqos,
    input  wire [AWUSER_WIDTH-1:0]  s21_axi_awuser,
    input  wire                     s21_axi_awvalid,
    output wire                     s21_axi_awready,
    input  wire [DATA_WIDTH-1:0]    s21_axi_wdata,
    input  wire [STRB_WIDTH-1:0]    s21_axi_wstrb,
    input  wire                     s21_axi_wlast,
    input  wire [WUSER_WIDTH-1:0]   s21_axi_wuser,
    input  wire                     s21_axi_wvalid,
    output wire                     s21_axi_wready,
    output wire [ID_WIDTH-1:0]      s21_axi_bid,
    output wire [1:0]               s21_axi_bresp,
    output wire [BUSER_WIDTH-1:0]   s21_axi_buser,
    output wire                     s21_axi_bvalid,
    input  wire                     s21_axi_bready,
    input  wire [ID_WIDTH-1:0]      s21_axi_arid,
    input  wire [ADDR_WIDTH-1:0]    s21_axi_araddr,
    input  wire [7:0]               s21_axi_arlen,
    input  wire [2:0]               s21_axi_arsize,
    input  wire [1:0]               s21_axi_arburst,
    input  wire                     s21_axi_arlock,
    input  wire [3:0]               s21_axi_arcache,
    input  wire [2:0]               s21_axi_arprot,
    input  wire [3:0]               s21_axi_arqos,
    input  wire [ARUSER_WIDTH-1:0]  s21_axi_aruser,
    input  wire                     s21_axi_arvalid,
    output wire                     s21_axi_arready,
    output wire [ID_WIDTH-1:0]      s21_axi_rid,
    output wire [DATA_WIDTH-1:0]    s21_axi_rdata,
    output wire [1:0]               s21_axi_rresp,
    output wire                     s21_axi_rlast,
    output wire [RUSER_WIDTH-1:0]   s21_axi_ruser,
    output wire                     s21_axi_rvalid,
    input  wire                     s21_axi_rready,

    input  wire [ID_WIDTH-1:0]      s22_axi_awid,
    input  wire [ADDR_WIDTH-1:0]    s22_axi_awaddr,
    input  wire [7:0]               s22_axi_awlen,
    input  wire [2:0]               s22_axi_awsize,
    input  wire [1:0]               s22_axi_awburst,
    input  wire                     s22_axi_awlock,
    input  wire [3:0]               s22_axi_awcache,
    input  wire [2:0]               s22_axi_awprot,
    input  wire [3:0]               s22_axi_awqos,
    input  wire [AWUSER_WIDTH-1:0]  s22_axi_awuser,
    input  wire                     s22_axi_awvalid,
    output wire                     s22_axi_awready,
    input  wire [DATA_WIDTH-1:0]    s22_axi_wdata,
    input  wire [STRB_WIDTH-1:0]    s22_axi_wstrb,
    input  wire                     s22_axi_wlast,
    input  wire [WUSER_WIDTH-1:0]   s22_axi_wuser,
    input  wire                     s22_axi_wvalid,
    output wire                     s22_axi_wready,
    output wire [ID_WIDTH-1:0]      s22_axi_bid,
    output wire [1:0]               s22_axi_bresp,
    output wire [BUSER_WIDTH-1:0]   s22_axi_buser,
    output wire                     s22_axi_bvalid,
    input  wire                     s22_axi_bready,
    input  wire [ID_WIDTH-1:0]      s22_axi_arid,
    input  wire [ADDR_WIDTH-1:0]    s22_axi_araddr,
    input  wire [7:0]               s22_axi_arlen,
    input  wire [2:0]               s22_axi_arsize,
    input  wire [1:0]               s22_axi_arburst,
    input  wire                     s22_axi_arlock,
    input  wire [3:0]               s22_axi_arcache,
    input  wire [2:0]               s22_axi_arprot,
    input  wire [3:0]               s22_axi_arqos,
    input  wire [ARUSER_WIDTH-1:0]  s22_axi_aruser,
    input  wire                     s22_axi_arvalid,
    output wire                     s22_axi_arready,
    output wire [ID_WIDTH-1:0]      s22_axi_rid,
    output wire [DATA_WIDTH-1:0]    s22_axi_rdata,
    output wire [1:0]               s22_axi_rresp,
    output wire                     s22_axi_rlast,
    output wire [RUSER_WIDTH-1:0]   s22_axi_ruser,
    output wire                     s22_axi_rvalid,
    input  wire                     s22_axi_rready,

    input  wire [ID_WIDTH-1:0]      s23_axi_awid,
    input  wire [ADDR_WIDTH-1:0]    s23_axi_awaddr,
    input  wire [7:0]               s23_axi_awlen,
    input  wire [2:0]               s23_axi_awsize,
    input  wire [1:0]               s23_axi_awburst,
    input  wire                     s23_axi_awlock,
    input  wire [3:0]               s23_axi_awcache,
    input  wire [2:0]               s23_axi_awprot,
    input  wire [3:0]               s23_axi_awqos,
    input  wire [AWUSER_WIDTH-1:0]  s23_axi_awuser,
    input  wire                     s23_axi_awvalid,
    output wire                     s23_axi_awready,
    input  wire [DATA_WIDTH-1:0]    s23_axi_wdata,
    input  wire [STRB_WIDTH-1:0]    s23_axi_wstrb,
    input  wire                     s23_axi_wlast,
    input  wire [WUSER_WIDTH-1:0]   s23_axi_wuser,
    input  wire                     s23_axi_wvalid,
    output wire                     s23_axi_wready,
    output wire [ID_WIDTH-1:0]      s23_axi_bid,
    output wire [1:0]               s23_axi_bresp,
    output wire [BUSER_WIDTH-1:0]   s23_axi_buser,
    output wire                     s23_axi_bvalid,
    input  wire                     s23_axi_bready,
    input  wire [ID_WIDTH-1:0]      s23_axi_arid,
    input  wire [ADDR_WIDTH-1:0]    s23_axi_araddr,
    input  wire [7:0]               s23_axi_arlen,
    input  wire [2:0]               s23_axi_arsize,
    input  wire [1:0]               s23_axi_arburst,
    input  wire                     s23_axi_arlock,
    input  wire [3:0]               s23_axi_arcache,
    input  wire [2:0]               s23_axi_arprot,
    input  wire [3:0]               s23_axi_arqos,
    input  wire [ARUSER_WIDTH-1:0]  s23_axi_aruser,
    input  wire                     s23_axi_arvalid,
    output wire                     s23_axi_arready,
    output wire [ID_WIDTH-1:0]      s23_axi_rid,
    output wire [DATA_WIDTH-1:0]    s23_axi_rdata,
    output wire [1:0]               s23_axi_rresp,
    output wire                     s23_axi_rlast,
    output wire [RUSER_WIDTH-1:0]   s23_axi_ruser,
    output wire                     s23_axi_rvalid,
    input  wire                     s23_axi_rready,

    input  wire [ID_WIDTH-1:0]      s24_axi_awid,
    input  wire [ADDR_WIDTH-1:0]    s24_axi_awaddr,
    input  wire [7:0]               s24_axi_awlen,
    input  wire [2:0]               s24_axi_awsize,
    input  wire [1:0]               s24_axi_awburst,
    input  wire                     s24_axi_awlock,
    input  wire [3:0]               s24_axi_awcache,
    input  wire [2:0]               s24_axi_awprot,
    input  wire [3:0]               s24_axi_awqos,
    input  wire [AWUSER_WIDTH-1:0]  s24_axi_awuser,
    input  wire                     s24_axi_awvalid,
    output wire                     s24_axi_awready,
    input  wire [DATA_WIDTH-1:0]    s24_axi_wdata,
    input  wire [STRB_WIDTH-1:0]    s24_axi_wstrb,
    input  wire                     s24_axi_wlast,
    input  wire [WUSER_WIDTH-1:0]   s24_axi_wuser,
    input  wire                     s24_axi_wvalid,
    output wire                     s24_axi_wready,
    output wire [ID_WIDTH-1:0]      s24_axi_bid,
    output wire [1:0]               s24_axi_bresp,
    output wire [BUSER_WIDTH-1:0]   s24_axi_buser,
    output wire                     s24_axi_bvalid,
    input  wire                     s24_axi_bready,
    input  wire [ID_WIDTH-1:0]      s24_axi_arid,
    input  wire [ADDR_WIDTH-1:0]    s24_axi_araddr,
    input  wire [7:0]               s24_axi_arlen,
    input  wire [2:0]               s24_axi_arsize,
    input  wire [1:0]               s24_axi_arburst,
    input  wire                     s24_axi_arlock,
    input  wire [3:0]               s24_axi_arcache,
    input  wire [2:0]               s24_axi_arprot,
    input  wire [3:0]               s24_axi_arqos,
    input  wire [ARUSER_WIDTH-1:0]  s24_axi_aruser,
    input  wire                     s24_axi_arvalid,
    output wire                     s24_axi_arready,
    output wire [ID_WIDTH-1:0]      s24_axi_rid,
    output wire [DATA_WIDTH-1:0]    s24_axi_rdata,
    output wire [1:0]               s24_axi_rresp,
    output wire                     s24_axi_rlast,
    output wire [RUSER_WIDTH-1:0]   s24_axi_ruser,
    output wire                     s24_axi_rvalid,
    input  wire                     s24_axi_rready,

    input  wire [ID_WIDTH-1:0]      s25_axi_awid,
    input  wire [ADDR_WIDTH-1:0]    s25_axi_awaddr,
    input  wire [7:0]               s25_axi_awlen,
    input  wire [2:0]               s25_axi_awsize,
    input  wire [1:0]               s25_axi_awburst,
    input  wire                     s25_axi_awlock,
    input  wire [3:0]               s25_axi_awcache,
    input  wire [2:0]               s25_axi_awprot,
    input  wire [3:0]               s25_axi_awqos,
    input  wire [AWUSER_WIDTH-1:0]  s25_axi_awuser,
    input  wire                     s25_axi_awvalid,
    output wire                     s25_axi_awready,
    input  wire [DATA_WIDTH-1:0]    s25_axi_wdata,
    input  wire [STRB_WIDTH-1:0]    s25_axi_wstrb,
    input  wire                     s25_axi_wlast,
    input  wire [WUSER_WIDTH-1:0]   s25_axi_wuser,
    input  wire                     s25_axi_wvalid,
    output wire                     s25_axi_wready,
    output wire [ID_WIDTH-1:0]      s25_axi_bid,
    output wire [1:0]               s25_axi_bresp,
    output wire [BUSER_WIDTH-1:0]   s25_axi_buser,
    output wire                     s25_axi_bvalid,
    input  wire                     s25_axi_bready,
    input  wire [ID_WIDTH-1:0]      s25_axi_arid,
    input  wire [ADDR_WIDTH-1:0]    s25_axi_araddr,
    input  wire [7:0]               s25_axi_arlen,
    input  wire [2:0]               s25_axi_arsize,
    input  wire [1:0]               s25_axi_arburst,
    input  wire                     s25_axi_arlock,
    input  wire [3:0]               s25_axi_arcache,
    input  wire [2:0]               s25_axi_arprot,
    input  wire [3:0]               s25_axi_arqos,
    input  wire [ARUSER_WIDTH-1:0]  s25_axi_aruser,
    input  wire                     s25_axi_arvalid,
    output wire                     s25_axi_arready,
    output wire [ID_WIDTH-1:0]      s25_axi_rid,
    output wire [DATA_WIDTH-1:0]    s25_axi_rdata,
    output wire [1:0]               s25_axi_rresp,
    output wire                     s25_axi_rlast,
    output wire [RUSER_WIDTH-1:0]   s25_axi_ruser,
    output wire                     s25_axi_rvalid,
    input  wire                     s25_axi_rready,

    input  wire [ID_WIDTH-1:0]      s26_axi_awid,
    input  wire [ADDR_WIDTH-1:0]    s26_axi_awaddr,
    input  wire [7:0]               s26_axi_awlen,
    input  wire [2:0]               s26_axi_awsize,
    input  wire [1:0]               s26_axi_awburst,
    input  wire                     s26_axi_awlock,
    input  wire [3:0]               s26_axi_awcache,
    input  wire [2:0]               s26_axi_awprot,
    input  wire [3:0]               s26_axi_awqos,
    input  wire [AWUSER_WIDTH-1:0]  s26_axi_awuser,
    input  wire                     s26_axi_awvalid,
    output wire                     s26_axi_awready,
    input  wire [DATA_WIDTH-1:0]    s26_axi_wdata,
    input  wire [STRB_WIDTH-1:0]    s26_axi_wstrb,
    input  wire                     s26_axi_wlast,
    input  wire [WUSER_WIDTH-1:0]   s26_axi_wuser,
    input  wire                     s26_axi_wvalid,
    output wire                     s26_axi_wready,
    output wire [ID_WIDTH-1:0]      s26_axi_bid,
    output wire [1:0]               s26_axi_bresp,
    output wire [BUSER_WIDTH-1:0]   s26_axi_buser,
    output wire                     s26_axi_bvalid,
    input  wire                     s26_axi_bready,
    input  wire [ID_WIDTH-1:0]      s26_axi_arid,
    input  wire [ADDR_WIDTH-1:0]    s26_axi_araddr,
    input  wire [7:0]               s26_axi_arlen,
    input  wire [2:0]               s26_axi_arsize,
    input  wire [1:0]               s26_axi_arburst,
    input  wire                     s26_axi_arlock,
    input  wire [3:0]               s26_axi_arcache,
    input  wire [2:0]               s26_axi_arprot,
    input  wire [3:0]               s26_axi_arqos,
    input  wire [ARUSER_WIDTH-1:0]  s26_axi_aruser,
    input  wire                     s26_axi_arvalid,
    output wire                     s26_axi_arready,
    output wire [ID_WIDTH-1:0]      s26_axi_rid,
    output wire [DATA_WIDTH-1:0]    s26_axi_rdata,
    output wire [1:0]               s26_axi_rresp,
    output wire                     s26_axi_rlast,
    output wire [RUSER_WIDTH-1:0]   s26_axi_ruser,
    output wire                     s26_axi_rvalid,
    input  wire                     s26_axi_rready,

    input  wire [ID_WIDTH-1:0]      s27_axi_awid,
    input  wire [ADDR_WIDTH-1:0]    s27_axi_awaddr,
    input  wire [7:0]               s27_axi_awlen,
    input  wire [2:0]               s27_axi_awsize,
    input  wire [1:0]               s27_axi_awburst,
    input  wire                     s27_axi_awlock,
    input  wire [3:0]               s27_axi_awcache,
    input  wire [2:0]               s27_axi_awprot,
    input  wire [3:0]               s27_axi_awqos,
    input  wire [AWUSER_WIDTH-1:0]  s27_axi_awuser,
    input  wire                     s27_axi_awvalid,
    output wire                     s27_axi_awready,
    input  wire [DATA_WIDTH-1:0]    s27_axi_wdata,
    input  wire [STRB_WIDTH-1:0]    s27_axi_wstrb,
    input  wire                     s27_axi_wlast,
    input  wire [WUSER_WIDTH-1:0]   s27_axi_wuser,
    input  wire                     s27_axi_wvalid,
    output wire                     s27_axi_wready,
    output wire [ID_WIDTH-1:0]      s27_axi_bid,
    output wire [1:0]               s27_axi_bresp,
    output wire [BUSER_WIDTH-1:0]   s27_axi_buser,
    output wire                     s27_axi_bvalid,
    input  wire                     s27_axi_bready,
    input  wire [ID_WIDTH-1:0]      s27_axi_arid,
    input  wire [ADDR_WIDTH-1:0]    s27_axi_araddr,
    input  wire [7:0]               s27_axi_arlen,
    input  wire [2:0]               s27_axi_arsize,
    input  wire [1:0]               s27_axi_arburst,
    input  wire                     s27_axi_arlock,
    input  wire [3:0]               s27_axi_arcache,
    input  wire [2:0]               s27_axi_arprot,
    input  wire [3:0]               s27_axi_arqos,
    input  wire [ARUSER_WIDTH-1:0]  s27_axi_aruser,
    input  wire                     s27_axi_arvalid,
    output wire                     s27_axi_arready,
    output wire [ID_WIDTH-1:0]      s27_axi_rid,
    output wire [DATA_WIDTH-1:0]    s27_axi_rdata,
    output wire [1:0]               s27_axi_rresp,
    output wire                     s27_axi_rlast,
    output wire [RUSER_WIDTH-1:0]   s27_axi_ruser,
    output wire                     s27_axi_rvalid,
    input  wire                     s27_axi_rready,

    /*
     * AXI master interface
     */
    output wire [ID_WIDTH-1:0]      m00_axi_awid,
    output wire [ADDR_WIDTH-1:0]    m00_axi_awaddr,
    output wire [7:0]               m00_axi_awlen,
    output wire [2:0]               m00_axi_awsize,
    output wire [1:0]               m00_axi_awburst,
    output wire                     m00_axi_awlock,
    output wire [3:0]               m00_axi_awcache,
    output wire [2:0]               m00_axi_awprot,
    output wire [3:0]               m00_axi_awqos,
    output wire [3:0]               m00_axi_awregion,
    output wire [AWUSER_WIDTH-1:0]  m00_axi_awuser,
    output wire                     m00_axi_awvalid,
    input  wire                     m00_axi_awready,
    output wire [DATA_WIDTH-1:0]    m00_axi_wdata,
    output wire [STRB_WIDTH-1:0]    m00_axi_wstrb,
    output wire                     m00_axi_wlast,
    output wire [WUSER_WIDTH-1:0]   m00_axi_wuser,
    output wire                     m00_axi_wvalid,
    input  wire                     m00_axi_wready,
    input  wire [ID_WIDTH-1:0]      m00_axi_bid,
    input  wire [1:0]               m00_axi_bresp,
    input  wire [BUSER_WIDTH-1:0]   m00_axi_buser,
    input  wire                     m00_axi_bvalid,
    output wire                     m00_axi_bready,
    output wire [ID_WIDTH-1:0]      m00_axi_arid,
    output wire [ADDR_WIDTH-1:0]    m00_axi_araddr,
    output wire [7:0]               m00_axi_arlen,
    output wire [2:0]               m00_axi_arsize,
    output wire [1:0]               m00_axi_arburst,
    output wire                     m00_axi_arlock,
    output wire [3:0]               m00_axi_arcache,
    output wire [2:0]               m00_axi_arprot,
    output wire [3:0]               m00_axi_arqos,
    output wire [3:0]               m00_axi_arregion,
    output wire [ARUSER_WIDTH-1:0]  m00_axi_aruser,
    output wire                     m00_axi_arvalid,
    input  wire                     m00_axi_arready,
    input  wire [ID_WIDTH-1:0]      m00_axi_rid,
    input  wire [DATA_WIDTH-1:0]    m00_axi_rdata,
    input  wire [1:0]               m00_axi_rresp,
    input  wire                     m00_axi_rlast,
    input  wire [RUSER_WIDTH-1:0]   m00_axi_ruser,
    input  wire                     m00_axi_rvalid,
    output wire                     m00_axi_rready,

    output wire [ID_WIDTH-1:0]      m01_axi_awid,
    output wire [ADDR_WIDTH-1:0]    m01_axi_awaddr,
    output wire [7:0]               m01_axi_awlen,
    output wire [2:0]               m01_axi_awsize,
    output wire [1:0]               m01_axi_awburst,
    output wire                     m01_axi_awlock,
    output wire [3:0]               m01_axi_awcache,
    output wire [2:0]               m01_axi_awprot,
    output wire [3:0]               m01_axi_awqos,
    output wire [3:0]               m01_axi_awregion,
    output wire [AWUSER_WIDTH-1:0]  m01_axi_awuser,
    output wire                     m01_axi_awvalid,
    input  wire                     m01_axi_awready,
    output wire [DATA_WIDTH-1:0]    m01_axi_wdata,
    output wire [STRB_WIDTH-1:0]    m01_axi_wstrb,
    output wire                     m01_axi_wlast,
    output wire [WUSER_WIDTH-1:0]   m01_axi_wuser,
    output wire                     m01_axi_wvalid,
    input  wire                     m01_axi_wready,
    input  wire [ID_WIDTH-1:0]      m01_axi_bid,
    input  wire [1:0]               m01_axi_bresp,
    input  wire [BUSER_WIDTH-1:0]   m01_axi_buser,
    input  wire                     m01_axi_bvalid,
    output wire                     m01_axi_bready,
    output wire [ID_WIDTH-1:0]      m01_axi_arid,
    output wire [ADDR_WIDTH-1:0]    m01_axi_araddr,
    output wire [7:0]               m01_axi_arlen,
    output wire [2:0]               m01_axi_arsize,
    output wire [1:0]               m01_axi_arburst,
    output wire                     m01_axi_arlock,
    output wire [3:0]               m01_axi_arcache,
    output wire [2:0]               m01_axi_arprot,
    output wire [3:0]               m01_axi_arqos,
    output wire [3:0]               m01_axi_arregion,
    output wire [ARUSER_WIDTH-1:0]  m01_axi_aruser,
    output wire                     m01_axi_arvalid,
    input  wire                     m01_axi_arready,
    input  wire [ID_WIDTH-1:0]      m01_axi_rid,
    input  wire [DATA_WIDTH-1:0]    m01_axi_rdata,
    input  wire [1:0]               m01_axi_rresp,
    input  wire                     m01_axi_rlast,
    input  wire [RUSER_WIDTH-1:0]   m01_axi_ruser,
    input  wire                     m01_axi_rvalid,
    output wire                     m01_axi_rready
);

localparam S_COUNT = 28;
localparam M_COUNT = 2;

// parameter sizing helpers
function [ADDR_WIDTH*M_REGIONS-1:0] w_a_r(input [ADDR_WIDTH*M_REGIONS-1:0] val);
    w_a_r = val;
endfunction

function [32*M_REGIONS-1:0] w_32_r(input [32*M_REGIONS-1:0] val);
    w_32_r = val;
endfunction

function [S_COUNT-1:0] w_s(input [S_COUNT-1:0] val);
    w_s = val;
endfunction

function w_1(input val);
    w_1 = val;
endfunction

axi_interconnect #(
    .S_COUNT(S_COUNT),
    .M_COUNT(M_COUNT),
    .DATA_WIDTH(DATA_WIDTH),
    .ADDR_WIDTH(ADDR_WIDTH),
    .STRB_WIDTH(STRB_WIDTH),
    .ID_WIDTH(ID_WIDTH),
    .AWUSER_ENABLE(AWUSER_ENABLE),
    .AWUSER_WIDTH(AWUSER_WIDTH),
    .WUSER_ENABLE(WUSER_ENABLE),
    .WUSER_WIDTH(WUSER_WIDTH),
    .BUSER_ENABLE(BUSER_ENABLE),
    .BUSER_WIDTH(BUSER_WIDTH),
    .ARUSER_ENABLE(ARUSER_ENABLE),
    .ARUSER_WIDTH(ARUSER_WIDTH),
    .RUSER_ENABLE(RUSER_ENABLE),
    .RUSER_WIDTH(RUSER_WIDTH),
    .FORWARD_ID(FORWARD_ID),
    .M_REGIONS(M_REGIONS),
    .M_BASE_ADDR({ w_a_r(M01_BASE_ADDR), w_a_r(M00_BASE_ADDR) }),
    .M_ADDR_WIDTH({ w_32_r(M01_ADDR_WIDTH), w_32_r(M00_ADDR_WIDTH) }),
    .M_CONNECT_READ({ w_s(M01_CONNECT_READ), w_s(M00_CONNECT_READ) }),
    .M_CONNECT_WRITE({ w_s(M01_CONNECT_WRITE), w_s(M00_CONNECT_WRITE) }),
    .M_SECURE({ w_1(M01_SECURE), w_1(M00_SECURE) })
)
axi_interconnect_inst (
    .clk(clk),
    .rst(rst),
    .s_axi_awid({ s27_axi_awid, s26_axi_awid, s25_axi_awid, s24_axi_awid, s23_axi_awid, s22_axi_awid, s21_axi_awid, s20_axi_awid, s19_axi_awid, s18_axi_awid, s17_axi_awid, s16_axi_awid, s15_axi_awid, s14_axi_awid, s13_axi_awid, s12_axi_awid, s11_axi_awid, s10_axi_awid, s09_axi_awid, s08_axi_awid, s07_axi_awid, s06_axi_awid, s05_axi_awid, s04_axi_awid, s03_axi_awid, s02_axi_awid, s01_axi_awid, s00_axi_awid }),
    .s_axi_awaddr({ s27_axi_awaddr, s26_axi_awaddr, s25_axi_awaddr, s24_axi_awaddr, s23_axi_awaddr, s22_axi_awaddr, s21_axi_awaddr, s20_axi_awaddr, s19_axi_awaddr, s18_axi_awaddr, s17_axi_awaddr, s16_axi_awaddr, s15_axi_awaddr, s14_axi_awaddr, s13_axi_awaddr, s12_axi_awaddr, s11_axi_awaddr, s10_axi_awaddr, s09_axi_awaddr, s08_axi_awaddr, s07_axi_awaddr, s06_axi_awaddr, s05_axi_awaddr, s04_axi_awaddr, s03_axi_awaddr, s02_axi_awaddr, s01_axi_awaddr, s00_axi_awaddr }),
    .s_axi_awlen({ s27_axi_awlen, s26_axi_awlen, s25_axi_awlen, s24_axi_awlen, s23_axi_awlen, s22_axi_awlen, s21_axi_awlen, s20_axi_awlen, s19_axi_awlen, s18_axi_awlen, s17_axi_awlen, s16_axi_awlen, s15_axi_awlen, s14_axi_awlen, s13_axi_awlen, s12_axi_awlen, s11_axi_awlen, s10_axi_awlen, s09_axi_awlen, s08_axi_awlen, s07_axi_awlen, s06_axi_awlen, s05_axi_awlen, s04_axi_awlen, s03_axi_awlen, s02_axi_awlen, s01_axi_awlen, s00_axi_awlen }),
    .s_axi_awsize({ s27_axi_awsize, s26_axi_awsize, s25_axi_awsize, s24_axi_awsize, s23_axi_awsize, s22_axi_awsize, s21_axi_awsize, s20_axi_awsize, s19_axi_awsize, s18_axi_awsize, s17_axi_awsize, s16_axi_awsize, s15_axi_awsize, s14_axi_awsize, s13_axi_awsize, s12_axi_awsize, s11_axi_awsize, s10_axi_awsize, s09_axi_awsize, s08_axi_awsize, s07_axi_awsize, s06_axi_awsize, s05_axi_awsize, s04_axi_awsize, s03_axi_awsize, s02_axi_awsize, s01_axi_awsize, s00_axi_awsize }),
    .s_axi_awburst({ s27_axi_awburst, s26_axi_awburst, s25_axi_awburst, s24_axi_awburst, s23_axi_awburst, s22_axi_awburst, s21_axi_awburst, s20_axi_awburst, s19_axi_awburst, s18_axi_awburst, s17_axi_awburst, s16_axi_awburst, s15_axi_awburst, s14_axi_awburst, s13_axi_awburst, s12_axi_awburst, s11_axi_awburst, s10_axi_awburst, s09_axi_awburst, s08_axi_awburst, s07_axi_awburst, s06_axi_awburst, s05_axi_awburst, s04_axi_awburst, s03_axi_awburst, s02_axi_awburst, s01_axi_awburst, s00_axi_awburst }),
    .s_axi_awlock({ s27_axi_awlock, s26_axi_awlock, s25_axi_awlock, s24_axi_awlock, s23_axi_awlock, s22_axi_awlock, s21_axi_awlock, s20_axi_awlock, s19_axi_awlock, s18_axi_awlock, s17_axi_awlock, s16_axi_awlock, s15_axi_awlock, s14_axi_awlock, s13_axi_awlock, s12_axi_awlock, s11_axi_awlock, s10_axi_awlock, s09_axi_awlock, s08_axi_awlock, s07_axi_awlock, s06_axi_awlock, s05_axi_awlock, s04_axi_awlock, s03_axi_awlock, s02_axi_awlock, s01_axi_awlock, s00_axi_awlock }),
    .s_axi_awcache({ s27_axi_awcache, s26_axi_awcache, s25_axi_awcache, s24_axi_awcache, s23_axi_awcache, s22_axi_awcache, s21_axi_awcache, s20_axi_awcache, s19_axi_awcache, s18_axi_awcache, s17_axi_awcache, s16_axi_awcache, s15_axi_awcache, s14_axi_awcache, s13_axi_awcache, s12_axi_awcache, s11_axi_awcache, s10_axi_awcache, s09_axi_awcache, s08_axi_awcache, s07_axi_awcache, s06_axi_awcache, s05_axi_awcache, s04_axi_awcache, s03_axi_awcache, s02_axi_awcache, s01_axi_awcache, s00_axi_awcache }),
    .s_axi_awprot({ s27_axi_awprot, s26_axi_awprot, s25_axi_awprot, s24_axi_awprot, s23_axi_awprot, s22_axi_awprot, s21_axi_awprot, s20_axi_awprot, s19_axi_awprot, s18_axi_awprot, s17_axi_awprot, s16_axi_awprot, s15_axi_awprot, s14_axi_awprot, s13_axi_awprot, s12_axi_awprot, s11_axi_awprot, s10_axi_awprot, s09_axi_awprot, s08_axi_awprot, s07_axi_awprot, s06_axi_awprot, s05_axi_awprot, s04_axi_awprot, s03_axi_awprot, s02_axi_awprot, s01_axi_awprot, s00_axi_awprot }),
    .s_axi_awqos({ s27_axi_awqos, s26_axi_awqos, s25_axi_awqos, s24_axi_awqos, s23_axi_awqos, s22_axi_awqos, s21_axi_awqos, s20_axi_awqos, s19_axi_awqos, s18_axi_awqos, s17_axi_awqos, s16_axi_awqos, s15_axi_awqos, s14_axi_awqos, s13_axi_awqos, s12_axi_awqos, s11_axi_awqos, s10_axi_awqos, s09_axi_awqos, s08_axi_awqos, s07_axi_awqos, s06_axi_awqos, s05_axi_awqos, s04_axi_awqos, s03_axi_awqos, s02_axi_awqos, s01_axi_awqos, s00_axi_awqos }),
    .s_axi_awuser({ s27_axi_awuser, s26_axi_awuser, s25_axi_awuser, s24_axi_awuser, s23_axi_awuser, s22_axi_awuser, s21_axi_awuser, s20_axi_awuser, s19_axi_awuser, s18_axi_awuser, s17_axi_awuser, s16_axi_awuser, s15_axi_awuser, s14_axi_awuser, s13_axi_awuser, s12_axi_awuser, s11_axi_awuser, s10_axi_awuser, s09_axi_awuser, s08_axi_awuser, s07_axi_awuser, s06_axi_awuser, s05_axi_awuser, s04_axi_awuser, s03_axi_awuser, s02_axi_awuser, s01_axi_awuser, s00_axi_awuser }),
    .s_axi_awvalid({ s27_axi_awvalid, s26_axi_awvalid, s25_axi_awvalid, s24_axi_awvalid, s23_axi_awvalid, s22_axi_awvalid, s21_axi_awvalid, s20_axi_awvalid, s19_axi_awvalid, s18_axi_awvalid, s17_axi_awvalid, s16_axi_awvalid, s15_axi_awvalid, s14_axi_awvalid, s13_axi_awvalid, s12_axi_awvalid, s11_axi_awvalid, s10_axi_awvalid, s09_axi_awvalid, s08_axi_awvalid, s07_axi_awvalid, s06_axi_awvalid, s05_axi_awvalid, s04_axi_awvalid, s03_axi_awvalid, s02_axi_awvalid, s01_axi_awvalid, s00_axi_awvalid }),
    .s_axi_awready({ s27_axi_awready, s26_axi_awready, s25_axi_awready, s24_axi_awready, s23_axi_awready, s22_axi_awready, s21_axi_awready, s20_axi_awready, s19_axi_awready, s18_axi_awready, s17_axi_awready, s16_axi_awready, s15_axi_awready, s14_axi_awready, s13_axi_awready, s12_axi_awready, s11_axi_awready, s10_axi_awready, s09_axi_awready, s08_axi_awready, s07_axi_awready, s06_axi_awready, s05_axi_awready, s04_axi_awready, s03_axi_awready, s02_axi_awready, s01_axi_awready, s00_axi_awready }),
    .s_axi_wdata({ s27_axi_wdata, s26_axi_wdata, s25_axi_wdata, s24_axi_wdata, s23_axi_wdata, s22_axi_wdata, s21_axi_wdata, s20_axi_wdata, s19_axi_wdata, s18_axi_wdata, s17_axi_wdata, s16_axi_wdata, s15_axi_wdata, s14_axi_wdata, s13_axi_wdata, s12_axi_wdata, s11_axi_wdata, s10_axi_wdata, s09_axi_wdata, s08_axi_wdata, s07_axi_wdata, s06_axi_wdata, s05_axi_wdata, s04_axi_wdata, s03_axi_wdata, s02_axi_wdata, s01_axi_wdata, s00_axi_wdata }),
    .s_axi_wstrb({ s27_axi_wstrb, s26_axi_wstrb, s25_axi_wstrb, s24_axi_wstrb, s23_axi_wstrb, s22_axi_wstrb, s21_axi_wstrb, s20_axi_wstrb, s19_axi_wstrb, s18_axi_wstrb, s17_axi_wstrb, s16_axi_wstrb, s15_axi_wstrb, s14_axi_wstrb, s13_axi_wstrb, s12_axi_wstrb, s11_axi_wstrb, s10_axi_wstrb, s09_axi_wstrb, s08_axi_wstrb, s07_axi_wstrb, s06_axi_wstrb, s05_axi_wstrb, s04_axi_wstrb, s03_axi_wstrb, s02_axi_wstrb, s01_axi_wstrb, s00_axi_wstrb }),
    .s_axi_wlast({ s27_axi_wlast, s26_axi_wlast, s25_axi_wlast, s24_axi_wlast, s23_axi_wlast, s22_axi_wlast, s21_axi_wlast, s20_axi_wlast, s19_axi_wlast, s18_axi_wlast, s17_axi_wlast, s16_axi_wlast, s15_axi_wlast, s14_axi_wlast, s13_axi_wlast, s12_axi_wlast, s11_axi_wlast, s10_axi_wlast, s09_axi_wlast, s08_axi_wlast, s07_axi_wlast, s06_axi_wlast, s05_axi_wlast, s04_axi_wlast, s03_axi_wlast, s02_axi_wlast, s01_axi_wlast, s00_axi_wlast }),
    .s_axi_wuser({ s27_axi_wuser, s26_axi_wuser, s25_axi_wuser, s24_axi_wuser, s23_axi_wuser, s22_axi_wuser, s21_axi_wuser, s20_axi_wuser, s19_axi_wuser, s18_axi_wuser, s17_axi_wuser, s16_axi_wuser, s15_axi_wuser, s14_axi_wuser, s13_axi_wuser, s12_axi_wuser, s11_axi_wuser, s10_axi_wuser, s09_axi_wuser, s08_axi_wuser, s07_axi_wuser, s06_axi_wuser, s05_axi_wuser, s04_axi_wuser, s03_axi_wuser, s02_axi_wuser, s01_axi_wuser, s00_axi_wuser }),
    .s_axi_wvalid({ s27_axi_wvalid, s26_axi_wvalid, s25_axi_wvalid, s24_axi_wvalid, s23_axi_wvalid, s22_axi_wvalid, s21_axi_wvalid, s20_axi_wvalid, s19_axi_wvalid, s18_axi_wvalid, s17_axi_wvalid, s16_axi_wvalid, s15_axi_wvalid, s14_axi_wvalid, s13_axi_wvalid, s12_axi_wvalid, s11_axi_wvalid, s10_axi_wvalid, s09_axi_wvalid, s08_axi_wvalid, s07_axi_wvalid, s06_axi_wvalid, s05_axi_wvalid, s04_axi_wvalid, s03_axi_wvalid, s02_axi_wvalid, s01_axi_wvalid, s00_axi_wvalid }),
    .s_axi_wready({ s27_axi_wready, s26_axi_wready, s25_axi_wready, s24_axi_wready, s23_axi_wready, s22_axi_wready, s21_axi_wready, s20_axi_wready, s19_axi_wready, s18_axi_wready, s17_axi_wready, s16_axi_wready, s15_axi_wready, s14_axi_wready, s13_axi_wready, s12_axi_wready, s11_axi_wready, s10_axi_wready, s09_axi_wready, s08_axi_wready, s07_axi_wready, s06_axi_wready, s05_axi_wready, s04_axi_wready, s03_axi_wready, s02_axi_wready, s01_axi_wready, s00_axi_wready }),
    .s_axi_bid({ s27_axi_bid, s26_axi_bid, s25_axi_bid, s24_axi_bid, s23_axi_bid, s22_axi_bid, s21_axi_bid, s20_axi_bid, s19_axi_bid, s18_axi_bid, s17_axi_bid, s16_axi_bid, s15_axi_bid, s14_axi_bid, s13_axi_bid, s12_axi_bid, s11_axi_bid, s10_axi_bid, s09_axi_bid, s08_axi_bid, s07_axi_bid, s06_axi_bid, s05_axi_bid, s04_axi_bid, s03_axi_bid, s02_axi_bid, s01_axi_bid, s00_axi_bid }),
    .s_axi_bresp({ s27_axi_bresp, s26_axi_bresp, s25_axi_bresp, s24_axi_bresp, s23_axi_bresp, s22_axi_bresp, s21_axi_bresp, s20_axi_bresp, s19_axi_bresp, s18_axi_bresp, s17_axi_bresp, s16_axi_bresp, s15_axi_bresp, s14_axi_bresp, s13_axi_bresp, s12_axi_bresp, s11_axi_bresp, s10_axi_bresp, s09_axi_bresp, s08_axi_bresp, s07_axi_bresp, s06_axi_bresp, s05_axi_bresp, s04_axi_bresp, s03_axi_bresp, s02_axi_bresp, s01_axi_bresp, s00_axi_bresp }),
    .s_axi_buser({ s27_axi_buser, s26_axi_buser, s25_axi_buser, s24_axi_buser, s23_axi_buser, s22_axi_buser, s21_axi_buser, s20_axi_buser, s19_axi_buser, s18_axi_buser, s17_axi_buser, s16_axi_buser, s15_axi_buser, s14_axi_buser, s13_axi_buser, s12_axi_buser, s11_axi_buser, s10_axi_buser, s09_axi_buser, s08_axi_buser, s07_axi_buser, s06_axi_buser, s05_axi_buser, s04_axi_buser, s03_axi_buser, s02_axi_buser, s01_axi_buser, s00_axi_buser }),
    .s_axi_bvalid({ s27_axi_bvalid, s26_axi_bvalid, s25_axi_bvalid, s24_axi_bvalid, s23_axi_bvalid, s22_axi_bvalid, s21_axi_bvalid, s20_axi_bvalid, s19_axi_bvalid, s18_axi_bvalid, s17_axi_bvalid, s16_axi_bvalid, s15_axi_bvalid, s14_axi_bvalid, s13_axi_bvalid, s12_axi_bvalid, s11_axi_bvalid, s10_axi_bvalid, s09_axi_bvalid, s08_axi_bvalid, s07_axi_bvalid, s06_axi_bvalid, s05_axi_bvalid, s04_axi_bvalid, s03_axi_bvalid, s02_axi_bvalid, s01_axi_bvalid, s00_axi_bvalid }),
    .s_axi_bready({ s27_axi_bready, s26_axi_bready, s25_axi_bready, s24_axi_bready, s23_axi_bready, s22_axi_bready, s21_axi_bready, s20_axi_bready, s19_axi_bready, s18_axi_bready, s17_axi_bready, s16_axi_bready, s15_axi_bready, s14_axi_bready, s13_axi_bready, s12_axi_bready, s11_axi_bready, s10_axi_bready, s09_axi_bready, s08_axi_bready, s07_axi_bready, s06_axi_bready, s05_axi_bready, s04_axi_bready, s03_axi_bready, s02_axi_bready, s01_axi_bready, s00_axi_bready }),
    .s_axi_arid({ s27_axi_arid, s26_axi_arid, s25_axi_arid, s24_axi_arid, s23_axi_arid, s22_axi_arid, s21_axi_arid, s20_axi_arid, s19_axi_arid, s18_axi_arid, s17_axi_arid, s16_axi_arid, s15_axi_arid, s14_axi_arid, s13_axi_arid, s12_axi_arid, s11_axi_arid, s10_axi_arid, s09_axi_arid, s08_axi_arid, s07_axi_arid, s06_axi_arid, s05_axi_arid, s04_axi_arid, s03_axi_arid, s02_axi_arid, s01_axi_arid, s00_axi_arid }),
    .s_axi_araddr({ s27_axi_araddr, s26_axi_araddr, s25_axi_araddr, s24_axi_araddr, s23_axi_araddr, s22_axi_araddr, s21_axi_araddr, s20_axi_araddr, s19_axi_araddr, s18_axi_araddr, s17_axi_araddr, s16_axi_araddr, s15_axi_araddr, s14_axi_araddr, s13_axi_araddr, s12_axi_araddr, s11_axi_araddr, s10_axi_araddr, s09_axi_araddr, s08_axi_araddr, s07_axi_araddr, s06_axi_araddr, s05_axi_araddr, s04_axi_araddr, s03_axi_araddr, s02_axi_araddr, s01_axi_araddr, s00_axi_araddr }),
    .s_axi_arlen({ s27_axi_arlen, s26_axi_arlen, s25_axi_arlen, s24_axi_arlen, s23_axi_arlen, s22_axi_arlen, s21_axi_arlen, s20_axi_arlen, s19_axi_arlen, s18_axi_arlen, s17_axi_arlen, s16_axi_arlen, s15_axi_arlen, s14_axi_arlen, s13_axi_arlen, s12_axi_arlen, s11_axi_arlen, s10_axi_arlen, s09_axi_arlen, s08_axi_arlen, s07_axi_arlen, s06_axi_arlen, s05_axi_arlen, s04_axi_arlen, s03_axi_arlen, s02_axi_arlen, s01_axi_arlen, s00_axi_arlen }),
    .s_axi_arsize({ s27_axi_arsize, s26_axi_arsize, s25_axi_arsize, s24_axi_arsize, s23_axi_arsize, s22_axi_arsize, s21_axi_arsize, s20_axi_arsize, s19_axi_arsize, s18_axi_arsize, s17_axi_arsize, s16_axi_arsize, s15_axi_arsize, s14_axi_arsize, s13_axi_arsize, s12_axi_arsize, s11_axi_arsize, s10_axi_arsize, s09_axi_arsize, s08_axi_arsize, s07_axi_arsize, s06_axi_arsize, s05_axi_arsize, s04_axi_arsize, s03_axi_arsize, s02_axi_arsize, s01_axi_arsize, s00_axi_arsize }),
    .s_axi_arburst({ s27_axi_arburst, s26_axi_arburst, s25_axi_arburst, s24_axi_arburst, s23_axi_arburst, s22_axi_arburst, s21_axi_arburst, s20_axi_arburst, s19_axi_arburst, s18_axi_arburst, s17_axi_arburst, s16_axi_arburst, s15_axi_arburst, s14_axi_arburst, s13_axi_arburst, s12_axi_arburst, s11_axi_arburst, s10_axi_arburst, s09_axi_arburst, s08_axi_arburst, s07_axi_arburst, s06_axi_arburst, s05_axi_arburst, s04_axi_arburst, s03_axi_arburst, s02_axi_arburst, s01_axi_arburst, s00_axi_arburst }),
    .s_axi_arlock({ s27_axi_arlock, s26_axi_arlock, s25_axi_arlock, s24_axi_arlock, s23_axi_arlock, s22_axi_arlock, s21_axi_arlock, s20_axi_arlock, s19_axi_arlock, s18_axi_arlock, s17_axi_arlock, s16_axi_arlock, s15_axi_arlock, s14_axi_arlock, s13_axi_arlock, s12_axi_arlock, s11_axi_arlock, s10_axi_arlock, s09_axi_arlock, s08_axi_arlock, s07_axi_arlock, s06_axi_arlock, s05_axi_arlock, s04_axi_arlock, s03_axi_arlock, s02_axi_arlock, s01_axi_arlock, s00_axi_arlock }),
    .s_axi_arcache({ s27_axi_arcache, s26_axi_arcache, s25_axi_arcache, s24_axi_arcache, s23_axi_arcache, s22_axi_arcache, s21_axi_arcache, s20_axi_arcache, s19_axi_arcache, s18_axi_arcache, s17_axi_arcache, s16_axi_arcache, s15_axi_arcache, s14_axi_arcache, s13_axi_arcache, s12_axi_arcache, s11_axi_arcache, s10_axi_arcache, s09_axi_arcache, s08_axi_arcache, s07_axi_arcache, s06_axi_arcache, s05_axi_arcache, s04_axi_arcache, s03_axi_arcache, s02_axi_arcache, s01_axi_arcache, s00_axi_arcache }),
    .s_axi_arprot({ s27_axi_arprot, s26_axi_arprot, s25_axi_arprot, s24_axi_arprot, s23_axi_arprot, s22_axi_arprot, s21_axi_arprot, s20_axi_arprot, s19_axi_arprot, s18_axi_arprot, s17_axi_arprot, s16_axi_arprot, s15_axi_arprot, s14_axi_arprot, s13_axi_arprot, s12_axi_arprot, s11_axi_arprot, s10_axi_arprot, s09_axi_arprot, s08_axi_arprot, s07_axi_arprot, s06_axi_arprot, s05_axi_arprot, s04_axi_arprot, s03_axi_arprot, s02_axi_arprot, s01_axi_arprot, s00_axi_arprot }),
    .s_axi_arqos({ s27_axi_arqos, s26_axi_arqos, s25_axi_arqos, s24_axi_arqos, s23_axi_arqos, s22_axi_arqos, s21_axi_arqos, s20_axi_arqos, s19_axi_arqos, s18_axi_arqos, s17_axi_arqos, s16_axi_arqos, s15_axi_arqos, s14_axi_arqos, s13_axi_arqos, s12_axi_arqos, s11_axi_arqos, s10_axi_arqos, s09_axi_arqos, s08_axi_arqos, s07_axi_arqos, s06_axi_arqos, s05_axi_arqos, s04_axi_arqos, s03_axi_arqos, s02_axi_arqos, s01_axi_arqos, s00_axi_arqos }),
    .s_axi_aruser({ s27_axi_aruser, s26_axi_aruser, s25_axi_aruser, s24_axi_aruser, s23_axi_aruser, s22_axi_aruser, s21_axi_aruser, s20_axi_aruser, s19_axi_aruser, s18_axi_aruser, s17_axi_aruser, s16_axi_aruser, s15_axi_aruser, s14_axi_aruser, s13_axi_aruser, s12_axi_aruser, s11_axi_aruser, s10_axi_aruser, s09_axi_aruser, s08_axi_aruser, s07_axi_aruser, s06_axi_aruser, s05_axi_aruser, s04_axi_aruser, s03_axi_aruser, s02_axi_aruser, s01_axi_aruser, s00_axi_aruser }),
    .s_axi_arvalid({ s27_axi_arvalid, s26_axi_arvalid, s25_axi_arvalid, s24_axi_arvalid, s23_axi_arvalid, s22_axi_arvalid, s21_axi_arvalid, s20_axi_arvalid, s19_axi_arvalid, s18_axi_arvalid, s17_axi_arvalid, s16_axi_arvalid, s15_axi_arvalid, s14_axi_arvalid, s13_axi_arvalid, s12_axi_arvalid, s11_axi_arvalid, s10_axi_arvalid, s09_axi_arvalid, s08_axi_arvalid, s07_axi_arvalid, s06_axi_arvalid, s05_axi_arvalid, s04_axi_arvalid, s03_axi_arvalid, s02_axi_arvalid, s01_axi_arvalid, s00_axi_arvalid }),
    .s_axi_arready({ s27_axi_arready, s26_axi_arready, s25_axi_arready, s24_axi_arready, s23_axi_arready, s22_axi_arready, s21_axi_arready, s20_axi_arready, s19_axi_arready, s18_axi_arready, s17_axi_arready, s16_axi_arready, s15_axi_arready, s14_axi_arready, s13_axi_arready, s12_axi_arready, s11_axi_arready, s10_axi_arready, s09_axi_arready, s08_axi_arready, s07_axi_arready, s06_axi_arready, s05_axi_arready, s04_axi_arready, s03_axi_arready, s02_axi_arready, s01_axi_arready, s00_axi_arready }),
    .s_axi_rid({ s27_axi_rid, s26_axi_rid, s25_axi_rid, s24_axi_rid, s23_axi_rid, s22_axi_rid, s21_axi_rid, s20_axi_rid, s19_axi_rid, s18_axi_rid, s17_axi_rid, s16_axi_rid, s15_axi_rid, s14_axi_rid, s13_axi_rid, s12_axi_rid, s11_axi_rid, s10_axi_rid, s09_axi_rid, s08_axi_rid, s07_axi_rid, s06_axi_rid, s05_axi_rid, s04_axi_rid, s03_axi_rid, s02_axi_rid, s01_axi_rid, s00_axi_rid }),
    .s_axi_rdata({ s27_axi_rdata, s26_axi_rdata, s25_axi_rdata, s24_axi_rdata, s23_axi_rdata, s22_axi_rdata, s21_axi_rdata, s20_axi_rdata, s19_axi_rdata, s18_axi_rdata, s17_axi_rdata, s16_axi_rdata, s15_axi_rdata, s14_axi_rdata, s13_axi_rdata, s12_axi_rdata, s11_axi_rdata, s10_axi_rdata, s09_axi_rdata, s08_axi_rdata, s07_axi_rdata, s06_axi_rdata, s05_axi_rdata, s04_axi_rdata, s03_axi_rdata, s02_axi_rdata, s01_axi_rdata, s00_axi_rdata }),
    .s_axi_rresp({ s27_axi_rresp, s26_axi_rresp, s25_axi_rresp, s24_axi_rresp, s23_axi_rresp, s22_axi_rresp, s21_axi_rresp, s20_axi_rresp, s19_axi_rresp, s18_axi_rresp, s17_axi_rresp, s16_axi_rresp, s15_axi_rresp, s14_axi_rresp, s13_axi_rresp, s12_axi_rresp, s11_axi_rresp, s10_axi_rresp, s09_axi_rresp, s08_axi_rresp, s07_axi_rresp, s06_axi_rresp, s05_axi_rresp, s04_axi_rresp, s03_axi_rresp, s02_axi_rresp, s01_axi_rresp, s00_axi_rresp }),
    .s_axi_rlast({ s27_axi_rlast, s26_axi_rlast, s25_axi_rlast, s24_axi_rlast, s23_axi_rlast, s22_axi_rlast, s21_axi_rlast, s20_axi_rlast, s19_axi_rlast, s18_axi_rlast, s17_axi_rlast, s16_axi_rlast, s15_axi_rlast, s14_axi_rlast, s13_axi_rlast, s12_axi_rlast, s11_axi_rlast, s10_axi_rlast, s09_axi_rlast, s08_axi_rlast, s07_axi_rlast, s06_axi_rlast, s05_axi_rlast, s04_axi_rlast, s03_axi_rlast, s02_axi_rlast, s01_axi_rlast, s00_axi_rlast }),
    .s_axi_ruser({ s27_axi_ruser, s26_axi_ruser, s25_axi_ruser, s24_axi_ruser, s23_axi_ruser, s22_axi_ruser, s21_axi_ruser, s20_axi_ruser, s19_axi_ruser, s18_axi_ruser, s17_axi_ruser, s16_axi_ruser, s15_axi_ruser, s14_axi_ruser, s13_axi_ruser, s12_axi_ruser, s11_axi_ruser, s10_axi_ruser, s09_axi_ruser, s08_axi_ruser, s07_axi_ruser, s06_axi_ruser, s05_axi_ruser, s04_axi_ruser, s03_axi_ruser, s02_axi_ruser, s01_axi_ruser, s00_axi_ruser }),
    .s_axi_rvalid({ s27_axi_rvalid, s26_axi_rvalid, s25_axi_rvalid, s24_axi_rvalid, s23_axi_rvalid, s22_axi_rvalid, s21_axi_rvalid, s20_axi_rvalid, s19_axi_rvalid, s18_axi_rvalid, s17_axi_rvalid, s16_axi_rvalid, s15_axi_rvalid, s14_axi_rvalid, s13_axi_rvalid, s12_axi_rvalid, s11_axi_rvalid, s10_axi_rvalid, s09_axi_rvalid, s08_axi_rvalid, s07_axi_rvalid, s06_axi_rvalid, s05_axi_rvalid, s04_axi_rvalid, s03_axi_rvalid, s02_axi_rvalid, s01_axi_rvalid, s00_axi_rvalid }),
    .s_axi_rready({ s27_axi_rready, s26_axi_rready, s25_axi_rready, s24_axi_rready, s23_axi_rready, s22_axi_rready, s21_axi_rready, s20_axi_rready, s19_axi_rready, s18_axi_rready, s17_axi_rready, s16_axi_rready, s15_axi_rready, s14_axi_rready, s13_axi_rready, s12_axi_rready, s11_axi_rready, s10_axi_rready, s09_axi_rready, s08_axi_rready, s07_axi_rready, s06_axi_rready, s05_axi_rready, s04_axi_rready, s03_axi_rready, s02_axi_rready, s01_axi_rready, s00_axi_rready }),
    .m_axi_awid({ m01_axi_awid, m00_axi_awid }),
    .m_axi_awaddr({ m01_axi_awaddr, m00_axi_awaddr }),
    .m_axi_awlen({ m01_axi_awlen, m00_axi_awlen }),
    .m_axi_awsize({ m01_axi_awsize, m00_axi_awsize }),
    .m_axi_awburst({ m01_axi_awburst, m00_axi_awburst }),
    .m_axi_awlock({ m01_axi_awlock, m00_axi_awlock }),
    .m_axi_awcache({ m01_axi_awcache, m00_axi_awcache }),
    .m_axi_awprot({ m01_axi_awprot, m00_axi_awprot }),
    .m_axi_awqos({ m01_axi_awqos, m00_axi_awqos }),
    .m_axi_awregion({ m01_axi_awregion, m00_axi_awregion }),
    .m_axi_awuser({ m01_axi_awuser, m00_axi_awuser }),
    .m_axi_awvalid({ m01_axi_awvalid, m00_axi_awvalid }),
    .m_axi_awready({ m01_axi_awready, m00_axi_awready }),
    .m_axi_wdata({ m01_axi_wdata, m00_axi_wdata }),
    .m_axi_wstrb({ m01_axi_wstrb, m00_axi_wstrb }),
    .m_axi_wlast({ m01_axi_wlast, m00_axi_wlast }),
    .m_axi_wuser({ m01_axi_wuser, m00_axi_wuser }),
    .m_axi_wvalid({ m01_axi_wvalid, m00_axi_wvalid }),
    .m_axi_wready({ m01_axi_wready, m00_axi_wready }),
    .m_axi_bid({ m01_axi_bid, m00_axi_bid }),
    .m_axi_bresp({ m01_axi_bresp, m00_axi_bresp }),
    .m_axi_buser({ m01_axi_buser, m00_axi_buser }),
    .m_axi_bvalid({ m01_axi_bvalid, m00_axi_bvalid }),
    .m_axi_bready({ m01_axi_bready, m00_axi_bready }),
    .m_axi_arid({ m01_axi_arid, m00_axi_arid }),
    .m_axi_araddr({ m01_axi_araddr, m00_axi_araddr }),
    .m_axi_arlen({ m01_axi_arlen, m00_axi_arlen }),
    .m_axi_arsize({ m01_axi_arsize, m00_axi_arsize }),
    .m_axi_arburst({ m01_axi_arburst, m00_axi_arburst }),
    .m_axi_arlock({ m01_axi_arlock, m00_axi_arlock }),
    .m_axi_arcache({ m01_axi_arcache, m00_axi_arcache }),
    .m_axi_arprot({ m01_axi_arprot, m00_axi_arprot }),
    .m_axi_arqos({ m01_axi_arqos, m00_axi_arqos }),
    .m_axi_arregion({ m01_axi_arregion, m00_axi_arregion }),
    .m_axi_aruser({ m01_axi_aruser, m00_axi_aruser }),
    .m_axi_arvalid({ m01_axi_arvalid, m00_axi_arvalid }),
    .m_axi_arready({ m01_axi_arready, m00_axi_arready }),
    .m_axi_rid({ m01_axi_rid, m00_axi_rid }),
    .m_axi_rdata({ m01_axi_rdata, m00_axi_rdata }),
    .m_axi_rresp({ m01_axi_rresp, m00_axi_rresp }),
    .m_axi_rlast({ m01_axi_rlast, m00_axi_rlast }),
    .m_axi_ruser({ m01_axi_ruser, m00_axi_ruser }),
    .m_axi_rvalid({ m01_axi_rvalid, m00_axi_rvalid }),
    .m_axi_rready({ m01_axi_rready, m00_axi_rready })
);

endmodule

`resetall
