/*
 * Ultra wide range test
*/

`define WIDTH 256
`define operator buf
`include "../.generic/range_any_width_unary_test.v"