/*
 * Ultra wide range test
*/

`define WIDTH 256
`define operator not
`include "range_any_width_unary_test.v"