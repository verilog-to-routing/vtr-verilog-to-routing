module test3(input a, output b);
    wire c;
    assign c = a;
    assign b = c;
endmodule