/*
 * Wide range test
*/

`define WIDTH 3
`define operator notif1
`include "../.generic/replicate_any_width_binary_test.v"