
 module ex2PM16_fir(clk, In_X, Out_Y); 

 input clk;
 input [11:0] In_X; 
 output [28 :0] Out_Y; 

 reg [11:0] x0 ;

 wire [14:0] x1 ;
 wire [16:0] x5 ;
 wire [21:0] x41 ;
 wire [21:0] x41_0_1 ;
 wire [21:0] y50 ;
 wire [21:0] x41_1_1 ;
 wire [21:0] y68 ;
 wire [22:0] x49 ;
 wire [22:0] x49_0_1 ;
 wire [22:0] y37 ;
 wire [22:0] x49_1_1 ;
 wire [22:0] y81 ;
 wire [22:0] x50 ;
 wire [22:0] x50_0_1 ;
 wire [22:0] y38 ;
 wire [22:0] x50_1_1 ;
 wire [22:0] y80 ;
 wire [24:0] x63 ;
 wire [24:0] x63_0_1 ;
 wire [24:0] y45 ;
 wire [24:0] x63_1_1 ;
 wire [24:0] y73 ;
 wire [28:0] x64 ;
 wire [28:0] x64_0_1 ;
 wire [28:0] y58 ;
 wire [28:0] x64_1_1 ;
 wire [28:0] y60 ;
 wire [19:0] x66 ;
 wire [19:0] x80 ;
 wire [20:0] y32 ;
 wire [19:0] x67 ;
 wire [19:0] x81 ;
 wire [19:0] y34 ;
 wire [21:0] x68 ;
 wire [21:0] x68_0_1 ;
 wire [23:0] y47 ;
 wire [21:0] x69 ;
 wire [21:0] x69_0_1 ;
 wire [23:0] y71 ;
 wire [19:0] x70 ;
 wire [19:0] x88 ;
 wire [19:0] y84 ;
 wire [19:0] x71 ;
 wire [19:0] x89 ;
 wire [20:0] y86 ;
 wire [19:0] x6 ;
 wire [22:0] x31 ;
 wire [22:0] x31_0_1 ;
 wire [23:0] y15 ;
 wire [22:0] x31_1_1 ;
 wire [23:0] y103 ;
 wire [23:0] x51 ;
 wire [23:0] x87 ;
 wire [25:0] y56 ;
 wire [25:0] y62 ;
 wire [26:0] x61 ;
 wire [26:0] x86 ;
 wire [26:0] y53 ;
 wire [26:0] y65 ;
 wire [19:0] x6_3_1 ;
 wire [19:0] x6_3_2 ;
 wire [22:0] y36 ;
 wire [19:0] x6_4_1 ;
 wire [19:0] x6_4_2 ;
 wire [22:0] y82 ;
 wire [18:0] x10 ;
 wire [18:0] x10_0_1 ;
 wire [18:0] x10_0_2 ;
 wire [20:0] y3 ;
 wire [18:0] x10_1_1 ;
 wire [18:0] x10_1_2 ;
 wire [20:0] y20 ;
 wire [18:0] x10_2_1 ;
 wire [18:0] x10_2_2 ;
 wire [20:0] y98 ;
 wire [18:0] x10_3_1 ;
 wire [18:0] x10_3_2 ;
 wire [20:0] y115 ;
 wire [22:0] x11 ;
 wire [23:0] x45 ;
 wire [23:0] x76 ;
 wire [23:0] y22 ;
 wire [23:0] y96 ;
 wire [23:0] x52 ;
 wire [23:0] x52_0_1 ;
 wire [23:0] y17 ;
 wire [23:0] x52_1_1 ;
 wire [23:0] y101 ;
 wire [17:0] x12 ;
 wire [22:0] x53 ;
 wire [22:0] x82 ;
 wire [22:0] y35 ;
 wire [22:0] y83 ;
 wire [24:0] x65 ;
 wire [24:0] x65_0_1 ;
 wire [24:0] y54 ;
 wire [24:0] x65_1_1 ;
 wire [24:0] y64 ;
 wire [20:0] x13 ;
 wire [25:0] x54 ;
 wire [25:0] x72 ;
 wire [25:0] y1 ;
 wire [25:0] y117 ;
 wire [20:0] x13_1_1 ;
 wire [20:0] x13_1_2 ;
 wire [21:0] y11 ;
 wire [20:0] x13_2_1 ;
 wire [20:0] x13_2_2 ;
 wire [21:0] y107 ;
 wire [24:0] x17 ;
 wire [25:0] x57 ;
 wire [25:0] x73 ;
 wire [25:0] y2 ;
 wire [25:0] y116 ;
 wire [20:0] x18 ;
 wire [20:0] x18_0_1 ;
 wire [20:0] x18_0_2 ;
 wire [20:0] y9 ;
 wire [20:0] x18_1_1 ;
 wire [20:0] x18_1_2 ;
 wire [20:0] y109 ;
 wire [21:0] x19 ;
 wire [22:0] x46 ;
 wire [22:0] x46_0_1 ;
 wire [22:0] y26 ;
 wire [22:0] x46_1_1 ;
 wire [22:0] y92 ;
 wire [23:0] x20 ;
 wire [22:0] x21 ;
 wire [22:0] x21_0_1 ;
 wire [22:0] x21_0_2 ;
 wire [22:0] y46 ;
 wire [22:0] x21_1_1 ;
 wire [22:0] x21_1_2 ;
 wire [22:0] y72 ;
 wire [16:0] x22 ;
 wire [20:0] x33 ;
 wire [20:0] x33_0_1 ;
 wire [20:0] x33_0_2 ;
 wire [22:0] y29 ;
 wire [20:0] x33_1_1 ;
 wire [20:0] x33_1_2 ;
 wire [22:0] y89 ;
 wire [21:0] x34 ;
 wire [26:0] x59 ;
 wire [26:0] x59_0_1 ;
 wire [26:0] y55 ;
 wire [26:0] x59_1_1 ;
 wire [26:0] y63 ;
 wire [25:0] x35 ;
 wire [26:0] x62 ;
 wire [26:0] x62_0_1 ;
 wire [26:0] y57 ;
 wire [26:0] x62_1_1 ;
 wire [26:0] y61 ;
 wire [23:0] x36 ;
 wire [23:0] x36_0_1 ;
 wire [23:0] x36_0_2 ;
 wire [23:0] y4 ;
 wire [23:0] x36_1_1 ;
 wire [23:0] x36_1_2 ;
 wire [23:0] y114 ;
 wire [20:0] x37 ;
 wire [20:0] x84 ;
 wire [20:0] x84_0_1 ;
 wire [23:0] y48 ;
 wire [20:0] x84_1_1 ;
 wire [23:0] y70 ;
 wire [20:0] x38 ;
 wire [20:0] x38_0_1 ;
 wire [20:0] x38_0_2 ;
 wire [21:0] y30 ;
 wire [20:0] x38_1_1 ;
 wire [20:0] x38_1_2 ;
 wire [21:0] y88 ;
 wire [20:0] x39 ;
 wire [20:0] x39_0_1 ;
 wire [20:0] x39_0_2 ;
 wire [22:0] y8 ;
 wire [20:0] x39_1_1 ;
 wire [20:0] x39_1_2 ;
 wire [22:0] y110 ;
 wire [21:0] x40 ;
 wire [21:0] x40_0_1 ;
 wire [21:0] x40_0_2 ;
 wire [24:0] y49 ;
 wire [21:0] x40_1_1 ;
 wire [21:0] x40_1_2 ;
 wire [24:0] y69 ;
 wire [21:0] x42 ;
 wire [21:0] x75 ;
 wire [21:0] x75_0_1 ;
 wire [22:0] y10 ;
 wire [21:0] x75_1_1 ;
 wire [22:0] y108 ;
 wire [22:0] x43 ;
 wire [22:0] x85 ;
 wire [22:0] x85_0_1 ;
 wire [23:0] y52 ;
 wire [22:0] x85_1_1 ;
 wire [23:0] y66 ;
 wire [23:0] x44 ;
 wire [23:0] x44_0_1 ;
 wire [23:0] y40 ;
 wire [23:0] x44_1_1 ;
 wire [23:0] y78 ;
 wire [14:0] x77 ;
 wire [14:0] x77_0_1 ;
 wire [14:0] x77_0_2 ;
 wire [20:0] y27 ;
 wire [14:0] x77_1_1 ;
 wire [14:0] x77_1_2 ;
 wire [20:0] y91 ;
 wire [14:0] x1_31_1 ;
 wire [14:0] x1_31_2 ;
 wire [14:0] x1_31_3 ;
 wire [16:0] y25 ;
 wire [14:0] x1_32_1 ;
 wire [14:0] x1_32_2 ;
 wire [14:0] x1_32_3 ;
 wire [16:0] y93 ;
 wire [14:0] x2 ;
 wire [17:0] x8 ;
 wire [17:0] x78 ;
 wire [17:0] x78_0_1 ;
 wire [21:0] y28 ;
 wire [17:0] x78_1_1 ;
 wire [21:0] y90 ;
 wire [17:0] x8_2_1 ;
 wire [17:0] x8_2_2 ;
 wire [19:0] y18 ;
 wire [17:0] x8_3_1 ;
 wire [17:0] x8_3_2 ;
 wire [19:0] y100 ;
 wire [17:0] x23 ;
 wire [17:0] x23_0_1 ;
 wire [17:0] x23_0_2 ;
 wire [19:0] y5 ;
 wire [17:0] x23_1_1 ;
 wire [17:0] x23_1_2 ;
 wire [19:0] y113 ;
 wire [18:0] x24 ;
 wire [18:0] x24_0_1 ;
 wire [18:0] x24_0_2 ;
 wire [20:0] y14 ;
 wire [18:0] x24_1_1 ;
 wire [18:0] x24_1_2 ;
 wire [20:0] y104 ;
 wire [19:0] x25 ;
 wire [19:0] x79 ;
 wire [19:0] x79_0_1 ;
 wire [21:0] y31 ;
 wire [19:0] x79_1_1 ;
 wire [21:0] y87 ;
 wire [22:0] x26 ;
 wire [23:0] x58 ;
 wire [23:0] x58_0_1 ;
 wire [23:0] y44 ;
 wire [23:0] x58_1_1 ;
 wire [23:0] y74 ;
 wire [20:0] x47 ;
 wire [20:0] x47_0_1 ;
 wire [20:0] x47_0_2 ;
 wire [20:0] y41 ;
 wire [20:0] x47_1_1 ;
 wire [20:0] x47_1_2 ;
 wire [20:0] y77 ;
 wire [21:0] x48 ;
 wire [21:0] x48_0_1 ;
 wire [21:0] x48_0_2 ;
 wire [21:0] y43 ;
 wire [21:0] x48_1_1 ;
 wire [21:0] x48_1_2 ;
 wire [21:0] y75 ;
 wire [21:0] x55 ;
 wire [21:0] x55_0_1 ;
 wire [21:0] x55_0_2 ;
 wire [21:0] y19 ;
 wire [21:0] x55_1_1 ;
 wire [21:0] x55_1_2 ;
 wire [21:0] y99 ;
 wire [23:0] x56 ;
 wire [23:0] x83 ;
 wire [23:0] x83_0_1 ;
 wire [23:0] y42 ;
 wire [23:0] x83_1_1 ;
 wire [23:0] y76 ;
 wire [14:0] x2_23_1 ;
 wire [14:0] x2_23_2 ;
 wire [14:0] x2_23_3 ;
 wire [21:0] y33 ;
 wire [14:0] x2_24_1 ;
 wire [14:0] x2_24_2 ;
 wire [14:0] x2_24_3 ;
 wire [21:0] y85 ;
 wire [15:0] x3 ;
 wire [20:0] x9 ;
 wire [20:0] x74 ;
 wire [20:0] x74_0_1 ;
 wire [21:0] y6 ;
 wire [20:0] x74_1_1 ;
 wire [20:0] y21 ;
 wire [20:0] x74_2_1 ;
 wire [20:0] y97 ;
 wire [20:0] x74_3_1 ;
 wire [21:0] y112 ;
 wire [20:0] x9_1_1 ;
 wire [20:0] x9_1_2 ;
 wire [20:0] y12 ;
 wire [20:0] x9_2_1 ;
 wire [20:0] x9_2_2 ;
 wire [20:0] y106 ;
 wire [21:0] x27 ;
 wire [21:0] x27_0_1 ;
 wire [21:0] x27_0_2 ;
 wire [21:0] y13 ;
 wire [21:0] x27_1_1 ;
 wire [21:0] x27_1_2 ;
 wire [21:0] y105 ;
 wire [18:0] x28 ;
 wire [18:0] x28_0_1 ;
 wire [18:0] x28_0_2 ;
 wire [21:0] y24 ;
 wire [18:0] x28_1_1 ;
 wire [18:0] x28_1_2 ;
 wire [21:0] y94 ;
 wire [27:0] x29 ;
 wire [24:0] x60 ;
 wire [24:0] x60_0_1 ;
 wire [24:0] x60_0_2 ;
 wire [24:0] y51 ;
 wire [24:0] x60_1_1 ;
 wire [24:0] x60_1_2 ;
 wire [24:0] y67 ;
 wire [15:0] x3_7_1 ;
 wire [15:0] x3_7_2 ;
 wire [15:0] x3_7_3 ;
 wire [19:0] y23 ;
 wire [15:0] x3_8_1 ;
 wire [15:0] x3_8_2 ;
 wire [15:0] x3_8_3 ;
 wire [19:0] y95 ;
 wire [15:0] x4 ;
 wire [21:0] x30 ;
 wire [21:0] x30_0_1 ;
 wire [21:0] x30_0_2 ;
 wire [22:0] y39 ;
 wire [21:0] x30_1_1 ;
 wire [21:0] x30_1_2 ;
 wire [22:0] y79 ;
 wire [15:0] x4_5_1 ;
 wire [15:0] x4_5_2 ;
 wire [15:0] x4_5_3 ;
 wire [17:0] y16 ;
 wire [15:0] x4_6_1 ;
 wire [15:0] x4_6_2 ;
 wire [15:0] x4_6_3 ;
 wire [17:0] y102 ;
 wire [16:0] x7 ;
 wire [20:0] x32 ;
 wire [20:0] x32_0_1 ;
 wire [20:0] x32_0_2 ;
 wire [21:0] y0 ;
 wire [20:0] x32_1_1 ;
 wire [20:0] x32_1_2 ;
 wire [21:0] y118 ;
 wire [16:0] x14 ;
 wire [17:0] x15 ;
 wire [17:0] x15_0_1 ;
 wire [17:0] x15_0_2 ;
 wire [17:0] x15_0_3 ;
 wire [17:0] y7 ;
 wire [17:0] x15_1_1 ;
 wire [17:0] x15_1_2 ;
 wire [17:0] x15_1_3 ;
 wire [17:0] y111 ;
 wire [22:0] x16 ;
 wire [11:0] x66_38_1 ;
 wire [11:0] x66_38_2 ;
 wire [11:0] x67_39_1 ;
 wire [11:0] x67_39_2 ;
 wire [11:0] x68_40_1 ;
 wire [11:0] x68_40_2 ;
 wire [11:0] x69_41_1 ;
 wire [11:0] x69_41_2 ;
 wire [11:0] x70_42_1 ;
 wire [11:0] x70_42_2 ;
 wire [11:0] x71_43_1 ;
 wire [11:0] x71_43_2 ;
 wire [11:0] x0_44_1 ;
 wire [11:0] x0_44_2 ;
 wire [11:0] x0_44_3 ;
 wire [11:0] x0_44_4 ;
 wire [26:0] y59 ;
 wire [21:0] x90 ;
 wire [26:0] x91 ;
 wire [26:0] x91_1 ;
 wire [27:0] x92 ;
 wire [27:0] x92_1 ;
 wire [28:0] x93 ;
 wire [28:0] x93_1 ;
 wire [28:0] x94 ;
 wire [28:0] x94_1 ;
 wire [28:0] x95 ;
 wire [28:0] x95_1 ;
 wire [28:0] x96 ;
 wire [28:0] x96_1 ;
 wire [28:0] x97 ;
 wire [28:0] x97_1 ;
 wire [28:0] x98 ;
 wire [28:0] x98_1 ;
 wire [28:0] x99 ;
 wire [28:0] x99_1 ;
 wire [28:0] x100 ;
 wire [28:0] x100_1 ;
 wire [28:0] x101 ;
 wire [28:0] x101_1 ;
 wire [28:0] x102 ;
 wire [28:0] x102_1 ;
 wire [28:0] x103 ;
 wire [28:0] x103_1 ;
 wire [28:0] x104 ;
 wire [28:0] x104_1 ;
 wire [28:0] x105 ;
 wire [28:0] x105_1 ;
 wire [28:0] x106 ;
 wire [28:0] x106_1 ;
 wire [28:0] x107 ;
 wire [28:0] x107_1 ;
 wire [28:0] x108 ;
 wire [28:0] x108_1 ;
 wire [28:0] x109 ;
 wire [28:0] x109_1 ;
 wire [28:0] x110 ;
 wire [28:0] x110_1 ;
 wire [28:0] x111 ;
 wire [28:0] x111_1 ;
 wire [28:0] x112 ;
 wire [28:0] x112_1 ;
 wire [28:0] x113 ;
 wire [28:0] x113_1 ;
 wire [28:0] x114 ;
 wire [28:0] x114_1 ;
 wire [28:0] x115 ;
 wire [28:0] x115_1 ;
 wire [28:0] x116 ;
 wire [28:0] x116_1 ;
 wire [28:0] x117 ;
 wire [28:0] x117_1 ;
 wire [28:0] x118 ;
 wire [28:0] x118_1 ;
 wire [28:0] x119 ;
 wire [28:0] x119_1 ;
 wire [28:0] x120 ;
 wire [28:0] x120_1 ;
 wire [28:0] x121 ;
 wire [28:0] x121_1 ;
 wire [28:0] x122 ;
 wire [28:0] x122_1 ;
 wire [28:0] x123 ;
 wire [28:0] x123_1 ;
 wire [28:0] x124 ;
 wire [28:0] x124_1 ;
 wire [28:0] x125 ;
 wire [28:0] x125_1 ;
 wire [28:0] x126 ;
 wire [28:0] x126_1 ;
 wire [28:0] x127 ;
 wire [28:0] x127_1 ;
 wire [28:0] x128 ;
 wire [28:0] x128_1 ;
 wire [28:0] x129 ;
 wire [28:0] x129_1 ;
 wire [28:0] x130 ;
 wire [28:0] x130_1 ;
 wire [28:0] x131 ;
 wire [28:0] x131_1 ;
 wire [28:0] x132 ;
 wire [28:0] x132_1 ;
 wire [28:0] x133 ;
 wire [28:0] x133_1 ;
 wire [28:0] x134 ;
 wire [28:0] x134_1 ;
 wire [28:0] x135 ;
 wire [28:0] x135_1 ;
 wire [28:0] x136 ;
 wire [28:0] x136_1 ;
 wire [28:0] x137 ;
 wire [28:0] x137_1 ;
 wire [28:0] x138 ;
 wire [28:0] x138_1 ;
 wire [28:0] x139 ;
 wire [28:0] x139_1 ;
 wire [28:0] x140 ;
 wire [28:0] x140_1 ;
 wire [28:0] x141 ;
 wire [28:0] x141_1 ;
 wire [28:0] x142 ;
 wire [28:0] x142_1 ;
 wire [28:0] x143 ;
 wire [28:0] x143_1 ;
 wire [28:0] x144 ;
 wire [28:0] x144_1 ;
 wire [28:0] x145 ;
 wire [28:0] x145_1 ;
 wire [28:0] x146 ;
 wire [28:0] x146_1 ;
 wire [28:0] x147 ;
 wire [28:0] x147_1 ;
 wire [28:0] x148 ;
 wire [28:0] x148_1 ;
 wire [28:0] x149 ;
 wire [28:0] x149_1 ;
 wire [28:0] x150 ;
 wire [28:0] x150_1 ;
 wire [28:0] x151 ;
 wire [28:0] x151_1 ;
 wire [28:0] x152 ;
 wire [28:0] x152_1 ;
 wire [28:0] x153 ;
 wire [28:0] x153_1 ;
 wire [28:0] x154 ;
 wire [28:0] x154_1 ;
 wire [28:0] x155 ;
 wire [28:0] x155_1 ;
 wire [28:0] x156 ;
 wire [28:0] x156_1 ;
 wire [28:0] x157 ;
 wire [28:0] x157_1 ;
 wire [28:0] x158 ;
 wire [28:0] x158_1 ;
 wire [28:0] x159 ;
 wire [28:0] x159_1 ;
 wire [28:0] x160 ;
 wire [28:0] x160_1 ;
 wire [28:0] x161 ;
 wire [28:0] x161_1 ;
 wire [28:0] x162 ;
 wire [28:0] x162_1 ;
 wire [28:0] x163 ;
 wire [28:0] x163_1 ;
 wire [28:0] x164 ;
 wire [28:0] x164_1 ;
 wire [28:0] x165 ;
 wire [28:0] x165_1 ;
 wire [28:0] x166 ;
 wire [28:0] x166_1 ;
 wire [28:0] x167 ;
 wire [28:0] x167_1 ;
 wire [28:0] x168 ;
 wire [28:0] x168_1 ;
 wire [28:0] x169 ;
 wire [28:0] x169_1 ;
 wire [28:0] x170 ;
 wire [28:0] x170_1 ;
 wire [28:0] x171 ;
 wire [28:0] x171_1 ;
 wire [28:0] x172 ;
 wire [28:0] x172_1 ;
 wire [28:0] x173 ;
 wire [28:0] x173_1 ;
 wire [28:0] x174 ;
 wire [28:0] x174_1 ;
 wire [28:0] x175 ;
 wire [28:0] x175_1 ;
 wire [28:0] x176 ;
 wire [28:0] x176_1 ;
 wire [28:0] x177 ;
 wire [28:0] x177_1 ;
 wire [28:0] x178 ;
 wire [28:0] x178_1 ;
 wire [28:0] x179 ;
 wire [28:0] x179_1 ;
 wire [28:0] x180 ;
 wire [28:0] x180_1 ;
 wire [28:0] x181 ;
 wire [28:0] x181_1 ;
 wire [28:0] x182 ;
 wire [28:0] x182_1 ;
 wire [28:0] x183 ;
 wire [28:0] x183_1 ;
 wire [28:0] x184 ;
 wire [28:0] x184_1 ;
 wire [28:0] x185 ;
 wire [28:0] x185_1 ;
 wire [28:0] x186 ;
 wire [28:0] x186_1 ;
 wire [28:0] x187 ;
 wire [28:0] x187_1 ;
 wire [28:0] x188 ;
 wire [28:0] x188_1 ;
 wire [28:0] x189 ;
 wire [28:0] x189_1 ;
 wire [28:0] x190 ;
 wire [28:0] x190_1 ;
 wire [28:0] x191 ;
 wire [28:0] x191_1 ;
 wire [28:0] x192 ;
 wire [28:0] x192_1 ;
 wire [28:0] x193 ;
 wire [28:0] x193_1 ;
 wire [28:0] x194 ;
 wire [28:0] x194_1 ;
 wire [28:0] x195 ;
 wire [28:0] x195_1 ;
 wire [28:0] x196 ;
 wire [28:0] x196_1 ;
 wire [28:0] x197 ;
 wire [28:0] x197_1 ;
 wire [28:0] x198 ;
 wire [28:0] x198_1 ;
 wire [28:0] x199 ;
 wire [28:0] x199_1 ;
 wire [28:0] x200 ;
 wire [28:0] x200_1 ;
 wire [28:0] x201 ;
 wire [28:0] x201_1 ;
 wire [28:0] x202 ;
 wire [28:0] x202_1 ;
 wire [28:0] x203 ;
 wire [28:0] x203_1 ;
 wire [28:0] x204 ;
 wire [28:0] x204_1 ;
 wire [28:0] x205 ;
 wire [28:0] x205_1 ;
 wire [28:0] x206 ;
 wire [28:0] x206_1 ;
 wire [28:0] x207 ;
 wire [28:0] x207_1 ;
 wire [28:0] Out_Y_wire ;
 reg [28:0] Out_Y;


 always @(posedge clk) 
 begin
 x0 <= In_X; 
 end 


 always @(posedge clk) 
 begin
 Out_Y = Out_Y_wire;
 end


 Subtractor14Bit Sub0(clk, { x0[11: 0], 2'b0 }, {x0[11],x0[11], x0[11: 0] }, x1); 


 Adder16Bit Adder0(clk,  { x0[11: 0], 4'b0 }, {x1[14], x1[14: 0]  }, x5); 


 Subtractor21Bit Sub1(clk, {x5[16],x5[16],x5[16],x5[16], x5[16: 0] },  { x1[14: 0], 6'b0 },x41); 

 Register22Bit Reg0 (clk,x41, x41_0_1 );
 Register22Bit Reg1 (clk,x41_0_1, y50 );
 Register22Bit Reg2 (clk,x41, x41_1_1 );
 Register22Bit Reg3 (clk,x41_1_1, y68 );

 Subtractor18Bit Sub2(clk, {x1[14],x1[14],x1[14], x1[14: 0] },  { x0[11: 0], 6'b0 },x10); 

 Register19Bit Reg4 (clk,x10, x10_0_1 );
 Register19Bit Reg5 (clk,x10_0_1, x10_0_2 );
 Register21Bit Reg6 (clk, {x10_0_2, 2'b0}, y3 );
 Register19Bit Reg7 (clk,x10, x10_1_1 );
 Register19Bit Reg8 (clk,x10_1_1, x10_1_2 );
 Register21Bit Reg9 (clk, {x10_1_2, 2'b0}, y20 );
 Register19Bit Reg10 (clk,x10, x10_2_1 );
 Register19Bit Reg11 (clk,x10_2_1, x10_2_2 );
 Register21Bit Reg12 (clk, {x10_2_2, 2'b0}, y98 );
 Register19Bit Reg13 (clk,x10, x10_3_1 );
 Register19Bit Reg14 (clk,x10_3_1, x10_3_2 );
 Register21Bit Reg15 (clk, {x10_3_2, 2'b0}, y115 );

 Subtractor22Bit Sub3(clk, {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] },  { x1[14: 0], 7'b0 },x11); 


 Adder23Bit Adder1(clk,  {x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0], 3'b0 }, { x11[22: 0]  }, x45); 

 Negator24Bit Neg0(clk, x45, x76 );
 Register24Bit Reg16 (clk,x76, y22 );
 Register24Bit Reg17 (clk,x76, y96 );

 Adder17Bit Adder2(clk,  { x0[11: 0], 5'b0 }, {x1[14],x1[14], x1[14: 0]  }, x12); 


 Adder20Bit Adder3(clk,  {x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0] },  { x1[14: 0], 5'b0 },x13); 

 Register21Bit Reg18 (clk,x13, x13_1_1 );
 Register21Bit Reg19 (clk,x13_1_1, x13_1_2 );
 Register22Bit Reg20 (clk, {x13_1_2, 1'b0}, y11 );
 Register21Bit Reg21 (clk,x13, x13_2_1 );
 Register21Bit Reg22 (clk,x13_2_1, x13_2_2 );
 Register22Bit Reg23 (clk, {x13_2_2, 1'b0}, y107 );

 Adder24Bit Adder4(clk,  {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] },  { x1[14: 0], 9'b0 },x17); 


 Subtractor20Bit Sub4(clk, {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] },  { x1[14: 0], 5'b0 },x18); 

 Register21Bit Reg24 (clk,x18, x18_0_1 );
 Register21Bit Reg25 (clk,x18_0_1, x18_0_2 );
 Register21Bit Reg26 (clk,x18_0_2, y9 );
 Register21Bit Reg27 (clk,x18, x18_1_1 );
 Register21Bit Reg28 (clk,x18_1_1, x18_1_2 );
 Register21Bit Reg29 (clk,x18_1_2, y109 );

 Adder21Bit Adder5(clk,  { x0[11: 0], 9'b0 }, {x1[14],x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0]  }, x19); 


 Subtractor22Bit Sub5(clk, { x19[21: 0] },  {x1[14],x1[14],x1[14], x1[14: 0], 4'b0 },x46); 

 Register23Bit Reg30 (clk,x46, x46_0_1 );
 Register23Bit Reg31 (clk,x46_0_1, y26 );
 Register23Bit Reg32 (clk,x46, x46_1_1 );
 Register23Bit Reg33 (clk,x46_1_1, y92 );

 Adder23Bit Adder6(clk,  {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] },  { x1[14: 0], 8'b0 },x20); 


 Subtractor24Bit Sub6(clk, {x5[16],x5[16],x5[16],x5[16],x5[16], x5[16: 0], 2'b0 }, { x20[23: 0] }, x63); 

 Register25Bit Reg34 (clk,x63, x63_0_1 );
 Register25Bit Reg35 (clk,x63_0_1, y45 );
 Register25Bit Reg36 (clk,x63, x63_1_1 );
 Register25Bit Reg37 (clk,x63_1_1, y73 );

 Subtractor22Bit Sub7(clk, {x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0] },  { x0[11: 0], 10'b0 },x21); 

 Register23Bit Reg38 (clk,x21, x21_0_1 );
 Register23Bit Reg39 (clk,x21_0_1, x21_0_2 );
 Register23Bit Reg40 (clk,x21_0_2, y46 );
 Register23Bit Reg41 (clk,x21, x21_1_1 );
 Register23Bit Reg42 (clk,x21_1_1, x21_1_2 );
 Register23Bit Reg43 (clk,x21_1_2, y72 );

 Subtractor16Bit Sub8(clk, { x0[11: 0], 4'b0 }, {x1[14], x1[14: 0] }, x22); 


 Adder24Bit Adder7(clk,  { x12[17: 0], 6'b0 }, {x22[16],x22[16],x22[16],x22[16],x22[16],x22[16],x22[16], x22[16: 0]  }, x65); 

 Register25Bit Reg44 (clk,x65, x65_0_1 );
 Register25Bit Reg45 (clk,x65_0_1, y54 );
 Register25Bit Reg46 (clk,x65, x65_1_1 );
 Register25Bit Reg47 (clk,x65_1_1, y64 );

 Subtractor20Bit Sub9(clk, { x1[14: 0], 5'b0 }, {x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0] }, x33); 

 Register21Bit Reg48 (clk,x33, x33_0_1 );
 Register21Bit Reg49 (clk,x33_0_1, x33_0_2 );
 Register23Bit Reg50 (clk, {x33_0_2, 2'b0}, y29 );
 Register21Bit Reg51 (clk,x33, x33_1_1 );
 Register21Bit Reg52 (clk,x33_1_1, x33_1_2 );
 Register23Bit Reg53 (clk, {x33_1_2, 2'b0}, y89 );

 Adder21Bit Adder8(clk,  {x1[14],x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0] },  { x1[14: 0], 6'b0 },x34); 


 Subtractor25Bit Sub10(clk, {x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0] },  { x1[14: 0], 10'b0 },x35); 

 Negator15Bit Neg1(clk, x1, x77 );
 Register15Bit Reg54 (clk,x77, x77_0_1 );
 Register15Bit Reg55 (clk,x77_0_1, x77_0_2 );
 Register21Bit Reg56 (clk, {x77_0_2, 6'b0}, y27 );
 Register15Bit Reg57 (clk,x77, x77_1_1 );
 Register15Bit Reg58 (clk,x77_1_1, x77_1_2 );
 Register21Bit Reg59 (clk, {x77_1_2, 6'b0}, y91 );
 Register15Bit Reg60 (clk,x1, x1_31_1 );
 Register15Bit Reg61 (clk,x1_31_1, x1_31_2 );
 Register15Bit Reg62 (clk,x1_31_2, x1_31_3 );
 Register17Bit Reg63 (clk, {x1_31_3, 2'b0}, y25 );
 Register15Bit Reg64 (clk,x1, x1_32_1 );
 Register15Bit Reg65 (clk,x1_32_1, x1_32_2 );
 Register15Bit Reg66 (clk,x1_32_2, x1_32_3 );
 Register17Bit Reg67 (clk, {x1_32_3, 2'b0}, y93 );

 Adder14Bit Adder9(clk,  {x0[11],x0[11], x0[11: 0] },  { x0[11: 0], 2'b0 },x2); 


 Subtractor19Bit Sub11(clk, { x1[14: 0], 4'b0 }, {x2[14],x2[14],x2[14],x2[14], x2[14: 0] }, x6); 


 Subtractor22Bit Sub12(clk, { x6[19: 0], 2'b0 }, {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] }, x31); 

 Register23Bit Reg68 (clk,x31, x31_0_1 );
 Register24Bit Reg69 (clk, {x31_0_1, 1'b0}, y15 );
 Register23Bit Reg70 (clk,x31, x31_1_1 );
 Register24Bit Reg71 (clk, {x31_1_1, 1'b0}, y103 );

 Adder23Bit Adder10(clk,  { x2[14: 0], 8'b0 }, {x6[19],x6[19],x6[19], x6[19: 0]  }, x51); 

 Negator24Bit Neg2(clk, x51, x87 );
 Register26Bit Reg72 (clk, {x87, 2'b0}, y56 );
 Register26Bit Reg73 (clk, {x87, 2'b0}, y62 );
 Register20Bit Reg74 (clk,x6, x6_3_1 );
 Register20Bit Reg75 (clk,x6_3_1, x6_3_2 );
 Register23Bit Reg76 (clk, {x6_3_2, 3'b0}, y36 );
 Register20Bit Reg77 (clk,x6, x6_4_1 );
 Register20Bit Reg78 (clk,x6_4_1, x6_4_2 );
 Register23Bit Reg79 (clk, {x6_4_2, 3'b0}, y82 );

 Subtractor17Bit Sub13(clk, { x0[11: 0], 5'b0 }, {x2[14],x2[14], x2[14: 0] }, x8); 


 Adder23Bit Adder11(clk,  {x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0] },  { x8[17: 0], 5'b0 },x44); 

 Register24Bit Reg80 (clk,x44, x44_0_1 );
 Register24Bit Reg81 (clk,x44_0_1, y40 );
 Register24Bit Reg82 (clk,x44, x44_1_1 );
 Register24Bit Reg83 (clk,x44_1_1, y78 );
 Negator18Bit Neg3(clk, x8, x78 );
 Register18Bit Reg84 (clk,x78, x78_0_1 );
 Register22Bit Reg85 (clk, {x78_0_1, 4'b0}, y28 );
 Register18Bit Reg86 (clk,x78, x78_1_1 );
 Register22Bit Reg87 (clk, {x78_1_1, 4'b0}, y90 );
 Register18Bit Reg88 (clk,x8, x8_2_1 );
 Register18Bit Reg89 (clk,x8_2_1, x8_2_2 );
 Register20Bit Reg90 (clk, {x8_2_2, 2'b0}, y18 );
 Register18Bit Reg91 (clk,x8, x8_3_1 );
 Register18Bit Reg92 (clk,x8_3_1, x8_3_2 );
 Register20Bit Reg93 (clk, {x8_3_2, 2'b0}, y100 );

 Adder17Bit Adder12(clk,  { x0[11: 0], 5'b0 }, {x2[14],x2[14], x2[14: 0]  }, x23); 

 Register18Bit Reg94 (clk,x23, x23_0_1 );
 Register18Bit Reg95 (clk,x23_0_1, x23_0_2 );
 Register20Bit Reg96 (clk, {x23_0_2, 2'b0}, y5 );
 Register18Bit Reg97 (clk,x23, x23_1_1 );
 Register18Bit Reg98 (clk,x23_1_1, x23_1_2 );
 Register20Bit Reg99 (clk, {x23_1_2, 2'b0}, y113 );

 Subtractor18Bit Sub14(clk, {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] },  { x2[14: 0], 3'b0 },x24); 

 Register19Bit Reg100 (clk,x24, x24_0_1 );
 Register19Bit Reg101 (clk,x24_0_1, x24_0_2 );
 Register21Bit Reg102 (clk, {x24_0_2, 2'b0}, y14 );
 Register19Bit Reg103 (clk,x24, x24_1_1 );
 Register19Bit Reg104 (clk,x24_1_1, x24_1_2 );
 Register21Bit Reg105 (clk, {x24_1_2, 2'b0}, y104 );

 Adder19Bit Adder13(clk,  { x0[11: 0], 7'b0 }, {x2[14],x2[14],x2[14],x2[14], x2[14: 0]  }, x25); 

 Negator20Bit Neg4(clk, x25, x79 );
 Register20Bit Reg106 (clk,x79, x79_0_1 );
 Register22Bit Reg107 (clk, {x79_0_1, 2'b0}, y31 );
 Register20Bit Reg108 (clk,x79, x79_1_1 );
 Register22Bit Reg109 (clk, {x79_1_1, 2'b0}, y87 );

 Adder22Bit Adder14(clk,  { x0[11: 0], 10'b0 }, {x2[14],x2[14],x2[14],x2[14],x2[14],x2[14],x2[14], x2[14: 0]  }, x26); 


 Adder23Bit Adder15(clk,  {x2[14],x2[14],x2[14],x2[14], x2[14: 0], 4'b0 }, { x26[22: 0]  }, x58); 

 Register24Bit Reg110 (clk,x58, x58_0_1 );
 Register24Bit Reg111 (clk,x58_0_1, y44 );
 Register24Bit Reg112 (clk,x58, x58_1_1 );
 Register24Bit Reg113 (clk,x58_1_1, y74 );

 Subtractor23Bit Sub15(clk, { x1[14: 0], 8'b0 }, {x2[14],x2[14],x2[14],x2[14],x2[14],x2[14],x2[14],x2[14], x2[14: 0] }, x36); 

 Register24Bit Reg114 (clk,x36, x36_0_1 );
 Register24Bit Reg115 (clk,x36_0_1, x36_0_2 );
 Register24Bit Reg116 (clk,x36_0_2, y4 );
 Register24Bit Reg117 (clk,x36, x36_1_1 );
 Register24Bit Reg118 (clk,x36_1_1, x36_1_2 );
 Register24Bit Reg119 (clk,x36_1_2, y114 );

 Subtractor20Bit Sub16(clk, {x2[14],x2[14],x2[14],x2[14],x2[14], x2[14: 0] },  { x1[14: 0], 5'b0 },x37); 

 Negator21Bit Neg5(clk, x37, x84 );
 Register21Bit Reg120 (clk,x84, x84_0_1 );
 Register24Bit Reg121 (clk, {x84_0_1, 3'b0}, y48 );
 Register21Bit Reg122 (clk,x84, x84_1_1 );
 Register24Bit Reg123 (clk, {x84_1_1, 3'b0}, y70 );

 Adder20Bit Adder16(clk,  {x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0] },  { x2[14: 0], 5'b0 },x38); 

 Register21Bit Reg124 (clk,x38, x38_0_1 );
 Register21Bit Reg125 (clk,x38_0_1, x38_0_2 );
 Register22Bit Reg126 (clk, {x38_0_2, 1'b0}, y30 );
 Register21Bit Reg127 (clk,x38, x38_1_1 );
 Register21Bit Reg128 (clk,x38_1_1, x38_1_2 );
 Register22Bit Reg129 (clk, {x38_1_2, 1'b0}, y88 );

 Adder20Bit Adder17(clk,  {x2[14],x2[14],x2[14],x2[14],x2[14], x2[14: 0] },  { x2[14: 0], 5'b0 },x47); 

 Register21Bit Reg130 (clk,x47, x47_0_1 );
 Register21Bit Reg131 (clk,x47_0_1, x47_0_2 );
 Register21Bit Reg132 (clk,x47_0_2, y41 );
 Register21Bit Reg133 (clk,x47, x47_1_1 );
 Register21Bit Reg134 (clk,x47_1_1, x47_1_2 );
 Register21Bit Reg135 (clk,x47_1_2, y77 );

 Adder22Bit Adder18(clk,  {x2[14],x2[14],x2[14],x2[14],x2[14],x2[14],x2[14], x2[14: 0] },  { x5[16: 0], 5'b0 },x49); 

 Register23Bit Reg136 (clk,x49, x49_0_1 );
 Register23Bit Reg137 (clk,x49_0_1, y37 );
 Register23Bit Reg138 (clk,x49, x49_1_1 );
 Register23Bit Reg139 (clk,x49_1_1, y81 );

 Subtractor22Bit Sub17(clk, {x5[16],x5[16],x5[16],x5[16],x5[16], x5[16: 0] },  { x2[14: 0], 7'b0 },x50); 

 Register23Bit Reg140 (clk,x50, x50_0_1 );
 Register23Bit Reg141 (clk,x50_0_1, y38 );
 Register23Bit Reg142 (clk,x50, x50_1_1 );
 Register23Bit Reg143 (clk,x50_1_1, y80 );

 Adder23Bit Adder19(clk,  {x2[14],x2[14],x2[14],x2[14],x2[14],x2[14], x2[14: 0], 2'b0 }, { x11[22: 0]  }, x52); 

 Register24Bit Reg144 (clk,x52, x52_0_1 );
 Register24Bit Reg145 (clk,x52_0_1, y17 );
 Register24Bit Reg146 (clk,x52, x52_1_1 );
 Register24Bit Reg147 (clk,x52_1_1, y101 );

 Adder22Bit Adder20(clk,  { x2[14: 0], 7'b0 }, {x12[17],x12[17],x12[17],x12[17], x12[17: 0]  }, x53); 

 Negator23Bit Neg6(clk, x53, x82 );
 Register23Bit Reg148 (clk,x82, y35 );
 Register23Bit Reg149 (clk,x82, y83 );

 Adder25Bit Adder21(clk,  {x2[14],x2[14],x2[14],x2[14],x2[14],x2[14],x2[14],x2[14],x2[14],x2[14], x2[14: 0] },  { x13[20: 0], 4'b0 },x54); 

 Negator26Bit Neg7(clk, x54, x72 );
 Register26Bit Reg150 (clk,x72, y1 );
 Register26Bit Reg151 (clk,x72, y117 );

 Adder25Bit Adder22(clk,  {x2[14],x2[14],x2[14],x2[14],x2[14],x2[14],x2[14], x2[14: 0], 3'b0 }, { x17[24: 0]  }, x57); 

 Negator26Bit Neg8(clk, x57, x73 );
 Register26Bit Reg152 (clk,x73, y2 );
 Register26Bit Reg153 (clk,x73, y116 );

 Adder26Bit Adder23(clk,  {x2[14],x2[14],x2[14],x2[14],x2[14],x2[14],x2[14],x2[14],x2[14],x2[14],x2[14], x2[14: 0] },  { x34[21: 0], 4'b0 },x59); 

 Register27Bit Reg154 (clk,x59, x59_0_1 );
 Register27Bit Reg155 (clk,x59_0_1, y55 );
 Register27Bit Reg156 (clk,x59, x59_1_1 );
 Register27Bit Reg157 (clk,x59_1_1, y63 );
 Register15Bit Reg158 (clk,x2, x2_23_1 );
 Register15Bit Reg159 (clk,x2_23_1, x2_23_2 );
 Register15Bit Reg160 (clk,x2_23_2, x2_23_3 );
 Register22Bit Reg161 (clk, {x2_23_3, 7'b0}, y33 );
 Register15Bit Reg162 (clk,x2, x2_24_1 );
 Register15Bit Reg163 (clk,x2_24_1, x2_24_2 );
 Register15Bit Reg164 (clk,x2_24_2, x2_24_3 );
 Register22Bit Reg165 (clk, {x2_24_3, 7'b0}, y85 );

 Adder15Bit Adder24(clk,  {x0[11],x0[11],x0[11], x0[11: 0] },  { x0[11: 0], 3'b0 },x3); 


 Adder20Bit Adder25(clk,  { x0[11: 0], 8'b0 }, {x3[15],x3[15],x3[15],x3[15], x3[15: 0]  }, x9); 

 Negator21Bit Neg9(clk, x9, x74 );
 Register21Bit Reg166 (clk,x74, x74_0_1 );
 Register22Bit Reg167 (clk, {x74_0_1, 1'b0}, y6 );
 Register21Bit Reg168 (clk,x74, x74_1_1 );
 Register21Bit Reg169 (clk,x74_1_1, y21 );
 Register21Bit Reg170 (clk,x74, x74_2_1 );
 Register21Bit Reg171 (clk,x74_2_1, y97 );
 Register21Bit Reg172 (clk,x74, x74_3_1 );
 Register22Bit Reg173 (clk, {x74_3_1, 1'b0}, y112 );
 Register21Bit Reg174 (clk,x9, x9_1_1 );
 Register21Bit Reg175 (clk,x9_1_1, x9_1_2 );
 Register21Bit Reg176 (clk,x9_1_2, y12 );
 Register21Bit Reg177 (clk,x9, x9_2_1 );
 Register21Bit Reg178 (clk,x9_2_1, x9_2_2 );
 Register21Bit Reg179 (clk,x9_2_2, y106 );

 Subtractor21Bit Sub18(clk, {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] },  { x3[15: 0], 5'b0 },x27); 

 Register22Bit Reg180 (clk,x27, x27_0_1 );
 Register22Bit Reg181 (clk,x27_0_1, x27_0_2 );
 Register22Bit Reg182 (clk,x27_0_2, y13 );
 Register22Bit Reg183 (clk,x27, x27_1_1 );
 Register22Bit Reg184 (clk,x27_1_1, x27_1_2 );
 Register22Bit Reg185 (clk,x27_1_2, y105 );

 Subtractor18Bit Sub19(clk, {x3[15],x3[15], x3[15: 0] },  { x0[11: 0], 6'b0 },x28); 

 Register19Bit Reg186 (clk,x28, x28_0_1 );
 Register19Bit Reg187 (clk,x28_0_1, x28_0_2 );
 Register22Bit Reg188 (clk, {x28_0_2, 3'b0}, y24 );
 Register19Bit Reg189 (clk,x28, x28_1_1 );
 Register19Bit Reg190 (clk,x28_1_1, x28_1_2 );
 Register22Bit Reg191 (clk, {x28_1_2, 3'b0}, y94 );

 Subtractor27Bit Sub20(clk, { x3[15: 0], 11'b0 }, {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] }, x29); 


 Subtractor28Bit Sub21(clk, { x29[27: 0] },  {x5[16],x5[16],x5[16],x5[16],x5[16],x5[16],x5[16],x5[16],x5[16], x5[16: 0], 2'b0 },x64); 

 Register29Bit Reg192 (clk,x64, x64_0_1 );
 Register29Bit Reg193 (clk,x64_0_1, y58 );
 Register29Bit Reg194 (clk,x64, x64_1_1 );
 Register29Bit Reg195 (clk,x64_1_1, y60 );

 Adder26Bit Adder26(clk,  {x3[15],x3[15],x3[15],x3[15],x3[15],x3[15],x3[15],x3[15],x3[15],x3[15], x3[15: 0] },  { x6[19: 0], 6'b0 },x61); 

 Negator27Bit Neg10(clk, x61, x86 );
 Register27Bit Reg196 (clk,x86, y53 );
 Register27Bit Reg197 (clk,x86, y65 );

 Subtractor26Bit Sub22(clk, { x35[25: 0] },  {x3[15],x3[15],x3[15],x3[15],x3[15], x3[15: 0], 5'b0 },x62); 

 Register27Bit Reg198 (clk,x62, x62_0_1 );
 Register27Bit Reg199 (clk,x62_0_1, y57 );
 Register27Bit Reg200 (clk,x62, x62_1_1 );
 Register27Bit Reg201 (clk,x62_1_1, y61 );
 Register16Bit Reg202 (clk,x3, x3_7_1 );
 Register16Bit Reg203 (clk,x3_7_1, x3_7_2 );
 Register16Bit Reg204 (clk,x3_7_2, x3_7_3 );
 Register20Bit Reg205 (clk, {x3_7_3, 4'b0}, y23 );
 Register16Bit Reg206 (clk,x3, x3_8_1 );
 Register16Bit Reg207 (clk,x3_8_1, x3_8_2 );
 Register16Bit Reg208 (clk,x3_8_2, x3_8_3 );
 Register20Bit Reg209 (clk, {x3_8_3, 4'b0}, y95 );

 Subtractor15Bit Sub23(clk, { x0[11: 0], 3'b0 }, {x0[11],x0[11],x0[11], x0[11: 0] }, x4); 


 Subtractor21Bit Sub24(clk, {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] },  { x4[15: 0], 5'b0 },x30); 

 Register22Bit Reg210 (clk,x30, x30_0_1 );
 Register22Bit Reg211 (clk,x30_0_1, x30_0_2 );
 Register23Bit Reg212 (clk, {x30_0_2, 1'b0}, y39 );
 Register22Bit Reg213 (clk,x30, x30_1_1 );
 Register22Bit Reg214 (clk,x30_1_1, x30_1_2 );
 Register23Bit Reg215 (clk, {x30_1_2, 1'b0}, y79 );

 Subtractor20Bit Sub25(clk, { x4[15: 0], 4'b0 }, {x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0] }, x39); 

 Register21Bit Reg216 (clk,x39, x39_0_1 );
 Register21Bit Reg217 (clk,x39_0_1, x39_0_2 );
 Register23Bit Reg218 (clk, {x39_0_2, 2'b0}, y8 );
 Register21Bit Reg219 (clk,x39, x39_1_1 );
 Register21Bit Reg220 (clk,x39_1_1, x39_1_2 );
 Register23Bit Reg221 (clk, {x39_1_2, 2'b0}, y110 );

 Subtractor21Bit Sub26(clk, {x1[14],x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0] },  { x4[15: 0], 5'b0 },x40); 

 Register22Bit Reg222 (clk,x40, x40_0_1 );
 Register22Bit Reg223 (clk,x40_0_1, x40_0_2 );
 Register25Bit Reg224 (clk, {x40_0_2, 3'b0}, y49 );
 Register22Bit Reg225 (clk,x40, x40_1_1 );
 Register22Bit Reg226 (clk,x40_1_1, x40_1_2 );
 Register25Bit Reg227 (clk, {x40_1_2, 3'b0}, y69 );

 Subtractor21Bit Sub27(clk, { x4[15: 0], 5'b0 }, {x2[14],x2[14],x2[14],x2[14],x2[14],x2[14], x2[14: 0] }, x48); 

 Register22Bit Reg228 (clk,x48, x48_0_1 );
 Register22Bit Reg229 (clk,x48_0_1, x48_0_2 );
 Register22Bit Reg230 (clk,x48_0_2, y43 );
 Register22Bit Reg231 (clk,x48, x48_1_1 );
 Register22Bit Reg232 (clk,x48_1_1, x48_1_2 );
 Register22Bit Reg233 (clk,x48_1_2, y75 );

 Subtractor24Bit Sub28(clk, { x3[15: 0], 8'b0 }, {x4[15],x4[15],x4[15],x4[15],x4[15],x4[15],x4[15],x4[15], x4[15: 0] }, x60); 

 Register25Bit Reg234 (clk,x60, x60_0_1 );
 Register25Bit Reg235 (clk,x60_0_1, x60_0_2 );
 Register25Bit Reg236 (clk,x60_0_2, y51 );
 Register25Bit Reg237 (clk,x60, x60_1_1 );
 Register25Bit Reg238 (clk,x60_1_1, x60_1_2 );
 Register25Bit Reg239 (clk,x60_1_2, y67 );
 Register16Bit Reg240 (clk,x4, x4_5_1 );
 Register16Bit Reg241 (clk,x4_5_1, x4_5_2 );
 Register16Bit Reg242 (clk,x4_5_2, x4_5_3 );
 Register18Bit Reg243 (clk, {x4_5_3, 2'b0}, y16 );
 Register16Bit Reg244 (clk,x4, x4_6_1 );
 Register16Bit Reg245 (clk,x4_6_1, x4_6_2 );
 Register16Bit Reg246 (clk,x4_6_2, x4_6_3 );
 Register18Bit Reg247 (clk, {x4_6_3, 2'b0}, y102 );

 Subtractor16Bit Sub29(clk, {x0[11],x0[11],x0[11],x0[11], x0[11: 0] },  { x0[11: 0], 4'b0 },x7); 


 Subtractor20Bit Sub30(clk, {x7[16],x7[16],x7[16], x7[16: 0] },  { x0[11: 0], 8'b0 },x32); 

 Register21Bit Reg248 (clk,x32, x32_0_1 );
 Register21Bit Reg249 (clk,x32_0_1, x32_0_2 );
 Register22Bit Reg250 (clk, {x32_0_2, 1'b0}, y0 );
 Register21Bit Reg251 (clk,x32, x32_1_1 );
 Register21Bit Reg252 (clk,x32_1_1, x32_1_2 );
 Register22Bit Reg253 (clk, {x32_1_2, 1'b0}, y118 );

 Adder21Bit Adder27(clk,  { x1[14: 0], 6'b0 }, {x7[16],x7[16],x7[16],x7[16], x7[16: 0]  }, x42); 

 Negator22Bit Neg11(clk, x42, x75 );
 Register22Bit Reg254 (clk,x75, x75_0_1 );
 Register23Bit Reg255 (clk, {x75_0_1, 1'b0}, y10 );
 Register22Bit Reg256 (clk,x75, x75_1_1 );
 Register23Bit Reg257 (clk, {x75_1_1, 1'b0}, y108 );

 Adder22Bit Adder28(clk,  { x1[14: 0], 7'b0 }, {x7[16],x7[16],x7[16],x7[16],x7[16], x7[16: 0]  }, x43); 

 Negator23Bit Neg12(clk, x43, x85 );
 Register23Bit Reg258 (clk,x85, x85_0_1 );
 Register24Bit Reg259 (clk, {x85_0_1, 1'b0}, y52 );
 Register23Bit Reg260 (clk,x85, x85_1_1 );
 Register24Bit Reg261 (clk, {x85_1_1, 1'b0}, y66 );

 Adder16Bit Adder29(clk,  {x0[11],x0[11],x0[11],x0[11], x0[11: 0] },  { x0[11: 0], 4'b0 },x14); 


 Adder21Bit Adder30(clk,  { x2[14: 0], 6'b0 }, {x14[16],x14[16],x14[16],x14[16], x14[16: 0]  }, x55); 

 Register22Bit Reg262 (clk,x55, x55_0_1 );
 Register22Bit Reg263 (clk,x55_0_1, x55_0_2 );
 Register22Bit Reg264 (clk,x55_0_2, y19 );
 Register22Bit Reg265 (clk,x55, x55_1_1 );
 Register22Bit Reg266 (clk,x55_1_1, x55_1_2 );
 Register22Bit Reg267 (clk,x55_1_2, y99 );

 Subtractor17Bit Sub31(clk, {x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] },  { x0[11: 0], 5'b0 },x15); 

 Register18Bit Reg268 (clk,x15, x15_0_1 );
 Register18Bit Reg269 (clk,x15_0_1, x15_0_2 );
 Register18Bit Reg270 (clk,x15_0_2, x15_0_3 );
 Register18Bit Reg271 (clk,x15_0_3, y7 );
 Register18Bit Reg272 (clk,x15, x15_1_1 );
 Register18Bit Reg273 (clk,x15_1_1, x15_1_2 );
 Register18Bit Reg274 (clk,x15_1_2, x15_1_3 );
 Register18Bit Reg275 (clk,x15_1_3, y111 );

 Adder22Bit Adder31(clk,  {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] },  { x0[11: 0], 10'b0 },x16); 


 Adder23Bit Adder32(clk,  {x2[14],x2[14],x2[14],x2[14],x2[14],x2[14], x2[14: 0], 2'b0 }, { x16[22: 0]  }, x56); 

 Negator24Bit Neg13(clk, x56, x83 );
 Register24Bit Reg276 (clk,x83, x83_0_1 );
 Register24Bit Reg277 (clk,x83_0_1, y42 );
 Register24Bit Reg278 (clk,x83, x83_1_1 );
 Register24Bit Reg279 (clk,x83_1_1, y76 );
 Register12Bit Reg280 (clk,x0, x66_38_1 );
 Register12Bit Reg281 (clk,x66_38_1, x66_38_2 );

 Adder19Bit Adder33(clk,  {x66_38_2[11],x66_38_2[11],x66_38_2[11],x66_38_2[11],x66_38_2[11],x66_38_2[11],x66_38_2[11], x66_38_2[11: 0] },  { x5[16: 0], 2'b0 },x66); 

 Negator20Bit Neg14(clk, x66, x80 );
 Register21Bit Reg282 (clk, {x80, 1'b0}, y32 );
 Register12Bit Reg283 (clk,x0, x67_39_1 );
 Register12Bit Reg284 (clk,x67_39_1, x67_39_2 );

 Adder19Bit Adder34(clk,  {x67_39_2[11],x67_39_2[11],x67_39_2[11],x67_39_2[11],x67_39_2[11],x67_39_2[11],x67_39_2[11], x67_39_2[11: 0] },  { x5[16: 0], 2'b0 },x67); 

 Negator20Bit Neg15(clk, x67, x81 );
 Register20Bit Reg285 (clk,x81, y34 );
 Register12Bit Reg286 (clk,x0, x68_40_1 );
 Register12Bit Reg287 (clk,x68_40_1, x68_40_2 );

 Adder21Bit Adder35(clk,  {x68_40_2[11],x68_40_2[11],x68_40_2[11],x68_40_2[11],x68_40_2[11],x68_40_2[11],x68_40_2[11],x68_40_2[11],x68_40_2[11], x68_40_2[11: 0] },  { x5[16: 0], 4'b0 },x68); 

 Register22Bit Reg288 (clk,x68, x68_0_1 );
 Register24Bit Reg289 (clk, {x68_0_1, 2'b0}, y47 );
 Register12Bit Reg290 (clk,x0, x69_41_1 );
 Register12Bit Reg291 (clk,x69_41_1, x69_41_2 );

 Adder21Bit Adder36(clk,  {x69_41_2[11],x69_41_2[11],x69_41_2[11],x69_41_2[11],x69_41_2[11],x69_41_2[11],x69_41_2[11],x69_41_2[11],x69_41_2[11], x69_41_2[11: 0] },  { x5[16: 0], 4'b0 },x69); 

 Register22Bit Reg292 (clk,x69, x69_0_1 );
 Register24Bit Reg293 (clk, {x69_0_1, 2'b0}, y71 );
 Register12Bit Reg294 (clk,x0, x70_42_1 );
 Register12Bit Reg295 (clk,x70_42_1, x70_42_2 );

 Adder19Bit Adder37(clk,  {x70_42_2[11],x70_42_2[11],x70_42_2[11],x70_42_2[11],x70_42_2[11],x70_42_2[11],x70_42_2[11], x70_42_2[11: 0] },  { x5[16: 0], 2'b0 },x70); 

 Negator20Bit Neg16(clk, x70, x88 );
 Register20Bit Reg296 (clk,x88, y84 );
 Register12Bit Reg297 (clk,x0, x71_43_1 );
 Register12Bit Reg298 (clk,x71_43_1, x71_43_2 );

 Adder19Bit Adder38(clk,  {x71_43_2[11],x71_43_2[11],x71_43_2[11],x71_43_2[11],x71_43_2[11],x71_43_2[11],x71_43_2[11], x71_43_2[11: 0] },  { x5[16: 0], 2'b0 },x71); 

 Negator20Bit Neg17(clk, x71, x89 );
 Register21Bit Reg299 (clk, {x89, 1'b0}, y86 );
 Register12Bit Reg300 (clk,x0, x0_44_1 );
 Register12Bit Reg301 (clk,x0_44_1, x0_44_2 );
 Register12Bit Reg302 (clk,x0_44_2, x0_44_3 );
 Register12Bit Reg303 (clk,x0_44_3, x0_44_4 );
 Register27Bit Reg304 (clk, {x0_44_4, 15'b0}, y59 );
 Register22Bit Reg305 (clk,y0, x90 );

 Adder26Bit Adder39(clk,  {x90[21],x90[21],x90[21],x90[21], x90[21: 0] },  { y1[25: 0]  }, x91); 

 Register27Bit Reg306 (clk,x91, x91_1 );

 Adder27Bit Adder40(clk,  { x91_1[26: 0] },  {y2[25], y2[25: 0]  }, x92); 

 Register28Bit Reg307 (clk,x92, x92_1 );

 Adder28Bit Adder41(clk,  { x92_1[27: 0] },  {y3[20],y3[20],y3[20],y3[20],y3[20],y3[20],y3[20], y3[20: 0]  }, x93); 

 Register29Bit Reg308 (clk,x93, x93_1 );

 Adder29Bit Adder42(clk,  { x93_1[28: 0] },  {y4[23],y4[23],y4[23],y4[23],y4[23], y4[23: 0]  }, x94); 

 Register29Bit Reg309 (clk,x94, x94_1 );

 Adder29Bit Adder43(clk,  { x94_1[28: 0] },  {y5[19],y5[19],y5[19],y5[19],y5[19],y5[19],y5[19],y5[19],y5[19], y5[19: 0]  }, x95); 

 Register29Bit Reg310 (clk,x95, x95_1 );

 Adder29Bit Adder44(clk,  { x95_1[28: 0] },  {y6[21],y6[21],y6[21],y6[21],y6[21],y6[21],y6[21], y6[21: 0]  }, x96); 

 Register29Bit Reg311 (clk,x96, x96_1 );

 Adder29Bit Adder45(clk,  { x96_1[28: 0] },  {y7[17],y7[17],y7[17],y7[17],y7[17],y7[17],y7[17],y7[17],y7[17],y7[17],y7[17], y7[17: 0]  }, x97); 

 Register29Bit Reg312 (clk,x97, x97_1 );

 Adder29Bit Adder46(clk,  { x97_1[28: 0] },  {y8[22],y8[22],y8[22],y8[22],y8[22],y8[22], y8[22: 0]  }, x98); 

 Register29Bit Reg313 (clk,x98, x98_1 );

 Adder29Bit Adder47(clk,  { x98_1[28: 0] },  {y9[20],y9[20],y9[20],y9[20],y9[20],y9[20],y9[20],y9[20], y9[20: 0]  }, x99); 

 Register29Bit Reg314 (clk,x99, x99_1 );

 Adder29Bit Adder48(clk,  { x99_1[28: 0] },  {y10[22],y10[22],y10[22],y10[22],y10[22],y10[22], y10[22: 0]  }, x100); 

 Register29Bit Reg315 (clk,x100, x100_1 );

 Adder29Bit Adder49(clk,  { x100_1[28: 0] },  {y11[21],y11[21],y11[21],y11[21],y11[21],y11[21],y11[21], y11[21: 0]  }, x101); 

 Register29Bit Reg316 (clk,x101, x101_1 );

 Adder29Bit Adder50(clk,  { x101_1[28: 0] },  {y12[20],y12[20],y12[20],y12[20],y12[20],y12[20],y12[20],y12[20], y12[20: 0]  }, x102); 

 Register29Bit Reg317 (clk,x102, x102_1 );

 Adder29Bit Adder51(clk,  { x102_1[28: 0] },  {y13[21],y13[21],y13[21],y13[21],y13[21],y13[21],y13[21], y13[21: 0]  }, x103); 

 Register29Bit Reg318 (clk,x103, x103_1 );

 Adder29Bit Adder52(clk,  { x103_1[28: 0] },  {y14[20],y14[20],y14[20],y14[20],y14[20],y14[20],y14[20],y14[20], y14[20: 0]  }, x104); 

 Register29Bit Reg319 (clk,x104, x104_1 );

 Adder29Bit Adder53(clk,  { x104_1[28: 0] },  {y15[23],y15[23],y15[23],y15[23],y15[23], y15[23: 0]  }, x105); 

 Register29Bit Reg320 (clk,x105, x105_1 );

 Adder29Bit Adder54(clk,  { x105_1[28: 0] },  {y16[17],y16[17],y16[17],y16[17],y16[17],y16[17],y16[17],y16[17],y16[17],y16[17],y16[17], y16[17: 0]  }, x106); 

 Register29Bit Reg321 (clk,x106, x106_1 );

 Adder29Bit Adder55(clk,  { x106_1[28: 0] },  {y17[23],y17[23],y17[23],y17[23],y17[23], y17[23: 0]  }, x107); 

 Register29Bit Reg322 (clk,x107, x107_1 );

 Adder29Bit Adder56(clk,  { x107_1[28: 0] },  {y18[19],y18[19],y18[19],y18[19],y18[19],y18[19],y18[19],y18[19],y18[19], y18[19: 0]  }, x108); 

 Register29Bit Reg323 (clk,x108, x108_1 );

 Adder29Bit Adder57(clk,  { x108_1[28: 0] },  {y19[21],y19[21],y19[21],y19[21],y19[21],y19[21],y19[21], y19[21: 0]  }, x109); 

 Register29Bit Reg324 (clk,x109, x109_1 );

 Adder29Bit Adder58(clk,  { x109_1[28: 0] },  {y20[20],y20[20],y20[20],y20[20],y20[20],y20[20],y20[20],y20[20], y20[20: 0]  }, x110); 

 Register29Bit Reg325 (clk,x110, x110_1 );

 Adder29Bit Adder59(clk,  { x110_1[28: 0] },  {y21[20],y21[20],y21[20],y21[20],y21[20],y21[20],y21[20],y21[20], y21[20: 0]  }, x111); 

 Register29Bit Reg326 (clk,x111, x111_1 );

 Adder29Bit Adder60(clk,  { x111_1[28: 0] },  {y22[23],y22[23],y22[23],y22[23],y22[23], y22[23: 0]  }, x112); 

 Register29Bit Reg327 (clk,x112, x112_1 );

 Adder29Bit Adder61(clk,  { x112_1[28: 0] },  {y23[19],y23[19],y23[19],y23[19],y23[19],y23[19],y23[19],y23[19],y23[19], y23[19: 0]  }, x113); 

 Register29Bit Reg328 (clk,x113, x113_1 );

 Adder29Bit Adder62(clk,  { x113_1[28: 0] },  {y24[21],y24[21],y24[21],y24[21],y24[21],y24[21],y24[21], y24[21: 0]  }, x114); 

 Register29Bit Reg329 (clk,x114, x114_1 );

 Adder29Bit Adder63(clk,  { x114_1[28: 0] },  {y25[16],y25[16],y25[16],y25[16],y25[16],y25[16],y25[16],y25[16],y25[16],y25[16],y25[16],y25[16], y25[16: 0]  }, x115); 

 Register29Bit Reg330 (clk,x115, x115_1 );

 Adder29Bit Adder64(clk,  { x115_1[28: 0] },  {y26[22],y26[22],y26[22],y26[22],y26[22],y26[22], y26[22: 0]  }, x116); 

 Register29Bit Reg331 (clk,x116, x116_1 );

 Adder29Bit Adder65(clk,  { x116_1[28: 0] },  {y27[20],y27[20],y27[20],y27[20],y27[20],y27[20],y27[20],y27[20], y27[20: 0]  }, x117); 

 Register29Bit Reg332 (clk,x117, x117_1 );

 Adder29Bit Adder66(clk,  { x117_1[28: 0] },  {y28[21],y28[21],y28[21],y28[21],y28[21],y28[21],y28[21], y28[21: 0]  }, x118); 

 Register29Bit Reg333 (clk,x118, x118_1 );

 Adder29Bit Adder67(clk,  { x118_1[28: 0] },  {y29[22],y29[22],y29[22],y29[22],y29[22],y29[22], y29[22: 0]  }, x119); 

 Register29Bit Reg334 (clk,x119, x119_1 );

 Adder29Bit Adder68(clk,  { x119_1[28: 0] },  {y30[21],y30[21],y30[21],y30[21],y30[21],y30[21],y30[21], y30[21: 0]  }, x120); 

 Register29Bit Reg335 (clk,x120, x120_1 );

 Adder29Bit Adder69(clk,  { x120_1[28: 0] },  {y31[21],y31[21],y31[21],y31[21],y31[21],y31[21],y31[21], y31[21: 0]  }, x121); 

 Register29Bit Reg336 (clk,x121, x121_1 );

 Adder29Bit Adder70(clk,  { x121_1[28: 0] },  {y32[20],y32[20],y32[20],y32[20],y32[20],y32[20],y32[20],y32[20], y32[20: 0]  }, x122); 

 Register29Bit Reg337 (clk,x122, x122_1 );

 Adder29Bit Adder71(clk,  { x122_1[28: 0] },  {y33[21],y33[21],y33[21],y33[21],y33[21],y33[21],y33[21], y33[21: 0]  }, x123); 

 Register29Bit Reg338 (clk,x123, x123_1 );

 Adder29Bit Adder72(clk,  { x123_1[28: 0] },  {y34[19],y34[19],y34[19],y34[19],y34[19],y34[19],y34[19],y34[19],y34[19], y34[19: 0]  }, x124); 

 Register29Bit Reg339 (clk,x124, x124_1 );

 Adder29Bit Adder73(clk,  { x124_1[28: 0] },  {y35[22],y35[22],y35[22],y35[22],y35[22],y35[22], y35[22: 0]  }, x125); 

 Register29Bit Reg340 (clk,x125, x125_1 );

 Adder29Bit Adder74(clk,  { x125_1[28: 0] },  {y36[22],y36[22],y36[22],y36[22],y36[22],y36[22], y36[22: 0]  }, x126); 

 Register29Bit Reg341 (clk,x126, x126_1 );

 Adder29Bit Adder75(clk,  { x126_1[28: 0] },  {y37[22],y37[22],y37[22],y37[22],y37[22],y37[22], y37[22: 0]  }, x127); 

 Register29Bit Reg342 (clk,x127, x127_1 );

 Adder29Bit Adder76(clk,  { x127_1[28: 0] },  {y38[22],y38[22],y38[22],y38[22],y38[22],y38[22], y38[22: 0]  }, x128); 

 Register29Bit Reg343 (clk,x128, x128_1 );

 Adder29Bit Adder77(clk,  { x128_1[28: 0] },  {y39[22],y39[22],y39[22],y39[22],y39[22],y39[22], y39[22: 0]  }, x129); 

 Register29Bit Reg344 (clk,x129, x129_1 );

 Adder29Bit Adder78(clk,  { x129_1[28: 0] },  {y40[23],y40[23],y40[23],y40[23],y40[23], y40[23: 0]  }, x130); 

 Register29Bit Reg345 (clk,x130, x130_1 );

 Adder29Bit Adder79(clk,  { x130_1[28: 0] },  {y41[20],y41[20],y41[20],y41[20],y41[20],y41[20],y41[20],y41[20], y41[20: 0]  }, x131); 

 Register29Bit Reg346 (clk,x131, x131_1 );

 Adder29Bit Adder80(clk,  { x131_1[28: 0] },  {y42[23],y42[23],y42[23],y42[23],y42[23], y42[23: 0]  }, x132); 

 Register29Bit Reg347 (clk,x132, x132_1 );

 Adder29Bit Adder81(clk,  { x132_1[28: 0] },  {y43[21],y43[21],y43[21],y43[21],y43[21],y43[21],y43[21], y43[21: 0]  }, x133); 

 Register29Bit Reg348 (clk,x133, x133_1 );

 Adder29Bit Adder82(clk,  { x133_1[28: 0] },  {y44[23],y44[23],y44[23],y44[23],y44[23], y44[23: 0]  }, x134); 

 Register29Bit Reg349 (clk,x134, x134_1 );

 Adder29Bit Adder83(clk,  { x134_1[28: 0] },  {y45[24],y45[24],y45[24],y45[24], y45[24: 0]  }, x135); 

 Register29Bit Reg350 (clk,x135, x135_1 );

 Adder29Bit Adder84(clk,  { x135_1[28: 0] },  {y46[22],y46[22],y46[22],y46[22],y46[22],y46[22], y46[22: 0]  }, x136); 

 Register29Bit Reg351 (clk,x136, x136_1 );

 Adder29Bit Adder85(clk,  { x136_1[28: 0] },  {y47[23],y47[23],y47[23],y47[23],y47[23], y47[23: 0]  }, x137); 

 Register29Bit Reg352 (clk,x137, x137_1 );

 Adder29Bit Adder86(clk,  { x137_1[28: 0] },  {y48[23],y48[23],y48[23],y48[23],y48[23], y48[23: 0]  }, x138); 

 Register29Bit Reg353 (clk,x138, x138_1 );

 Adder29Bit Adder87(clk,  { x138_1[28: 0] },  {y49[24],y49[24],y49[24],y49[24], y49[24: 0]  }, x139); 

 Register29Bit Reg354 (clk,x139, x139_1 );

 Adder29Bit Adder88(clk,  { x139_1[28: 0] },  {y50[21],y50[21],y50[21],y50[21],y50[21],y50[21],y50[21], y50[21: 0]  }, x140); 

 Register29Bit Reg355 (clk,x140, x140_1 );

 Adder29Bit Adder89(clk,  { x140_1[28: 0] },  {y51[24],y51[24],y51[24],y51[24], y51[24: 0]  }, x141); 

 Register29Bit Reg356 (clk,x141, x141_1 );

 Adder29Bit Adder90(clk,  { x141_1[28: 0] },  {y52[23],y52[23],y52[23],y52[23],y52[23], y52[23: 0]  }, x142); 

 Register29Bit Reg357 (clk,x142, x142_1 );

 Adder29Bit Adder91(clk,  { x142_1[28: 0] },  {y53[26],y53[26], y53[26: 0]  }, x143); 

 Register29Bit Reg358 (clk,x143, x143_1 );

 Adder29Bit Adder92(clk,  { x143_1[28: 0] },  {y54[24],y54[24],y54[24],y54[24], y54[24: 0]  }, x144); 

 Register29Bit Reg359 (clk,x144, x144_1 );

 Adder29Bit Adder93(clk,  { x144_1[28: 0] },  {y55[26],y55[26], y55[26: 0]  }, x145); 

 Register29Bit Reg360 (clk,x145, x145_1 );

 Adder29Bit Adder94(clk,  { x145_1[28: 0] },  {y56[25],y56[25],y56[25], y56[25: 0]  }, x146); 

 Register29Bit Reg361 (clk,x146, x146_1 );

 Adder29Bit Adder95(clk,  { x146_1[28: 0] },  {y57[26],y57[26], y57[26: 0]  }, x147); 

 Register29Bit Reg362 (clk,x147, x147_1 );

 Adder29Bit Adder96(clk,  { x147_1[28: 0] },  { y58[28: 0]  }, x148); 

 Register29Bit Reg363 (clk,x148, x148_1 );

 Adder29Bit Adder97(clk,  { x148_1[28: 0] },  {y59[26],y59[26], y59[26: 0]  }, x149); 

 Register29Bit Reg364 (clk,x149, x149_1 );

 Adder29Bit Adder98(clk,  { x149_1[28: 0] },  { y60[28: 0]  }, x150); 

 Register29Bit Reg365 (clk,x150, x150_1 );

 Adder29Bit Adder99(clk,  { x150_1[28: 0] },  {y61[26],y61[26], y61[26: 0]  }, x151); 

 Register29Bit Reg366 (clk,x151, x151_1 );

 Adder29Bit Adder100(clk,  { x151_1[28: 0] },  {y62[25],y62[25],y62[25], y62[25: 0]  }, x152); 

 Register29Bit Reg367 (clk,x152, x152_1 );

 Adder29Bit Adder101(clk,  { x152_1[28: 0] },  {y63[26],y63[26], y63[26: 0]  }, x153); 

 Register29Bit Reg368 (clk,x153, x153_1 );

 Adder29Bit Adder102(clk,  { x153_1[28: 0] },  {y64[24],y64[24],y64[24],y64[24], y64[24: 0]  }, x154); 

 Register29Bit Reg369 (clk,x154, x154_1 );

 Adder29Bit Adder103(clk,  { x154_1[28: 0] },  {y65[26],y65[26], y65[26: 0]  }, x155); 

 Register29Bit Reg370 (clk,x155, x155_1 );

 Adder29Bit Adder104(clk,  { x155_1[28: 0] },  {y66[23],y66[23],y66[23],y66[23],y66[23], y66[23: 0]  }, x156); 

 Register29Bit Reg371 (clk,x156, x156_1 );

 Adder29Bit Adder105(clk,  { x156_1[28: 0] },  {y67[24],y67[24],y67[24],y67[24], y67[24: 0]  }, x157); 

 Register29Bit Reg372 (clk,x157, x157_1 );

 Adder29Bit Adder106(clk,  { x157_1[28: 0] },  {y68[21],y68[21],y68[21],y68[21],y68[21],y68[21],y68[21], y68[21: 0]  }, x158); 

 Register29Bit Reg373 (clk,x158, x158_1 );

 Adder29Bit Adder107(clk,  { x158_1[28: 0] },  {y69[24],y69[24],y69[24],y69[24], y69[24: 0]  }, x159); 

 Register29Bit Reg374 (clk,x159, x159_1 );

 Adder29Bit Adder108(clk,  { x159_1[28: 0] },  {y70[23],y70[23],y70[23],y70[23],y70[23], y70[23: 0]  }, x160); 

 Register29Bit Reg375 (clk,x160, x160_1 );

 Adder29Bit Adder109(clk,  { x160_1[28: 0] },  {y71[23],y71[23],y71[23],y71[23],y71[23], y71[23: 0]  }, x161); 

 Register29Bit Reg376 (clk,x161, x161_1 );

 Adder29Bit Adder110(clk,  { x161_1[28: 0] },  {y72[22],y72[22],y72[22],y72[22],y72[22],y72[22], y72[22: 0]  }, x162); 

 Register29Bit Reg377 (clk,x162, x162_1 );

 Adder29Bit Adder111(clk,  { x162_1[28: 0] },  {y73[24],y73[24],y73[24],y73[24], y73[24: 0]  }, x163); 

 Register29Bit Reg378 (clk,x163, x163_1 );

 Adder29Bit Adder112(clk,  { x163_1[28: 0] },  {y74[23],y74[23],y74[23],y74[23],y74[23], y74[23: 0]  }, x164); 

 Register29Bit Reg379 (clk,x164, x164_1 );

 Adder29Bit Adder113(clk,  { x164_1[28: 0] },  {y75[21],y75[21],y75[21],y75[21],y75[21],y75[21],y75[21], y75[21: 0]  }, x165); 

 Register29Bit Reg380 (clk,x165, x165_1 );

 Adder29Bit Adder114(clk,  { x165_1[28: 0] },  {y76[23],y76[23],y76[23],y76[23],y76[23], y76[23: 0]  }, x166); 

 Register29Bit Reg381 (clk,x166, x166_1 );

 Adder29Bit Adder115(clk,  { x166_1[28: 0] },  {y77[20],y77[20],y77[20],y77[20],y77[20],y77[20],y77[20],y77[20], y77[20: 0]  }, x167); 

 Register29Bit Reg382 (clk,x167, x167_1 );

 Adder29Bit Adder116(clk,  { x167_1[28: 0] },  {y78[23],y78[23],y78[23],y78[23],y78[23], y78[23: 0]  }, x168); 

 Register29Bit Reg383 (clk,x168, x168_1 );

 Adder29Bit Adder117(clk,  { x168_1[28: 0] },  {y79[22],y79[22],y79[22],y79[22],y79[22],y79[22], y79[22: 0]  }, x169); 

 Register29Bit Reg384 (clk,x169, x169_1 );

 Adder29Bit Adder118(clk,  { x169_1[28: 0] },  {y80[22],y80[22],y80[22],y80[22],y80[22],y80[22], y80[22: 0]  }, x170); 

 Register29Bit Reg385 (clk,x170, x170_1 );

 Adder29Bit Adder119(clk,  { x170_1[28: 0] },  {y81[22],y81[22],y81[22],y81[22],y81[22],y81[22], y81[22: 0]  }, x171); 

 Register29Bit Reg386 (clk,x171, x171_1 );

 Adder29Bit Adder120(clk,  { x171_1[28: 0] },  {y82[22],y82[22],y82[22],y82[22],y82[22],y82[22], y82[22: 0]  }, x172); 

 Register29Bit Reg387 (clk,x172, x172_1 );

 Adder29Bit Adder121(clk,  { x172_1[28: 0] },  {y83[22],y83[22],y83[22],y83[22],y83[22],y83[22], y83[22: 0]  }, x173); 

 Register29Bit Reg388 (clk,x173, x173_1 );

 Adder29Bit Adder122(clk,  { x173_1[28: 0] },  {y84[19],y84[19],y84[19],y84[19],y84[19],y84[19],y84[19],y84[19],y84[19], y84[19: 0]  }, x174); 

 Register29Bit Reg389 (clk,x174, x174_1 );

 Adder29Bit Adder123(clk,  { x174_1[28: 0] },  {y85[21],y85[21],y85[21],y85[21],y85[21],y85[21],y85[21], y85[21: 0]  }, x175); 

 Register29Bit Reg390 (clk,x175, x175_1 );

 Adder29Bit Adder124(clk,  { x175_1[28: 0] },  {y86[20],y86[20],y86[20],y86[20],y86[20],y86[20],y86[20],y86[20], y86[20: 0]  }, x176); 

 Register29Bit Reg391 (clk,x176, x176_1 );

 Adder29Bit Adder125(clk,  { x176_1[28: 0] },  {y87[21],y87[21],y87[21],y87[21],y87[21],y87[21],y87[21], y87[21: 0]  }, x177); 

 Register29Bit Reg392 (clk,x177, x177_1 );

 Adder29Bit Adder126(clk,  { x177_1[28: 0] },  {y88[21],y88[21],y88[21],y88[21],y88[21],y88[21],y88[21], y88[21: 0]  }, x178); 

 Register29Bit Reg393 (clk,x178, x178_1 );

 Adder29Bit Adder127(clk,  { x178_1[28: 0] },  {y89[22],y89[22],y89[22],y89[22],y89[22],y89[22], y89[22: 0]  }, x179); 

 Register29Bit Reg394 (clk,x179, x179_1 );

 Adder29Bit Adder128(clk,  { x179_1[28: 0] },  {y90[21],y90[21],y90[21],y90[21],y90[21],y90[21],y90[21], y90[21: 0]  }, x180); 

 Register29Bit Reg395 (clk,x180, x180_1 );

 Adder29Bit Adder129(clk,  { x180_1[28: 0] },  {y91[20],y91[20],y91[20],y91[20],y91[20],y91[20],y91[20],y91[20], y91[20: 0]  }, x181); 

 Register29Bit Reg396 (clk,x181, x181_1 );

 Adder29Bit Adder130(clk,  { x181_1[28: 0] },  {y92[22],y92[22],y92[22],y92[22],y92[22],y92[22], y92[22: 0]  }, x182); 

 Register29Bit Reg397 (clk,x182, x182_1 );

 Adder29Bit Adder131(clk,  { x182_1[28: 0] },  {y93[16],y93[16],y93[16],y93[16],y93[16],y93[16],y93[16],y93[16],y93[16],y93[16],y93[16],y93[16], y93[16: 0]  }, x183); 

 Register29Bit Reg398 (clk,x183, x183_1 );

 Adder29Bit Adder132(clk,  { x183_1[28: 0] },  {y94[21],y94[21],y94[21],y94[21],y94[21],y94[21],y94[21], y94[21: 0]  }, x184); 

 Register29Bit Reg399 (clk,x184, x184_1 );

 Adder29Bit Adder133(clk,  { x184_1[28: 0] },  {y95[19],y95[19],y95[19],y95[19],y95[19],y95[19],y95[19],y95[19],y95[19], y95[19: 0]  }, x185); 

 Register29Bit Reg400 (clk,x185, x185_1 );

 Adder29Bit Adder134(clk,  { x185_1[28: 0] },  {y96[23],y96[23],y96[23],y96[23],y96[23], y96[23: 0]  }, x186); 

 Register29Bit Reg401 (clk,x186, x186_1 );

 Adder29Bit Adder135(clk,  { x186_1[28: 0] },  {y97[20],y97[20],y97[20],y97[20],y97[20],y97[20],y97[20],y97[20], y97[20: 0]  }, x187); 

 Register29Bit Reg402 (clk,x187, x187_1 );

 Adder29Bit Adder136(clk,  { x187_1[28: 0] },  {y98[20],y98[20],y98[20],y98[20],y98[20],y98[20],y98[20],y98[20], y98[20: 0]  }, x188); 

 Register29Bit Reg403 (clk,x188, x188_1 );

 Adder29Bit Adder137(clk,  { x188_1[28: 0] },  {y99[21],y99[21],y99[21],y99[21],y99[21],y99[21],y99[21], y99[21: 0]  }, x189); 

 Register29Bit Reg404 (clk,x189, x189_1 );

 Adder29Bit Adder138(clk,  { x189_1[28: 0] },  {y100[19],y100[19],y100[19],y100[19],y100[19],y100[19],y100[19],y100[19],y100[19], y100[19: 0]  }, x190); 

 Register29Bit Reg405 (clk,x190, x190_1 );

 Adder29Bit Adder139(clk,  { x190_1[28: 0] },  {y101[23],y101[23],y101[23],y101[23],y101[23], y101[23: 0]  }, x191); 

 Register29Bit Reg406 (clk,x191, x191_1 );

 Adder29Bit Adder140(clk,  { x191_1[28: 0] },  {y102[17],y102[17],y102[17],y102[17],y102[17],y102[17],y102[17],y102[17],y102[17],y102[17],y102[17], y102[17: 0]  }, x192); 

 Register29Bit Reg407 (clk,x192, x192_1 );

 Adder29Bit Adder141(clk,  { x192_1[28: 0] },  {y103[23],y103[23],y103[23],y103[23],y103[23], y103[23: 0]  }, x193); 

 Register29Bit Reg408 (clk,x193, x193_1 );

 Adder29Bit Adder142(clk,  { x193_1[28: 0] },  {y104[20],y104[20],y104[20],y104[20],y104[20],y104[20],y104[20],y104[20], y104[20: 0]  }, x194); 

 Register29Bit Reg409 (clk,x194, x194_1 );

 Adder29Bit Adder143(clk,  { x194_1[28: 0] },  {y105[21],y105[21],y105[21],y105[21],y105[21],y105[21],y105[21], y105[21: 0]  }, x195); 

 Register29Bit Reg410 (clk,x195, x195_1 );

 Adder29Bit Adder144(clk,  { x195_1[28: 0] },  {y106[20],y106[20],y106[20],y106[20],y106[20],y106[20],y106[20],y106[20], y106[20: 0]  }, x196); 

 Register29Bit Reg411 (clk,x196, x196_1 );

 Adder29Bit Adder145(clk,  { x196_1[28: 0] },  {y107[21],y107[21],y107[21],y107[21],y107[21],y107[21],y107[21], y107[21: 0]  }, x197); 

 Register29Bit Reg412 (clk,x197, x197_1 );

 Adder29Bit Adder146(clk,  { x197_1[28: 0] },  {y108[22],y108[22],y108[22],y108[22],y108[22],y108[22], y108[22: 0]  }, x198); 

 Register29Bit Reg413 (clk,x198, x198_1 );

 Adder29Bit Adder147(clk,  { x198_1[28: 0] },  {y109[20],y109[20],y109[20],y109[20],y109[20],y109[20],y109[20],y109[20], y109[20: 0]  }, x199); 

 Register29Bit Reg414 (clk,x199, x199_1 );

 Adder29Bit Adder148(clk,  { x199_1[28: 0] },  {y110[22],y110[22],y110[22],y110[22],y110[22],y110[22], y110[22: 0]  }, x200); 

 Register29Bit Reg415 (clk,x200, x200_1 );

 Adder29Bit Adder149(clk,  { x200_1[28: 0] },  {y111[17],y111[17],y111[17],y111[17],y111[17],y111[17],y111[17],y111[17],y111[17],y111[17],y111[17], y111[17: 0]  }, x201); 

 Register29Bit Reg416 (clk,x201, x201_1 );

 Adder29Bit Adder150(clk,  { x201_1[28: 0] },  {y112[21],y112[21],y112[21],y112[21],y112[21],y112[21],y112[21], y112[21: 0]  }, x202); 

 Register29Bit Reg417 (clk,x202, x202_1 );

 Adder29Bit Adder151(clk,  { x202_1[28: 0] },  {y113[19],y113[19],y113[19],y113[19],y113[19],y113[19],y113[19],y113[19],y113[19], y113[19: 0]  }, x203); 

 Register29Bit Reg418 (clk,x203, x203_1 );

 Adder29Bit Adder152(clk,  { x203_1[28: 0] },  {y114[23],y114[23],y114[23],y114[23],y114[23], y114[23: 0]  }, x204); 

 Register29Bit Reg419 (clk,x204, x204_1 );

 Adder29Bit Adder153(clk,  { x204_1[28: 0] },  {y115[20],y115[20],y115[20],y115[20],y115[20],y115[20],y115[20],y115[20], y115[20: 0]  }, x205); 

 Register29Bit Reg420 (clk,x205, x205_1 );

 Adder29Bit Adder154(clk,  { x205_1[28: 0] },  {y116[25],y116[25],y116[25], y116[25: 0]  }, x206); 

 Register29Bit Reg421 (clk,x206, x206_1 );

 Adder29Bit Adder155(clk,  { x206_1[28: 0] },  {y117[25],y117[25],y117[25], y117[25: 0]  }, x207); 

 Register29Bit Reg422 (clk,x207, x207_1 );

 Adder29Bit Adder156(clk,  { x207_1[28: 0] },  {y118[21],y118[21],y118[21],y118[21],y118[21],y118[21],y118[21], y118[21: 0]  }, Out_Y_wire); 

 endmodule 



module Adder16Bit (clk, In1, In2, AddOut);
 input clk;
 input [15:0] In1, In2; 

 output [16:0] AddOut;

 reg [16 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder22Bit (clk, In1, In2, AddOut);
 input clk;
 input [21:0] In1, In2; 

 output [22:0] AddOut;

 reg [22 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder19Bit (clk, In1, In2, AddOut);
 input clk;
 input [18:0] In1, In2; 

 output [19:0] AddOut;

 reg [19 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder21Bit (clk, In1, In2, AddOut);
 input clk;
 input [20:0] In1, In2; 

 output [21:0] AddOut;

 reg [21 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder23Bit (clk, In1, In2, AddOut);
 input clk;
 input [22:0] In1, In2; 

 output [23:0] AddOut;

 reg [23 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder26Bit (clk, In1, In2, AddOut);
 input clk;
 input [25:0] In1, In2; 

 output [26:0] AddOut;

 reg [26 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder17Bit (clk, In1, In2, AddOut);
 input clk;
 input [16:0] In1, In2; 

 output [17:0] AddOut;

 reg [17 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder24Bit (clk, In1, In2, AddOut);
 input clk;
 input [23:0] In1, In2; 

 output [24:0] AddOut;

 reg [24 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder20Bit (clk, In1, In2, AddOut);
 input clk;
 input [19:0] In1, In2; 

 output [20:0] AddOut;

 reg [20 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder25Bit (clk, In1, In2, AddOut);
 input clk;
 input [24:0] In1, In2; 

 output [25:0] AddOut;

 reg [25 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder14Bit (clk, In1, In2, AddOut);
 input clk;
 input [13:0] In1, In2; 

 output [14:0] AddOut;

 reg [14 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder15Bit (clk, In1, In2, AddOut);
 input clk;
 input [14:0] In1, In2; 

 output [15:0] AddOut;

 reg [15 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder27Bit (clk, In1, In2, AddOut);
 input clk;
 input [26:0] In1, In2; 

 output [27:0] AddOut;

 reg [27 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder28Bit (clk, In1, In2, AddOut);
 input clk;
 input [27:0] In1, In2; 

 output [28:0] AddOut;

 reg [28 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder29Bit (clk, In1, In2, AddOut);
 input clk;
 input [28:0] In1, In2; 

 output [28:0] AddOut;

 reg [28 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule



module Subtractor14Bit (clk, In1, In2, SubOut);
 input clk;
 input [13:0] In1, In2;
 output [14 :0] SubOut;

 reg [14 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule

module Subtractor21Bit (clk, In1, In2, SubOut);
 input clk;
 input [20:0] In1, In2;
 output [21 :0] SubOut;

 reg [21 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule

module Subtractor22Bit (clk, In1, In2, SubOut);
 input clk;
 input [21:0] In1, In2;
 output [22 :0] SubOut;

 reg [22 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule

module Subtractor24Bit (clk, In1, In2, SubOut);
 input clk;
 input [23:0] In1, In2;
 output [24 :0] SubOut;

 reg [24 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule

module Subtractor28Bit (clk, In1, In2, SubOut);
 input clk;
 input [27:0] In1, In2;
 output [28 :0] SubOut;

 reg [28 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule

module Subtractor19Bit (clk, In1, In2, SubOut);
 input clk;
 input [18:0] In1, In2;
 output [19 :0] SubOut;

 reg [19 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule

module Subtractor18Bit (clk, In1, In2, SubOut);
 input clk;
 input [17:0] In1, In2;
 output [18 :0] SubOut;

 reg [18 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule

module Subtractor20Bit (clk, In1, In2, SubOut);
 input clk;
 input [19:0] In1, In2;
 output [20 :0] SubOut;

 reg [20 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule

module Subtractor16Bit (clk, In1, In2, SubOut);
 input clk;
 input [15:0] In1, In2;
 output [16 :0] SubOut;

 reg [16 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule

module Subtractor25Bit (clk, In1, In2, SubOut);
 input clk;
 input [24:0] In1, In2;
 output [25 :0] SubOut;

 reg [25 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule

module Subtractor26Bit (clk, In1, In2, SubOut);
 input clk;
 input [25:0] In1, In2;
 output [26 :0] SubOut;

 reg [26 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule

module Subtractor23Bit (clk, In1, In2, SubOut);
 input clk;
 input [22:0] In1, In2;
 output [23 :0] SubOut;

 reg [23 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule

module Subtractor17Bit (clk, In1, In2, SubOut);
 input clk;
 input [16:0] In1, In2;
 output [17 :0] SubOut;

 reg [17 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule

module Subtractor27Bit (clk, In1, In2, SubOut);
 input clk;
 input [26:0] In1, In2;
 output [27 :0] SubOut;

 reg [27 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule

module Subtractor15Bit (clk, In1, In2, SubOut);
 input clk;
 input [14:0] In1, In2;
 output [15 :0] SubOut;

 reg [15 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule



module Register22Bit (clk, In1, RegOut);
 input clk;
 input [21:0] In1;
 output [21 :0] RegOut;

 reg [21 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register23Bit (clk, In1, RegOut);
 input clk;
 input [22:0] In1;
 output [22 :0] RegOut;

 reg [22 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register25Bit (clk, In1, RegOut);
 input clk;
 input [24:0] In1;
 output [24 :0] RegOut;

 reg [24 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register29Bit (clk, In1, RegOut);
 input clk;
 input [28:0] In1;
 output [28 :0] RegOut;

 reg [28 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register21Bit (clk, In1, RegOut);
 input clk;
 input [20:0] In1;
 output [20 :0] RegOut;

 reg [20 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register20Bit (clk, In1, RegOut);
 input clk;
 input [19:0] In1;
 output [19 :0] RegOut;

 reg [19 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register24Bit (clk, In1, RegOut);
 input clk;
 input [23:0] In1;
 output [23 :0] RegOut;

 reg [23 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register26Bit (clk, In1, RegOut);
 input clk;
 input [25:0] In1;
 output [25 :0] RegOut;

 reg [25 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register27Bit (clk, In1, RegOut);
 input clk;
 input [26:0] In1;
 output [26 :0] RegOut;

 reg [26 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register19Bit (clk, In1, RegOut);
 input clk;
 input [18:0] In1;
 output [18 :0] RegOut;

 reg [18 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register15Bit (clk, In1, RegOut);
 input clk;
 input [14:0] In1;
 output [14 :0] RegOut;

 reg [14 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register17Bit (clk, In1, RegOut);
 input clk;
 input [16:0] In1;
 output [16 :0] RegOut;

 reg [16 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register18Bit (clk, In1, RegOut);
 input clk;
 input [17:0] In1;
 output [17 :0] RegOut;

 reg [17 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register16Bit (clk, In1, RegOut);
 input clk;
 input [15:0] In1;
 output [15 :0] RegOut;

 reg [15 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register12Bit (clk, In1, RegOut);
 input clk;
 input [11:0] In1;
 output [11 :0] RegOut;

 reg [11 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register28Bit (clk, In1, RegOut);
 input clk;
 input [27:0] In1;
 output [27 :0] RegOut;

 reg [27 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule



module Negator20Bit (clk, In1, NegOut);
 input clk;
 input [19:0] In1;
 output [19 :0] NegOut;

 reg [19 :0] NegOut; 

always @(posedge clk)
begin
NegOut <= -(In1);
end
endmodule

module Negator24Bit (clk, In1, NegOut);
 input clk;
 input [23:0] In1;
 output [23 :0] NegOut;

 reg [23 :0] NegOut; 

always @(posedge clk)
begin
NegOut <= -(In1);
end
endmodule

module Negator27Bit (clk, In1, NegOut);
 input clk;
 input [26:0] In1;
 output [26 :0] NegOut;

 reg [26 :0] NegOut; 

always @(posedge clk)
begin
NegOut <= -(In1);
end
endmodule

module Negator23Bit (clk, In1, NegOut);
 input clk;
 input [22:0] In1;
 output [22 :0] NegOut;

 reg [22 :0] NegOut; 

always @(posedge clk)
begin
NegOut <= -(In1);
end
endmodule

module Negator26Bit (clk, In1, NegOut);
 input clk;
 input [25:0] In1;
 output [25 :0] NegOut;

 reg [25 :0] NegOut; 

always @(posedge clk)
begin
NegOut <= -(In1);
end
endmodule

module Negator21Bit (clk, In1, NegOut);
 input clk;
 input [20:0] In1;
 output [20 :0] NegOut;

 reg [20 :0] NegOut; 

always @(posedge clk)
begin
NegOut <= -(In1);
end
endmodule

module Negator22Bit (clk, In1, NegOut);
 input clk;
 input [21:0] In1;
 output [21 :0] NegOut;

 reg [21 :0] NegOut; 

always @(posedge clk)
begin
NegOut <= -(In1);
end
endmodule

module Negator15Bit (clk, In1, NegOut);
 input clk;
 input [14:0] In1;
 output [14 :0] NegOut;

 reg [14 :0] NegOut; 

always @(posedge clk)
begin
NegOut <= -(In1);
end
endmodule

module Negator18Bit (clk, In1, NegOut);
 input clk;
 input [17:0] In1;
 output [17 :0] NegOut;

 reg [17 :0] NegOut; 

always @(posedge clk)
begin
NegOut <= -(In1);
end
endmodule
