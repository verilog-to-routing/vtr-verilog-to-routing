/*
 * Ultra wide range test
*/

`define WIDTH 256
`define operator and
`include "replicate_any_width_binary_test.v"