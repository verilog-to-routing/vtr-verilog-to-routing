module simple_op ( input in,
                                output out );

    assign out = in >> 1;

endmodule
