`define BINARY_OP(out,a,b) bufif0(out, a, b);
`include "../.generic/wire_test.v"