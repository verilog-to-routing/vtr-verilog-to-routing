/*
 * Ultra wide range test
*/

`define WIDTH 256
`define operator notif0
`include "../.generic/range_any_width_binary_test.v"