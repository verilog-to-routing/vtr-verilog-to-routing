`define UNARY_OP(out,a) buf(out, a);
`include "../.generic/wire_test.v"