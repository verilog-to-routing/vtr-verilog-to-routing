module simple_op ( input [2:0] in,
                                output [2:0] out );

    assign out = in >> 2;

endmodule
