/*
 * Integer wide range test
*/

`define WIDTH 32
`define operator xor
`include "replicate_any_width_binary_test.v"