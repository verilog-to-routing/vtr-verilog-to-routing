module simple_op(a,c);
input a;

output c;

wire a,c;

assign c = a;

endmodule