
    // RC4 PRGA module implementation
    // Copyright 2012 - Alfredo Ortega
	// aortega@alu.itba.edu.ar
	// aortega@groundworkstech.com

 // This library is free software: you can redistribute it and/or
 // modify it under the terms of the GNU Lesser General Public
 // License as published by the Free Software Foundation, either
 // version 3 of the License, or (at your option) any later version.

 // This library is distributed in the hope that it will be useful,
 // but WITHOUT ANY WARRANTY; without even the implied warranty of
 // MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
 // Lesser General Public License for more details.

 // You should have received a copy of the GNU Lesser General Public
 // License along with this library.  If not, see <http://www.gnu.org/licenses/>.



	// RC4 PRGA constants
	// Copyright 2012 - Alfredo Ortega
	// aortega@alu.itba.edu.ar

 // This library is free software: you can redistribute it and/or
 // modify it under the terms of the GNU Lesser General Public
 // License as published by the Free Software Foundation, either
 // version 3 of the License, or (at your option) any later version.

 // This library is distributed in the hope that it will be useful,
 // but WITHOUT ANY WARRANTY; without even the implied warranty of
 // MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
 // Lesser General Public License for more details.

 // You should have received a copy of the GNU Lesser General Public
 // License along with this library.  If not, see <http://www.gnu.org/licenses/>.

//%%GENDEFINE%% (choose_to,   nonblocking, 0, 256 )
//%%GENDEFINE%% (choose_from, blocking,    0, 256 )
//%%GENDEFINE%% (choose_from, nonblocking, 0, 256 )
//%%GENDEFINE%% (choose_to,   nonblocking, 0, 255 )
//%%GENDEFINE%% (choose_from, blocking,    0, 255 )
//%%GENDEFINE%% (choose_from, nonblocking, 0, 255 )

//%%GENDEFINE%% (choose_to,   nonblocking, 0, 6   )
//%%GENDEFINE%% (choose_from, blocking,    0, 6   )
//%%GENDEFINE%% (choose_from, blocking,    0, 6   )

//%%GENDEFINE%% (always_list, 0, 256)
//%%GENDEFINE%% (always_list, 0, 255)
//%%GENDEFINE%% (always_list, 0, 6)

//%%GENDEFINE%% (mod_op, blocking, 7, 0, 255)



module rc4(clk,
rst,
output_ready,
password_input,
K);


input clk; // Clock
input rst; // Reset
input [7:0] password_input; // Password input
output output_ready; // Output valid
output [7:0] K; // Output port


wire clk, rst; // clock, reset
reg output_ready;
wire [7:0] password_input;


 // RC4 PRGA

// Key
reg [7:0] key_0;
reg [7:0] key_1;
reg [7:0] key_2;
reg [7:0] key_3;
reg [7:0] key_4;
reg [7:0] key_5;
reg [7:0] key_6;

// S array
reg [7:0] S_0;
reg [7:0] S_1;
reg [7:0] S_2;
reg [7:0] S_3;
reg [7:0] S_4;
reg [7:0] S_5;
reg [7:0] S_6;
reg [7:0] S_7;
reg [7:0] S_8;
reg [7:0] S_9;
reg [7:0] S_10;
reg [7:0] S_11;
reg [7:0] S_12;
reg [7:0] S_13;
reg [7:0] S_14;
reg [7:0] S_15;
reg [7:0] S_16;
reg [7:0] S_17;
reg [7:0] S_18;
reg [7:0] S_19;
reg [7:0] S_20;
reg [7:0] S_21;
reg [7:0] S_22;
reg [7:0] S_23;
reg [7:0] S_24;
reg [7:0] S_25;
reg [7:0] S_26;
reg [7:0] S_27;
reg [7:0] S_28;
reg [7:0] S_29;
reg [7:0] S_30;
reg [7:0] S_31;
reg [7:0] S_32;
reg [7:0] S_33;
reg [7:0] S_34;
reg [7:0] S_35;
reg [7:0] S_36;
reg [7:0] S_37;
reg [7:0] S_38;
reg [7:0] S_39;
reg [7:0] S_40;
reg [7:0] S_41;
reg [7:0] S_42;
reg [7:0] S_43;
reg [7:0] S_44;
reg [7:0] S_45;
reg [7:0] S_46;
reg [7:0] S_47;
reg [7:0] S_48;
reg [7:0] S_49;
reg [7:0] S_50;
reg [7:0] S_51;
reg [7:0] S_52;
reg [7:0] S_53;
reg [7:0] S_54;
reg [7:0] S_55;
reg [7:0] S_56;
reg [7:0] S_57;
reg [7:0] S_58;
reg [7:0] S_59;
reg [7:0] S_60;
reg [7:0] S_61;
reg [7:0] S_62;
reg [7:0] S_63;
reg [7:0] S_64;
reg [7:0] S_65;
reg [7:0] S_66;
reg [7:0] S_67;
reg [7:0] S_68;
reg [7:0] S_69;
reg [7:0] S_70;
reg [7:0] S_71;
reg [7:0] S_72;
reg [7:0] S_73;
reg [7:0] S_74;
reg [7:0] S_75;
reg [7:0] S_76;
reg [7:0] S_77;
reg [7:0] S_78;
reg [7:0] S_79;
reg [7:0] S_80;
reg [7:0] S_81;
reg [7:0] S_82;
reg [7:0] S_83;
reg [7:0] S_84;
reg [7:0] S_85;
reg [7:0] S_86;
reg [7:0] S_87;
reg [7:0] S_88;
reg [7:0] S_89;
reg [7:0] S_90;
reg [7:0] S_91;
reg [7:0] S_92;
reg [7:0] S_93;
reg [7:0] S_94;
reg [7:0] S_95;
reg [7:0] S_96;
reg [7:0] S_97;
reg [7:0] S_98;
reg [7:0] S_99;
reg [7:0] S_100;
reg [7:0] S_101;
reg [7:0] S_102;
reg [7:0] S_103;
reg [7:0] S_104;
reg [7:0] S_105;
reg [7:0] S_106;
reg [7:0] S_107;
reg [7:0] S_108;
reg [7:0] S_109;
reg [7:0] S_110;
reg [7:0] S_111;
reg [7:0] S_112;
reg [7:0] S_113;
reg [7:0] S_114;
reg [7:0] S_115;
reg [7:0] S_116;
reg [7:0] S_117;
reg [7:0] S_118;
reg [7:0] S_119;
reg [7:0] S_120;
reg [7:0] S_121;
reg [7:0] S_122;
reg [7:0] S_123;
reg [7:0] S_124;
reg [7:0] S_125;
reg [7:0] S_126;
reg [7:0] S_127;
reg [7:0] S_128;
reg [7:0] S_129;
reg [7:0] S_130;
reg [7:0] S_131;
reg [7:0] S_132;
reg [7:0] S_133;
reg [7:0] S_134;
reg [7:0] S_135;
reg [7:0] S_136;
reg [7:0] S_137;
reg [7:0] S_138;
reg [7:0] S_139;
reg [7:0] S_140;
reg [7:0] S_141;
reg [7:0] S_142;
reg [7:0] S_143;
reg [7:0] S_144;
reg [7:0] S_145;
reg [7:0] S_146;
reg [7:0] S_147;
reg [7:0] S_148;
reg [7:0] S_149;
reg [7:0] S_150;
reg [7:0] S_151;
reg [7:0] S_152;
reg [7:0] S_153;
reg [7:0] S_154;
reg [7:0] S_155;
reg [7:0] S_156;
reg [7:0] S_157;
reg [7:0] S_158;
reg [7:0] S_159;
reg [7:0] S_160;
reg [7:0] S_161;
reg [7:0] S_162;
reg [7:0] S_163;
reg [7:0] S_164;
reg [7:0] S_165;
reg [7:0] S_166;
reg [7:0] S_167;
reg [7:0] S_168;
reg [7:0] S_169;
reg [7:0] S_170;
reg [7:0] S_171;
reg [7:0] S_172;
reg [7:0] S_173;
reg [7:0] S_174;
reg [7:0] S_175;
reg [7:0] S_176;
reg [7:0] S_177;
reg [7:0] S_178;
reg [7:0] S_179;
reg [7:0] S_180;
reg [7:0] S_181;
reg [7:0] S_182;
reg [7:0] S_183;
reg [7:0] S_184;
reg [7:0] S_185;
reg [7:0] S_186;
reg [7:0] S_187;
reg [7:0] S_188;
reg [7:0] S_189;
reg [7:0] S_190;
reg [7:0] S_191;
reg [7:0] S_192;
reg [7:0] S_193;
reg [7:0] S_194;
reg [7:0] S_195;
reg [7:0] S_196;
reg [7:0] S_197;
reg [7:0] S_198;
reg [7:0] S_199;
reg [7:0] S_200;
reg [7:0] S_201;
reg [7:0] S_202;
reg [7:0] S_203;
reg [7:0] S_204;
reg [7:0] S_205;
reg [7:0] S_206;
reg [7:0] S_207;
reg [7:0] S_208;
reg [7:0] S_209;
reg [7:0] S_210;
reg [7:0] S_211;
reg [7:0] S_212;
reg [7:0] S_213;
reg [7:0] S_214;
reg [7:0] S_215;
reg [7:0] S_216;
reg [7:0] S_217;
reg [7:0] S_218;
reg [7:0] S_219;
reg [7:0] S_220;
reg [7:0] S_221;
reg [7:0] S_222;
reg [7:0] S_223;
reg [7:0] S_224;
reg [7:0] S_225;
reg [7:0] S_226;
reg [7:0] S_227;
reg [7:0] S_228;
reg [7:0] S_229;
reg [7:0] S_230;
reg [7:0] S_231;
reg [7:0] S_232;
reg [7:0] S_233;
reg [7:0] S_234;
reg [7:0] S_235;
reg [7:0] S_236;
reg [7:0] S_237;
reg [7:0] S_238;
reg [7:0] S_239;
reg [7:0] S_240;
reg [7:0] S_241;
reg [7:0] S_242;
reg [7:0] S_243;
reg [7:0] S_244;
reg [7:0] S_245;
reg [7:0] S_246;
reg [7:0] S_247;
reg [7:0] S_248;
reg [7:0] S_249;
reg [7:0] S_250;
reg [7:0] S_251;
reg [7:0] S_252;
reg [7:0] S_253;
reg [7:0] S_254;
reg [7:0] S_255;
reg [7:0] S_256;

reg [10:0] discardCount;

// Key-scheduling state

// Variable names from http://en.wikipedia.org/wiki/RC4
reg [3:0] KSState;
reg [7:0] i; // Counter
reg [7:0] j;
reg [7:0] K;


reg [7:0] S_of_i;
reg [7:0] S_of_i_plus_1;
reg [7:0] S_of_j;
wire [7:0] S_of_i_plus_S_of_j;

reg [7:0] prev_i;
reg [7:0] prev_S_of_j;

reg [7:0]  key_of_i_mod_KEYSIZE;
reg [7:0] i_mod_KEYSIZE;

always @ (i or S_0 or S_1 or S_2 or S_3 or S_4 or S_5 or S_6 or S_7 or S_8 or S_9 or S_10 or S_11 or S_12 or S_13 or S_14 or S_15 or S_16 or S_17 or S_18 or S_19 or S_20 or S_21 or S_22 or S_23 or S_24 or S_25 or S_26 or S_27 or S_28 or S_29 or S_30 or S_31 or S_32 or S_33 or S_34 or S_35 or S_36 or S_37 or S_38 or S_39 or S_40 or S_41 or S_42 or S_43 or S_44 or S_45 or S_46 or S_47 or S_48 or S_49 or S_50 or S_51 or S_52 or S_53 or S_54 or S_55 or S_56 or S_57 or S_58 or S_59 or S_60 or S_61 or S_62 or S_63 or S_64 or S_65 or S_66 or S_67 or S_68 or S_69 or S_70 or S_71 or S_72 or S_73 or S_74 or S_75 or S_76 or S_77 or S_78 or S_79 or S_80 or S_81 or S_82 or S_83 or S_84 or S_85 or S_86 or S_87 or S_88 or S_89 or S_90 or S_91 or S_92 or S_93 or S_94 or S_95 or S_96 or S_97 or S_98 or S_99 or S_100 or S_101 or S_102 or S_103 or S_104 or S_105 or S_106 or S_107 or S_108 or S_109 or S_110 or S_111 or S_112 or S_113 or S_114 or S_115 or S_116 or S_117 or S_118 or S_119 or S_120 or S_121 or S_122 or S_123 or S_124 or S_125 or S_126 or S_127 or S_128 or S_129 or S_130 or S_131 or S_132 or S_133 or S_134 or S_135 or S_136 or S_137 or S_138 or S_139 or S_140 or S_141 or S_142 or S_143 or S_144 or S_145 or S_146 or S_147 or S_148 or S_149 or S_150 or S_151 or S_152 or S_153 or S_154 or S_155 or S_156 or S_157 or S_158 or S_159 or S_160 or S_161 or S_162 or S_163 or S_164 or S_165 or S_166 or S_167 or S_168 or S_169 or S_170 or S_171 or S_172 or S_173 or S_174 or S_175 or S_176 or S_177 or S_178 or S_179 or S_180 or S_181 or S_182 or S_183 or S_184 or S_185 or S_186 or S_187 or S_188 or S_189 or S_190 or S_191 or S_192 or S_193 or S_194 or S_195 or S_196 or S_197 or S_198 or S_199 or S_200 or S_201 or S_202 or S_203 or S_204 or S_205 or S_206 or S_207 or S_208 or S_209 or S_210 or S_211 or S_212 or S_213 or S_214 or S_215 or S_216 or S_217 or S_218 or S_219 or S_220 or S_221 or S_222 or S_223 or S_224 or S_225 or S_226 or S_227 or S_228 or S_229 or S_230 or S_231 or S_232 or S_233 or S_234 or S_235 or S_236 or S_237 or S_238 or S_239 or S_240 or S_241 or S_242 or S_243 or S_244 or S_245 or S_246 or S_247 or S_248 or S_249 or S_250 or S_251 or S_252 or S_253 or S_254 or S_255) begin
	case (i) 
		'd0:S_of_i = S_0; 
		'd1:S_of_i = S_1; 
		'd2:S_of_i = S_2; 
		'd3:S_of_i = S_3; 
		'd4:S_of_i = S_4; 
		'd5:S_of_i = S_5; 
		'd6:S_of_i = S_6; 
		'd7:S_of_i = S_7; 
		'd8:S_of_i = S_8; 
		'd9:S_of_i = S_9; 
		'd10:S_of_i = S_10; 
		'd11:S_of_i = S_11; 
		'd12:S_of_i = S_12; 
		'd13:S_of_i = S_13; 
		'd14:S_of_i = S_14; 
		'd15:S_of_i = S_15; 
		'd16:S_of_i = S_16; 
		'd17:S_of_i = S_17; 
		'd18:S_of_i = S_18; 
		'd19:S_of_i = S_19; 
		'd20:S_of_i = S_20; 
		'd21:S_of_i = S_21; 
		'd22:S_of_i = S_22; 
		'd23:S_of_i = S_23; 
		'd24:S_of_i = S_24; 
		'd25:S_of_i = S_25; 
		'd26:S_of_i = S_26; 
		'd27:S_of_i = S_27; 
		'd28:S_of_i = S_28; 
		'd29:S_of_i = S_29; 
		'd30:S_of_i = S_30; 
		'd31:S_of_i = S_31; 
		'd32:S_of_i = S_32; 
		'd33:S_of_i = S_33; 
		'd34:S_of_i = S_34; 
		'd35:S_of_i = S_35; 
		'd36:S_of_i = S_36; 
		'd37:S_of_i = S_37; 
		'd38:S_of_i = S_38; 
		'd39:S_of_i = S_39; 
		'd40:S_of_i = S_40; 
		'd41:S_of_i = S_41; 
		'd42:S_of_i = S_42; 
		'd43:S_of_i = S_43; 
		'd44:S_of_i = S_44; 
		'd45:S_of_i = S_45; 
		'd46:S_of_i = S_46; 
		'd47:S_of_i = S_47; 
		'd48:S_of_i = S_48; 
		'd49:S_of_i = S_49; 
		'd50:S_of_i = S_50; 
		'd51:S_of_i = S_51; 
		'd52:S_of_i = S_52; 
		'd53:S_of_i = S_53; 
		'd54:S_of_i = S_54; 
		'd55:S_of_i = S_55; 
		'd56:S_of_i = S_56; 
		'd57:S_of_i = S_57; 
		'd58:S_of_i = S_58; 
		'd59:S_of_i = S_59; 
		'd60:S_of_i = S_60; 
		'd61:S_of_i = S_61; 
		'd62:S_of_i = S_62; 
		'd63:S_of_i = S_63; 
		'd64:S_of_i = S_64; 
		'd65:S_of_i = S_65; 
		'd66:S_of_i = S_66; 
		'd67:S_of_i = S_67; 
		'd68:S_of_i = S_68; 
		'd69:S_of_i = S_69; 
		'd70:S_of_i = S_70; 
		'd71:S_of_i = S_71; 
		'd72:S_of_i = S_72; 
		'd73:S_of_i = S_73; 
		'd74:S_of_i = S_74; 
		'd75:S_of_i = S_75; 
		'd76:S_of_i = S_76; 
		'd77:S_of_i = S_77; 
		'd78:S_of_i = S_78; 
		'd79:S_of_i = S_79; 
		'd80:S_of_i = S_80; 
		'd81:S_of_i = S_81; 
		'd82:S_of_i = S_82; 
		'd83:S_of_i = S_83; 
		'd84:S_of_i = S_84; 
		'd85:S_of_i = S_85; 
		'd86:S_of_i = S_86; 
		'd87:S_of_i = S_87; 
		'd88:S_of_i = S_88; 
		'd89:S_of_i = S_89; 
		'd90:S_of_i = S_90; 
		'd91:S_of_i = S_91; 
		'd92:S_of_i = S_92; 
		'd93:S_of_i = S_93; 
		'd94:S_of_i = S_94; 
		'd95:S_of_i = S_95; 
		'd96:S_of_i = S_96; 
		'd97:S_of_i = S_97; 
		'd98:S_of_i = S_98; 
		'd99:S_of_i = S_99; 
		'd100:S_of_i = S_100; 
		'd101:S_of_i = S_101; 
		'd102:S_of_i = S_102; 
		'd103:S_of_i = S_103; 
		'd104:S_of_i = S_104; 
		'd105:S_of_i = S_105; 
		'd106:S_of_i = S_106; 
		'd107:S_of_i = S_107; 
		'd108:S_of_i = S_108; 
		'd109:S_of_i = S_109; 
		'd110:S_of_i = S_110; 
		'd111:S_of_i = S_111; 
		'd112:S_of_i = S_112; 
		'd113:S_of_i = S_113; 
		'd114:S_of_i = S_114; 
		'd115:S_of_i = S_115; 
		'd116:S_of_i = S_116; 
		'd117:S_of_i = S_117; 
		'd118:S_of_i = S_118; 
		'd119:S_of_i = S_119; 
		'd120:S_of_i = S_120; 
		'd121:S_of_i = S_121; 
		'd122:S_of_i = S_122; 
		'd123:S_of_i = S_123; 
		'd124:S_of_i = S_124; 
		'd125:S_of_i = S_125; 
		'd126:S_of_i = S_126; 
		'd127:S_of_i = S_127; 
		'd128:S_of_i = S_128; 
		'd129:S_of_i = S_129; 
		'd130:S_of_i = S_130; 
		'd131:S_of_i = S_131; 
		'd132:S_of_i = S_132; 
		'd133:S_of_i = S_133; 
		'd134:S_of_i = S_134; 
		'd135:S_of_i = S_135; 
		'd136:S_of_i = S_136; 
		'd137:S_of_i = S_137; 
		'd138:S_of_i = S_138; 
		'd139:S_of_i = S_139; 
		'd140:S_of_i = S_140; 
		'd141:S_of_i = S_141; 
		'd142:S_of_i = S_142; 
		'd143:S_of_i = S_143; 
		'd144:S_of_i = S_144; 
		'd145:S_of_i = S_145; 
		'd146:S_of_i = S_146; 
		'd147:S_of_i = S_147; 
		'd148:S_of_i = S_148; 
		'd149:S_of_i = S_149; 
		'd150:S_of_i = S_150; 
		'd151:S_of_i = S_151; 
		'd152:S_of_i = S_152; 
		'd153:S_of_i = S_153; 
		'd154:S_of_i = S_154; 
		'd155:S_of_i = S_155; 
		'd156:S_of_i = S_156; 
		'd157:S_of_i = S_157; 
		'd158:S_of_i = S_158; 
		'd159:S_of_i = S_159; 
		'd160:S_of_i = S_160; 
		'd161:S_of_i = S_161; 
		'd162:S_of_i = S_162; 
		'd163:S_of_i = S_163; 
		'd164:S_of_i = S_164; 
		'd165:S_of_i = S_165; 
		'd166:S_of_i = S_166; 
		'd167:S_of_i = S_167; 
		'd168:S_of_i = S_168; 
		'd169:S_of_i = S_169; 
		'd170:S_of_i = S_170; 
		'd171:S_of_i = S_171; 
		'd172:S_of_i = S_172; 
		'd173:S_of_i = S_173; 
		'd174:S_of_i = S_174; 
		'd175:S_of_i = S_175; 
		'd176:S_of_i = S_176; 
		'd177:S_of_i = S_177; 
		'd178:S_of_i = S_178; 
		'd179:S_of_i = S_179; 
		'd180:S_of_i = S_180; 
		'd181:S_of_i = S_181; 
		'd182:S_of_i = S_182; 
		'd183:S_of_i = S_183; 
		'd184:S_of_i = S_184; 
		'd185:S_of_i = S_185; 
		'd186:S_of_i = S_186; 
		'd187:S_of_i = S_187; 
		'd188:S_of_i = S_188; 
		'd189:S_of_i = S_189; 
		'd190:S_of_i = S_190; 
		'd191:S_of_i = S_191; 
		'd192:S_of_i = S_192; 
		'd193:S_of_i = S_193; 
		'd194:S_of_i = S_194; 
		'd195:S_of_i = S_195; 
		'd196:S_of_i = S_196; 
		'd197:S_of_i = S_197; 
		'd198:S_of_i = S_198; 
		'd199:S_of_i = S_199; 
		'd200:S_of_i = S_200; 
		'd201:S_of_i = S_201; 
		'd202:S_of_i = S_202; 
		'd203:S_of_i = S_203; 
		'd204:S_of_i = S_204; 
		'd205:S_of_i = S_205; 
		'd206:S_of_i = S_206; 
		'd207:S_of_i = S_207; 
		'd208:S_of_i = S_208; 
		'd209:S_of_i = S_209; 
		'd210:S_of_i = S_210; 
		'd211:S_of_i = S_211; 
		'd212:S_of_i = S_212; 
		'd213:S_of_i = S_213; 
		'd214:S_of_i = S_214; 
		'd215:S_of_i = S_215; 
		'd216:S_of_i = S_216; 
		'd217:S_of_i = S_217; 
		'd218:S_of_i = S_218; 
		'd219:S_of_i = S_219; 
		'd220:S_of_i = S_220; 
		'd221:S_of_i = S_221; 
		'd222:S_of_i = S_222; 
		'd223:S_of_i = S_223; 
		'd224:S_of_i = S_224; 
		'd225:S_of_i = S_225; 
		'd226:S_of_i = S_226; 
		'd227:S_of_i = S_227; 
		'd228:S_of_i = S_228; 
		'd229:S_of_i = S_229; 
		'd230:S_of_i = S_230; 
		'd231:S_of_i = S_231; 
		'd232:S_of_i = S_232; 
		'd233:S_of_i = S_233; 
		'd234:S_of_i = S_234; 
		'd235:S_of_i = S_235; 
		'd236:S_of_i = S_236; 
		'd237:S_of_i = S_237; 
		'd238:S_of_i = S_238; 
		'd239:S_of_i = S_239; 
		'd240:S_of_i = S_240; 
		'd241:S_of_i = S_241; 
		'd242:S_of_i = S_242; 
		'd243:S_of_i = S_243; 
		'd244:S_of_i = S_244; 
		'd245:S_of_i = S_245; 
		'd246:S_of_i = S_246; 
		'd247:S_of_i = S_247; 
		'd248:S_of_i = S_248; 
		'd249:S_of_i = S_249; 
		'd250:S_of_i = S_250; 
		'd251:S_of_i = S_251; 
		'd252:S_of_i = S_252; 
		'd253:S_of_i = S_253; 
		'd254:S_of_i = S_254; 
		default:S_of_i = S_255; 
	endcase
end
always @ (i or S_0 or S_1 or S_2 or S_3 or S_4 or S_5 or S_6 or S_7 or S_8 or S_9 or S_10 or S_11 or S_12 or S_13 or S_14 or S_15 or S_16 or S_17 or S_18 or S_19 or S_20 or S_21 or S_22 or S_23 or S_24 or S_25 or S_26 or S_27 or S_28 or S_29 or S_30 or S_31 or S_32 or S_33 or S_34 or S_35 or S_36 or S_37 or S_38 or S_39 or S_40 or S_41 or S_42 or S_43 or S_44 or S_45 or S_46 or S_47 or S_48 or S_49 or S_50 or S_51 or S_52 or S_53 or S_54 or S_55 or S_56 or S_57 or S_58 or S_59 or S_60 or S_61 or S_62 or S_63 or S_64 or S_65 or S_66 or S_67 or S_68 or S_69 or S_70 or S_71 or S_72 or S_73 or S_74 or S_75 or S_76 or S_77 or S_78 or S_79 or S_80 or S_81 or S_82 or S_83 or S_84 or S_85 or S_86 or S_87 or S_88 or S_89 or S_90 or S_91 or S_92 or S_93 or S_94 or S_95 or S_96 or S_97 or S_98 or S_99 or S_100 or S_101 or S_102 or S_103 or S_104 or S_105 or S_106 or S_107 or S_108 or S_109 or S_110 or S_111 or S_112 or S_113 or S_114 or S_115 or S_116 or S_117 or S_118 or S_119 or S_120 or S_121 or S_122 or S_123 or S_124 or S_125 or S_126 or S_127 or S_128 or S_129 or S_130 or S_131 or S_132 or S_133 or S_134 or S_135 or S_136 or S_137 or S_138 or S_139 or S_140 or S_141 or S_142 or S_143 or S_144 or S_145 or S_146 or S_147 or S_148 or S_149 or S_150 or S_151 or S_152 or S_153 or S_154 or S_155 or S_156 or S_157 or S_158 or S_159 or S_160 or S_161 or S_162 or S_163 or S_164 or S_165 or S_166 or S_167 or S_168 or S_169 or S_170 or S_171 or S_172 or S_173 or S_174 or S_175 or S_176 or S_177 or S_178 or S_179 or S_180 or S_181 or S_182 or S_183 or S_184 or S_185 or S_186 or S_187 or S_188 or S_189 or S_190 or S_191 or S_192 or S_193 or S_194 or S_195 or S_196 or S_197 or S_198 or S_199 or S_200 or S_201 or S_202 or S_203 or S_204 or S_205 or S_206 or S_207 or S_208 or S_209 or S_210 or S_211 or S_212 or S_213 or S_214 or S_215 or S_216 or S_217 or S_218 or S_219 or S_220 or S_221 or S_222 or S_223 or S_224 or S_225 or S_226 or S_227 or S_228 or S_229 or S_230 or S_231 or S_232 or S_233 or S_234 or S_235 or S_236 or S_237 or S_238 or S_239 or S_240 or S_241 or S_242 or S_243 or S_244 or S_245 or S_246 or S_247 or S_248 or S_249 or S_250 or S_251 or S_252 or S_253 or S_254 or S_255 or S_256) begin
	case (i+1) 
		'd0:S_of_i_plus_1 = S_0; 
		'd1:S_of_i_plus_1 = S_1; 
		'd2:S_of_i_plus_1 = S_2; 
		'd3:S_of_i_plus_1 = S_3; 
		'd4:S_of_i_plus_1 = S_4; 
		'd5:S_of_i_plus_1 = S_5; 
		'd6:S_of_i_plus_1 = S_6; 
		'd7:S_of_i_plus_1 = S_7; 
		'd8:S_of_i_plus_1 = S_8; 
		'd9:S_of_i_plus_1 = S_9; 
		'd10:S_of_i_plus_1 = S_10; 
		'd11:S_of_i_plus_1 = S_11; 
		'd12:S_of_i_plus_1 = S_12; 
		'd13:S_of_i_plus_1 = S_13; 
		'd14:S_of_i_plus_1 = S_14; 
		'd15:S_of_i_plus_1 = S_15; 
		'd16:S_of_i_plus_1 = S_16; 
		'd17:S_of_i_plus_1 = S_17; 
		'd18:S_of_i_plus_1 = S_18; 
		'd19:S_of_i_plus_1 = S_19; 
		'd20:S_of_i_plus_1 = S_20; 
		'd21:S_of_i_plus_1 = S_21; 
		'd22:S_of_i_plus_1 = S_22; 
		'd23:S_of_i_plus_1 = S_23; 
		'd24:S_of_i_plus_1 = S_24; 
		'd25:S_of_i_plus_1 = S_25; 
		'd26:S_of_i_plus_1 = S_26; 
		'd27:S_of_i_plus_1 = S_27; 
		'd28:S_of_i_plus_1 = S_28; 
		'd29:S_of_i_plus_1 = S_29; 
		'd30:S_of_i_plus_1 = S_30; 
		'd31:S_of_i_plus_1 = S_31; 
		'd32:S_of_i_plus_1 = S_32; 
		'd33:S_of_i_plus_1 = S_33; 
		'd34:S_of_i_plus_1 = S_34; 
		'd35:S_of_i_plus_1 = S_35; 
		'd36:S_of_i_plus_1 = S_36; 
		'd37:S_of_i_plus_1 = S_37; 
		'd38:S_of_i_plus_1 = S_38; 
		'd39:S_of_i_plus_1 = S_39; 
		'd40:S_of_i_plus_1 = S_40; 
		'd41:S_of_i_plus_1 = S_41; 
		'd42:S_of_i_plus_1 = S_42; 
		'd43:S_of_i_plus_1 = S_43; 
		'd44:S_of_i_plus_1 = S_44; 
		'd45:S_of_i_plus_1 = S_45; 
		'd46:S_of_i_plus_1 = S_46; 
		'd47:S_of_i_plus_1 = S_47; 
		'd48:S_of_i_plus_1 = S_48; 
		'd49:S_of_i_plus_1 = S_49; 
		'd50:S_of_i_plus_1 = S_50; 
		'd51:S_of_i_plus_1 = S_51; 
		'd52:S_of_i_plus_1 = S_52; 
		'd53:S_of_i_plus_1 = S_53; 
		'd54:S_of_i_plus_1 = S_54; 
		'd55:S_of_i_plus_1 = S_55; 
		'd56:S_of_i_plus_1 = S_56; 
		'd57:S_of_i_plus_1 = S_57; 
		'd58:S_of_i_plus_1 = S_58; 
		'd59:S_of_i_plus_1 = S_59; 
		'd60:S_of_i_plus_1 = S_60; 
		'd61:S_of_i_plus_1 = S_61; 
		'd62:S_of_i_plus_1 = S_62; 
		'd63:S_of_i_plus_1 = S_63; 
		'd64:S_of_i_plus_1 = S_64; 
		'd65:S_of_i_plus_1 = S_65; 
		'd66:S_of_i_plus_1 = S_66; 
		'd67:S_of_i_plus_1 = S_67; 
		'd68:S_of_i_plus_1 = S_68; 
		'd69:S_of_i_plus_1 = S_69; 
		'd70:S_of_i_plus_1 = S_70; 
		'd71:S_of_i_plus_1 = S_71; 
		'd72:S_of_i_plus_1 = S_72; 
		'd73:S_of_i_plus_1 = S_73; 
		'd74:S_of_i_plus_1 = S_74; 
		'd75:S_of_i_plus_1 = S_75; 
		'd76:S_of_i_plus_1 = S_76; 
		'd77:S_of_i_plus_1 = S_77; 
		'd78:S_of_i_plus_1 = S_78; 
		'd79:S_of_i_plus_1 = S_79; 
		'd80:S_of_i_plus_1 = S_80; 
		'd81:S_of_i_plus_1 = S_81; 
		'd82:S_of_i_plus_1 = S_82; 
		'd83:S_of_i_plus_1 = S_83; 
		'd84:S_of_i_plus_1 = S_84; 
		'd85:S_of_i_plus_1 = S_85; 
		'd86:S_of_i_plus_1 = S_86; 
		'd87:S_of_i_plus_1 = S_87; 
		'd88:S_of_i_plus_1 = S_88; 
		'd89:S_of_i_plus_1 = S_89; 
		'd90:S_of_i_plus_1 = S_90; 
		'd91:S_of_i_plus_1 = S_91; 
		'd92:S_of_i_plus_1 = S_92; 
		'd93:S_of_i_plus_1 = S_93; 
		'd94:S_of_i_plus_1 = S_94; 
		'd95:S_of_i_plus_1 = S_95; 
		'd96:S_of_i_plus_1 = S_96; 
		'd97:S_of_i_plus_1 = S_97; 
		'd98:S_of_i_plus_1 = S_98; 
		'd99:S_of_i_plus_1 = S_99; 
		'd100:S_of_i_plus_1 = S_100; 
		'd101:S_of_i_plus_1 = S_101; 
		'd102:S_of_i_plus_1 = S_102; 
		'd103:S_of_i_plus_1 = S_103; 
		'd104:S_of_i_plus_1 = S_104; 
		'd105:S_of_i_plus_1 = S_105; 
		'd106:S_of_i_plus_1 = S_106; 
		'd107:S_of_i_plus_1 = S_107; 
		'd108:S_of_i_plus_1 = S_108; 
		'd109:S_of_i_plus_1 = S_109; 
		'd110:S_of_i_plus_1 = S_110; 
		'd111:S_of_i_plus_1 = S_111; 
		'd112:S_of_i_plus_1 = S_112; 
		'd113:S_of_i_plus_1 = S_113; 
		'd114:S_of_i_plus_1 = S_114; 
		'd115:S_of_i_plus_1 = S_115; 
		'd116:S_of_i_plus_1 = S_116; 
		'd117:S_of_i_plus_1 = S_117; 
		'd118:S_of_i_plus_1 = S_118; 
		'd119:S_of_i_plus_1 = S_119; 
		'd120:S_of_i_plus_1 = S_120; 
		'd121:S_of_i_plus_1 = S_121; 
		'd122:S_of_i_plus_1 = S_122; 
		'd123:S_of_i_plus_1 = S_123; 
		'd124:S_of_i_plus_1 = S_124; 
		'd125:S_of_i_plus_1 = S_125; 
		'd126:S_of_i_plus_1 = S_126; 
		'd127:S_of_i_plus_1 = S_127; 
		'd128:S_of_i_plus_1 = S_128; 
		'd129:S_of_i_plus_1 = S_129; 
		'd130:S_of_i_plus_1 = S_130; 
		'd131:S_of_i_plus_1 = S_131; 
		'd132:S_of_i_plus_1 = S_132; 
		'd133:S_of_i_plus_1 = S_133; 
		'd134:S_of_i_plus_1 = S_134; 
		'd135:S_of_i_plus_1 = S_135; 
		'd136:S_of_i_plus_1 = S_136; 
		'd137:S_of_i_plus_1 = S_137; 
		'd138:S_of_i_plus_1 = S_138; 
		'd139:S_of_i_plus_1 = S_139; 
		'd140:S_of_i_plus_1 = S_140; 
		'd141:S_of_i_plus_1 = S_141; 
		'd142:S_of_i_plus_1 = S_142; 
		'd143:S_of_i_plus_1 = S_143; 
		'd144:S_of_i_plus_1 = S_144; 
		'd145:S_of_i_plus_1 = S_145; 
		'd146:S_of_i_plus_1 = S_146; 
		'd147:S_of_i_plus_1 = S_147; 
		'd148:S_of_i_plus_1 = S_148; 
		'd149:S_of_i_plus_1 = S_149; 
		'd150:S_of_i_plus_1 = S_150; 
		'd151:S_of_i_plus_1 = S_151; 
		'd152:S_of_i_plus_1 = S_152; 
		'd153:S_of_i_plus_1 = S_153; 
		'd154:S_of_i_plus_1 = S_154; 
		'd155:S_of_i_plus_1 = S_155; 
		'd156:S_of_i_plus_1 = S_156; 
		'd157:S_of_i_plus_1 = S_157; 
		'd158:S_of_i_plus_1 = S_158; 
		'd159:S_of_i_plus_1 = S_159; 
		'd160:S_of_i_plus_1 = S_160; 
		'd161:S_of_i_plus_1 = S_161; 
		'd162:S_of_i_plus_1 = S_162; 
		'd163:S_of_i_plus_1 = S_163; 
		'd164:S_of_i_plus_1 = S_164; 
		'd165:S_of_i_plus_1 = S_165; 
		'd166:S_of_i_plus_1 = S_166; 
		'd167:S_of_i_plus_1 = S_167; 
		'd168:S_of_i_plus_1 = S_168; 
		'd169:S_of_i_plus_1 = S_169; 
		'd170:S_of_i_plus_1 = S_170; 
		'd171:S_of_i_plus_1 = S_171; 
		'd172:S_of_i_plus_1 = S_172; 
		'd173:S_of_i_plus_1 = S_173; 
		'd174:S_of_i_plus_1 = S_174; 
		'd175:S_of_i_plus_1 = S_175; 
		'd176:S_of_i_plus_1 = S_176; 
		'd177:S_of_i_plus_1 = S_177; 
		'd178:S_of_i_plus_1 = S_178; 
		'd179:S_of_i_plus_1 = S_179; 
		'd180:S_of_i_plus_1 = S_180; 
		'd181:S_of_i_plus_1 = S_181; 
		'd182:S_of_i_plus_1 = S_182; 
		'd183:S_of_i_plus_1 = S_183; 
		'd184:S_of_i_plus_1 = S_184; 
		'd185:S_of_i_plus_1 = S_185; 
		'd186:S_of_i_plus_1 = S_186; 
		'd187:S_of_i_plus_1 = S_187; 
		'd188:S_of_i_plus_1 = S_188; 
		'd189:S_of_i_plus_1 = S_189; 
		'd190:S_of_i_plus_1 = S_190; 
		'd191:S_of_i_plus_1 = S_191; 
		'd192:S_of_i_plus_1 = S_192; 
		'd193:S_of_i_plus_1 = S_193; 
		'd194:S_of_i_plus_1 = S_194; 
		'd195:S_of_i_plus_1 = S_195; 
		'd196:S_of_i_plus_1 = S_196; 
		'd197:S_of_i_plus_1 = S_197; 
		'd198:S_of_i_plus_1 = S_198; 
		'd199:S_of_i_plus_1 = S_199; 
		'd200:S_of_i_plus_1 = S_200; 
		'd201:S_of_i_plus_1 = S_201; 
		'd202:S_of_i_plus_1 = S_202; 
		'd203:S_of_i_plus_1 = S_203; 
		'd204:S_of_i_plus_1 = S_204; 
		'd205:S_of_i_plus_1 = S_205; 
		'd206:S_of_i_plus_1 = S_206; 
		'd207:S_of_i_plus_1 = S_207; 
		'd208:S_of_i_plus_1 = S_208; 
		'd209:S_of_i_plus_1 = S_209; 
		'd210:S_of_i_plus_1 = S_210; 
		'd211:S_of_i_plus_1 = S_211; 
		'd212:S_of_i_plus_1 = S_212; 
		'd213:S_of_i_plus_1 = S_213; 
		'd214:S_of_i_plus_1 = S_214; 
		'd215:S_of_i_plus_1 = S_215; 
		'd216:S_of_i_plus_1 = S_216; 
		'd217:S_of_i_plus_1 = S_217; 
		'd218:S_of_i_plus_1 = S_218; 
		'd219:S_of_i_plus_1 = S_219; 
		'd220:S_of_i_plus_1 = S_220; 
		'd221:S_of_i_plus_1 = S_221; 
		'd222:S_of_i_plus_1 = S_222; 
		'd223:S_of_i_plus_1 = S_223; 
		'd224:S_of_i_plus_1 = S_224; 
		'd225:S_of_i_plus_1 = S_225; 
		'd226:S_of_i_plus_1 = S_226; 
		'd227:S_of_i_plus_1 = S_227; 
		'd228:S_of_i_plus_1 = S_228; 
		'd229:S_of_i_plus_1 = S_229; 
		'd230:S_of_i_plus_1 = S_230; 
		'd231:S_of_i_plus_1 = S_231; 
		'd232:S_of_i_plus_1 = S_232; 
		'd233:S_of_i_plus_1 = S_233; 
		'd234:S_of_i_plus_1 = S_234; 
		'd235:S_of_i_plus_1 = S_235; 
		'd236:S_of_i_plus_1 = S_236; 
		'd237:S_of_i_plus_1 = S_237; 
		'd238:S_of_i_plus_1 = S_238; 
		'd239:S_of_i_plus_1 = S_239; 
		'd240:S_of_i_plus_1 = S_240; 
		'd241:S_of_i_plus_1 = S_241; 
		'd242:S_of_i_plus_1 = S_242; 
		'd243:S_of_i_plus_1 = S_243; 
		'd244:S_of_i_plus_1 = S_244; 
		'd245:S_of_i_plus_1 = S_245; 
		'd246:S_of_i_plus_1 = S_246; 
		'd247:S_of_i_plus_1 = S_247; 
		'd248:S_of_i_plus_1 = S_248; 
		'd249:S_of_i_plus_1 = S_249; 
		'd250:S_of_i_plus_1 = S_250; 
		'd251:S_of_i_plus_1 = S_251; 
		'd252:S_of_i_plus_1 = S_252; 
		'd253:S_of_i_plus_1 = S_253; 
		'd254:S_of_i_plus_1 = S_254; 
		'd255:S_of_i_plus_1 = S_255; 
		default:S_of_i_plus_1 = S_256; 
	endcase
end
always @ (j or S_0 or S_1 or S_2 or S_3 or S_4 or S_5 or S_6 or S_7 or S_8 or S_9 or S_10 or S_11 or S_12 or S_13 or S_14 or S_15 or S_16 or S_17 or S_18 or S_19 or S_20 or S_21 or S_22 or S_23 or S_24 or S_25 or S_26 or S_27 or S_28 or S_29 or S_30 or S_31 or S_32 or S_33 or S_34 or S_35 or S_36 or S_37 or S_38 or S_39 or S_40 or S_41 or S_42 or S_43 or S_44 or S_45 or S_46 or S_47 or S_48 or S_49 or S_50 or S_51 or S_52 or S_53 or S_54 or S_55 or S_56 or S_57 or S_58 or S_59 or S_60 or S_61 or S_62 or S_63 or S_64 or S_65 or S_66 or S_67 or S_68 or S_69 or S_70 or S_71 or S_72 or S_73 or S_74 or S_75 or S_76 or S_77 or S_78 or S_79 or S_80 or S_81 or S_82 or S_83 or S_84 or S_85 or S_86 or S_87 or S_88 or S_89 or S_90 or S_91 or S_92 or S_93 or S_94 or S_95 or S_96 or S_97 or S_98 or S_99 or S_100 or S_101 or S_102 or S_103 or S_104 or S_105 or S_106 or S_107 or S_108 or S_109 or S_110 or S_111 or S_112 or S_113 or S_114 or S_115 or S_116 or S_117 or S_118 or S_119 or S_120 or S_121 or S_122 or S_123 or S_124 or S_125 or S_126 or S_127 or S_128 or S_129 or S_130 or S_131 or S_132 or S_133 or S_134 or S_135 or S_136 or S_137 or S_138 or S_139 or S_140 or S_141 or S_142 or S_143 or S_144 or S_145 or S_146 or S_147 or S_148 or S_149 or S_150 or S_151 or S_152 or S_153 or S_154 or S_155 or S_156 or S_157 or S_158 or S_159 or S_160 or S_161 or S_162 or S_163 or S_164 or S_165 or S_166 or S_167 or S_168 or S_169 or S_170 or S_171 or S_172 or S_173 or S_174 or S_175 or S_176 or S_177 or S_178 or S_179 or S_180 or S_181 or S_182 or S_183 or S_184 or S_185 or S_186 or S_187 or S_188 or S_189 or S_190 or S_191 or S_192 or S_193 or S_194 or S_195 or S_196 or S_197 or S_198 or S_199 or S_200 or S_201 or S_202 or S_203 or S_204 or S_205 or S_206 or S_207 or S_208 or S_209 or S_210 or S_211 or S_212 or S_213 or S_214 or S_215 or S_216 or S_217 or S_218 or S_219 or S_220 or S_221 or S_222 or S_223 or S_224 or S_225 or S_226 or S_227 or S_228 or S_229 or S_230 or S_231 or S_232 or S_233 or S_234 or S_235 or S_236 or S_237 or S_238 or S_239 or S_240 or S_241 or S_242 or S_243 or S_244 or S_245 or S_246 or S_247 or S_248 or S_249 or S_250 or S_251 or S_252 or S_253 or S_254 or S_255) begin
	case (j) 
		'd0:S_of_j = S_0; 
		'd1:S_of_j = S_1; 
		'd2:S_of_j = S_2; 
		'd3:S_of_j = S_3; 
		'd4:S_of_j = S_4; 
		'd5:S_of_j = S_5; 
		'd6:S_of_j = S_6; 
		'd7:S_of_j = S_7; 
		'd8:S_of_j = S_8; 
		'd9:S_of_j = S_9; 
		'd10:S_of_j = S_10; 
		'd11:S_of_j = S_11; 
		'd12:S_of_j = S_12; 
		'd13:S_of_j = S_13; 
		'd14:S_of_j = S_14; 
		'd15:S_of_j = S_15; 
		'd16:S_of_j = S_16; 
		'd17:S_of_j = S_17; 
		'd18:S_of_j = S_18; 
		'd19:S_of_j = S_19; 
		'd20:S_of_j = S_20; 
		'd21:S_of_j = S_21; 
		'd22:S_of_j = S_22; 
		'd23:S_of_j = S_23; 
		'd24:S_of_j = S_24; 
		'd25:S_of_j = S_25; 
		'd26:S_of_j = S_26; 
		'd27:S_of_j = S_27; 
		'd28:S_of_j = S_28; 
		'd29:S_of_j = S_29; 
		'd30:S_of_j = S_30; 
		'd31:S_of_j = S_31; 
		'd32:S_of_j = S_32; 
		'd33:S_of_j = S_33; 
		'd34:S_of_j = S_34; 
		'd35:S_of_j = S_35; 
		'd36:S_of_j = S_36; 
		'd37:S_of_j = S_37; 
		'd38:S_of_j = S_38; 
		'd39:S_of_j = S_39; 
		'd40:S_of_j = S_40; 
		'd41:S_of_j = S_41; 
		'd42:S_of_j = S_42; 
		'd43:S_of_j = S_43; 
		'd44:S_of_j = S_44; 
		'd45:S_of_j = S_45; 
		'd46:S_of_j = S_46; 
		'd47:S_of_j = S_47; 
		'd48:S_of_j = S_48; 
		'd49:S_of_j = S_49; 
		'd50:S_of_j = S_50; 
		'd51:S_of_j = S_51; 
		'd52:S_of_j = S_52; 
		'd53:S_of_j = S_53; 
		'd54:S_of_j = S_54; 
		'd55:S_of_j = S_55; 
		'd56:S_of_j = S_56; 
		'd57:S_of_j = S_57; 
		'd58:S_of_j = S_58; 
		'd59:S_of_j = S_59; 
		'd60:S_of_j = S_60; 
		'd61:S_of_j = S_61; 
		'd62:S_of_j = S_62; 
		'd63:S_of_j = S_63; 
		'd64:S_of_j = S_64; 
		'd65:S_of_j = S_65; 
		'd66:S_of_j = S_66; 
		'd67:S_of_j = S_67; 
		'd68:S_of_j = S_68; 
		'd69:S_of_j = S_69; 
		'd70:S_of_j = S_70; 
		'd71:S_of_j = S_71; 
		'd72:S_of_j = S_72; 
		'd73:S_of_j = S_73; 
		'd74:S_of_j = S_74; 
		'd75:S_of_j = S_75; 
		'd76:S_of_j = S_76; 
		'd77:S_of_j = S_77; 
		'd78:S_of_j = S_78; 
		'd79:S_of_j = S_79; 
		'd80:S_of_j = S_80; 
		'd81:S_of_j = S_81; 
		'd82:S_of_j = S_82; 
		'd83:S_of_j = S_83; 
		'd84:S_of_j = S_84; 
		'd85:S_of_j = S_85; 
		'd86:S_of_j = S_86; 
		'd87:S_of_j = S_87; 
		'd88:S_of_j = S_88; 
		'd89:S_of_j = S_89; 
		'd90:S_of_j = S_90; 
		'd91:S_of_j = S_91; 
		'd92:S_of_j = S_92; 
		'd93:S_of_j = S_93; 
		'd94:S_of_j = S_94; 
		'd95:S_of_j = S_95; 
		'd96:S_of_j = S_96; 
		'd97:S_of_j = S_97; 
		'd98:S_of_j = S_98; 
		'd99:S_of_j = S_99; 
		'd100:S_of_j = S_100; 
		'd101:S_of_j = S_101; 
		'd102:S_of_j = S_102; 
		'd103:S_of_j = S_103; 
		'd104:S_of_j = S_104; 
		'd105:S_of_j = S_105; 
		'd106:S_of_j = S_106; 
		'd107:S_of_j = S_107; 
		'd108:S_of_j = S_108; 
		'd109:S_of_j = S_109; 
		'd110:S_of_j = S_110; 
		'd111:S_of_j = S_111; 
		'd112:S_of_j = S_112; 
		'd113:S_of_j = S_113; 
		'd114:S_of_j = S_114; 
		'd115:S_of_j = S_115; 
		'd116:S_of_j = S_116; 
		'd117:S_of_j = S_117; 
		'd118:S_of_j = S_118; 
		'd119:S_of_j = S_119; 
		'd120:S_of_j = S_120; 
		'd121:S_of_j = S_121; 
		'd122:S_of_j = S_122; 
		'd123:S_of_j = S_123; 
		'd124:S_of_j = S_124; 
		'd125:S_of_j = S_125; 
		'd126:S_of_j = S_126; 
		'd127:S_of_j = S_127; 
		'd128:S_of_j = S_128; 
		'd129:S_of_j = S_129; 
		'd130:S_of_j = S_130; 
		'd131:S_of_j = S_131; 
		'd132:S_of_j = S_132; 
		'd133:S_of_j = S_133; 
		'd134:S_of_j = S_134; 
		'd135:S_of_j = S_135; 
		'd136:S_of_j = S_136; 
		'd137:S_of_j = S_137; 
		'd138:S_of_j = S_138; 
		'd139:S_of_j = S_139; 
		'd140:S_of_j = S_140; 
		'd141:S_of_j = S_141; 
		'd142:S_of_j = S_142; 
		'd143:S_of_j = S_143; 
		'd144:S_of_j = S_144; 
		'd145:S_of_j = S_145; 
		'd146:S_of_j = S_146; 
		'd147:S_of_j = S_147; 
		'd148:S_of_j = S_148; 
		'd149:S_of_j = S_149; 
		'd150:S_of_j = S_150; 
		'd151:S_of_j = S_151; 
		'd152:S_of_j = S_152; 
		'd153:S_of_j = S_153; 
		'd154:S_of_j = S_154; 
		'd155:S_of_j = S_155; 
		'd156:S_of_j = S_156; 
		'd157:S_of_j = S_157; 
		'd158:S_of_j = S_158; 
		'd159:S_of_j = S_159; 
		'd160:S_of_j = S_160; 
		'd161:S_of_j = S_161; 
		'd162:S_of_j = S_162; 
		'd163:S_of_j = S_163; 
		'd164:S_of_j = S_164; 
		'd165:S_of_j = S_165; 
		'd166:S_of_j = S_166; 
		'd167:S_of_j = S_167; 
		'd168:S_of_j = S_168; 
		'd169:S_of_j = S_169; 
		'd170:S_of_j = S_170; 
		'd171:S_of_j = S_171; 
		'd172:S_of_j = S_172; 
		'd173:S_of_j = S_173; 
		'd174:S_of_j = S_174; 
		'd175:S_of_j = S_175; 
		'd176:S_of_j = S_176; 
		'd177:S_of_j = S_177; 
		'd178:S_of_j = S_178; 
		'd179:S_of_j = S_179; 
		'd180:S_of_j = S_180; 
		'd181:S_of_j = S_181; 
		'd182:S_of_j = S_182; 
		'd183:S_of_j = S_183; 
		'd184:S_of_j = S_184; 
		'd185:S_of_j = S_185; 
		'd186:S_of_j = S_186; 
		'd187:S_of_j = S_187; 
		'd188:S_of_j = S_188; 
		'd189:S_of_j = S_189; 
		'd190:S_of_j = S_190; 
		'd191:S_of_j = S_191; 
		'd192:S_of_j = S_192; 
		'd193:S_of_j = S_193; 
		'd194:S_of_j = S_194; 
		'd195:S_of_j = S_195; 
		'd196:S_of_j = S_196; 
		'd197:S_of_j = S_197; 
		'd198:S_of_j = S_198; 
		'd199:S_of_j = S_199; 
		'd200:S_of_j = S_200; 
		'd201:S_of_j = S_201; 
		'd202:S_of_j = S_202; 
		'd203:S_of_j = S_203; 
		'd204:S_of_j = S_204; 
		'd205:S_of_j = S_205; 
		'd206:S_of_j = S_206; 
		'd207:S_of_j = S_207; 
		'd208:S_of_j = S_208; 
		'd209:S_of_j = S_209; 
		'd210:S_of_j = S_210; 
		'd211:S_of_j = S_211; 
		'd212:S_of_j = S_212; 
		'd213:S_of_j = S_213; 
		'd214:S_of_j = S_214; 
		'd215:S_of_j = S_215; 
		'd216:S_of_j = S_216; 
		'd217:S_of_j = S_217; 
		'd218:S_of_j = S_218; 
		'd219:S_of_j = S_219; 
		'd220:S_of_j = S_220; 
		'd221:S_of_j = S_221; 
		'd222:S_of_j = S_222; 
		'd223:S_of_j = S_223; 
		'd224:S_of_j = S_224; 
		'd225:S_of_j = S_225; 
		'd226:S_of_j = S_226; 
		'd227:S_of_j = S_227; 
		'd228:S_of_j = S_228; 
		'd229:S_of_j = S_229; 
		'd230:S_of_j = S_230; 
		'd231:S_of_j = S_231; 
		'd232:S_of_j = S_232; 
		'd233:S_of_j = S_233; 
		'd234:S_of_j = S_234; 
		'd235:S_of_j = S_235; 
		'd236:S_of_j = S_236; 
		'd237:S_of_j = S_237; 
		'd238:S_of_j = S_238; 
		'd239:S_of_j = S_239; 
		'd240:S_of_j = S_240; 
		'd241:S_of_j = S_241; 
		'd242:S_of_j = S_242; 
		'd243:S_of_j = S_243; 
		'd244:S_of_j = S_244; 
		'd245:S_of_j = S_245; 
		'd246:S_of_j = S_246; 
		'd247:S_of_j = S_247; 
		'd248:S_of_j = S_248; 
		'd249:S_of_j = S_249; 
		'd250:S_of_j = S_250; 
		'd251:S_of_j = S_251; 
		'd252:S_of_j = S_252; 
		'd253:S_of_j = S_253; 
		'd254:S_of_j = S_254; 
		default:S_of_j = S_255; 
	endcase
end
always @ (i_mod_KEYSIZE or key_0 or key_1 or key_2 or key_3 or key_4 or key_5 or key_6) begin
	case (i_mod_KEYSIZE) 
		'd0:key_of_i_mod_KEYSIZE = key_0; 
		'd1:key_of_i_mod_KEYSIZE = key_1; 
		'd2:key_of_i_mod_KEYSIZE = key_2; 
		'd3:key_of_i_mod_KEYSIZE = key_3; 
		'd4:key_of_i_mod_KEYSIZE = key_4; 
		'd5:key_of_i_mod_KEYSIZE = key_5; 
		default:key_of_i_mod_KEYSIZE = key_6; 
	endcase
end
always @ (i) begin
	case (i) 
		'd0: i_mod_KEYSIZE = 0; 
		'd1: i_mod_KEYSIZE = 1; 
		'd2: i_mod_KEYSIZE = 2; 
		'd3: i_mod_KEYSIZE = 3; 
		'd4: i_mod_KEYSIZE = 4; 
		'd5: i_mod_KEYSIZE = 5; 
		'd6: i_mod_KEYSIZE = 6; 
		'd7: i_mod_KEYSIZE = 0; 
		'd8: i_mod_KEYSIZE = 1; 
		'd9: i_mod_KEYSIZE = 2; 
		'd10: i_mod_KEYSIZE = 3; 
		'd11: i_mod_KEYSIZE = 4; 
		'd12: i_mod_KEYSIZE = 5; 
		'd13: i_mod_KEYSIZE = 6; 
		'd14: i_mod_KEYSIZE = 0; 
		'd15: i_mod_KEYSIZE = 1; 
		'd16: i_mod_KEYSIZE = 2; 
		'd17: i_mod_KEYSIZE = 3; 
		'd18: i_mod_KEYSIZE = 4; 
		'd19: i_mod_KEYSIZE = 5; 
		'd20: i_mod_KEYSIZE = 6; 
		'd21: i_mod_KEYSIZE = 0; 
		'd22: i_mod_KEYSIZE = 1; 
		'd23: i_mod_KEYSIZE = 2; 
		'd24: i_mod_KEYSIZE = 3; 
		'd25: i_mod_KEYSIZE = 4; 
		'd26: i_mod_KEYSIZE = 5; 
		'd27: i_mod_KEYSIZE = 6; 
		'd28: i_mod_KEYSIZE = 0; 
		'd29: i_mod_KEYSIZE = 1; 
		'd30: i_mod_KEYSIZE = 2; 
		'd31: i_mod_KEYSIZE = 3; 
		'd32: i_mod_KEYSIZE = 4; 
		'd33: i_mod_KEYSIZE = 5; 
		'd34: i_mod_KEYSIZE = 6; 
		'd35: i_mod_KEYSIZE = 0; 
		'd36: i_mod_KEYSIZE = 1; 
		'd37: i_mod_KEYSIZE = 2; 
		'd38: i_mod_KEYSIZE = 3; 
		'd39: i_mod_KEYSIZE = 4; 
		'd40: i_mod_KEYSIZE = 5; 
		'd41: i_mod_KEYSIZE = 6; 
		'd42: i_mod_KEYSIZE = 0; 
		'd43: i_mod_KEYSIZE = 1; 
		'd44: i_mod_KEYSIZE = 2; 
		'd45: i_mod_KEYSIZE = 3; 
		'd46: i_mod_KEYSIZE = 4; 
		'd47: i_mod_KEYSIZE = 5; 
		'd48: i_mod_KEYSIZE = 6; 
		'd49: i_mod_KEYSIZE = 0; 
		'd50: i_mod_KEYSIZE = 1; 
		'd51: i_mod_KEYSIZE = 2; 
		'd52: i_mod_KEYSIZE = 3; 
		'd53: i_mod_KEYSIZE = 4; 
		'd54: i_mod_KEYSIZE = 5; 
		'd55: i_mod_KEYSIZE = 6; 
		'd56: i_mod_KEYSIZE = 0; 
		'd57: i_mod_KEYSIZE = 1; 
		'd58: i_mod_KEYSIZE = 2; 
		'd59: i_mod_KEYSIZE = 3; 
		'd60: i_mod_KEYSIZE = 4; 
		'd61: i_mod_KEYSIZE = 5; 
		'd62: i_mod_KEYSIZE = 6; 
		'd63: i_mod_KEYSIZE = 0; 
		'd64: i_mod_KEYSIZE = 1; 
		'd65: i_mod_KEYSIZE = 2; 
		'd66: i_mod_KEYSIZE = 3; 
		'd67: i_mod_KEYSIZE = 4; 
		'd68: i_mod_KEYSIZE = 5; 
		'd69: i_mod_KEYSIZE = 6; 
		'd70: i_mod_KEYSIZE = 0; 
		'd71: i_mod_KEYSIZE = 1; 
		'd72: i_mod_KEYSIZE = 2; 
		'd73: i_mod_KEYSIZE = 3; 
		'd74: i_mod_KEYSIZE = 4; 
		'd75: i_mod_KEYSIZE = 5; 
		'd76: i_mod_KEYSIZE = 6; 
		'd77: i_mod_KEYSIZE = 0; 
		'd78: i_mod_KEYSIZE = 1; 
		'd79: i_mod_KEYSIZE = 2; 
		'd80: i_mod_KEYSIZE = 3; 
		'd81: i_mod_KEYSIZE = 4; 
		'd82: i_mod_KEYSIZE = 5; 
		'd83: i_mod_KEYSIZE = 6; 
		'd84: i_mod_KEYSIZE = 0; 
		'd85: i_mod_KEYSIZE = 1; 
		'd86: i_mod_KEYSIZE = 2; 
		'd87: i_mod_KEYSIZE = 3; 
		'd88: i_mod_KEYSIZE = 4; 
		'd89: i_mod_KEYSIZE = 5; 
		'd90: i_mod_KEYSIZE = 6; 
		'd91: i_mod_KEYSIZE = 0; 
		'd92: i_mod_KEYSIZE = 1; 
		'd93: i_mod_KEYSIZE = 2; 
		'd94: i_mod_KEYSIZE = 3; 
		'd95: i_mod_KEYSIZE = 4; 
		'd96: i_mod_KEYSIZE = 5; 
		'd97: i_mod_KEYSIZE = 6; 
		'd98: i_mod_KEYSIZE = 0; 
		'd99: i_mod_KEYSIZE = 1; 
		'd100: i_mod_KEYSIZE = 2; 
		'd101: i_mod_KEYSIZE = 3; 
		'd102: i_mod_KEYSIZE = 4; 
		'd103: i_mod_KEYSIZE = 5; 
		'd104: i_mod_KEYSIZE = 6; 
		'd105: i_mod_KEYSIZE = 0; 
		'd106: i_mod_KEYSIZE = 1; 
		'd107: i_mod_KEYSIZE = 2; 
		'd108: i_mod_KEYSIZE = 3; 
		'd109: i_mod_KEYSIZE = 4; 
		'd110: i_mod_KEYSIZE = 5; 
		'd111: i_mod_KEYSIZE = 6; 
		'd112: i_mod_KEYSIZE = 0; 
		'd113: i_mod_KEYSIZE = 1; 
		'd114: i_mod_KEYSIZE = 2; 
		'd115: i_mod_KEYSIZE = 3; 
		'd116: i_mod_KEYSIZE = 4; 
		'd117: i_mod_KEYSIZE = 5; 
		'd118: i_mod_KEYSIZE = 6; 
		'd119: i_mod_KEYSIZE = 0; 
		'd120: i_mod_KEYSIZE = 1; 
		'd121: i_mod_KEYSIZE = 2; 
		'd122: i_mod_KEYSIZE = 3; 
		'd123: i_mod_KEYSIZE = 4; 
		'd124: i_mod_KEYSIZE = 5; 
		'd125: i_mod_KEYSIZE = 6; 
		'd126: i_mod_KEYSIZE = 0; 
		'd127: i_mod_KEYSIZE = 1; 
		'd128: i_mod_KEYSIZE = 2; 
		'd129: i_mod_KEYSIZE = 3; 
		'd130: i_mod_KEYSIZE = 4; 
		'd131: i_mod_KEYSIZE = 5; 
		'd132: i_mod_KEYSIZE = 6; 
		'd133: i_mod_KEYSIZE = 0; 
		'd134: i_mod_KEYSIZE = 1; 
		'd135: i_mod_KEYSIZE = 2; 
		'd136: i_mod_KEYSIZE = 3; 
		'd137: i_mod_KEYSIZE = 4; 
		'd138: i_mod_KEYSIZE = 5; 
		'd139: i_mod_KEYSIZE = 6; 
		'd140: i_mod_KEYSIZE = 0; 
		'd141: i_mod_KEYSIZE = 1; 
		'd142: i_mod_KEYSIZE = 2; 
		'd143: i_mod_KEYSIZE = 3; 
		'd144: i_mod_KEYSIZE = 4; 
		'd145: i_mod_KEYSIZE = 5; 
		'd146: i_mod_KEYSIZE = 6; 
		'd147: i_mod_KEYSIZE = 0; 
		'd148: i_mod_KEYSIZE = 1; 
		'd149: i_mod_KEYSIZE = 2; 
		'd150: i_mod_KEYSIZE = 3; 
		'd151: i_mod_KEYSIZE = 4; 
		'd152: i_mod_KEYSIZE = 5; 
		'd153: i_mod_KEYSIZE = 6; 
		'd154: i_mod_KEYSIZE = 0; 
		'd155: i_mod_KEYSIZE = 1; 
		'd156: i_mod_KEYSIZE = 2; 
		'd157: i_mod_KEYSIZE = 3; 
		'd158: i_mod_KEYSIZE = 4; 
		'd159: i_mod_KEYSIZE = 5; 
		'd160: i_mod_KEYSIZE = 6; 
		'd161: i_mod_KEYSIZE = 0; 
		'd162: i_mod_KEYSIZE = 1; 
		'd163: i_mod_KEYSIZE = 2; 
		'd164: i_mod_KEYSIZE = 3; 
		'd165: i_mod_KEYSIZE = 4; 
		'd166: i_mod_KEYSIZE = 5; 
		'd167: i_mod_KEYSIZE = 6; 
		'd168: i_mod_KEYSIZE = 0; 
		'd169: i_mod_KEYSIZE = 1; 
		'd170: i_mod_KEYSIZE = 2; 
		'd171: i_mod_KEYSIZE = 3; 
		'd172: i_mod_KEYSIZE = 4; 
		'd173: i_mod_KEYSIZE = 5; 
		'd174: i_mod_KEYSIZE = 6; 
		'd175: i_mod_KEYSIZE = 0; 
		'd176: i_mod_KEYSIZE = 1; 
		'd177: i_mod_KEYSIZE = 2; 
		'd178: i_mod_KEYSIZE = 3; 
		'd179: i_mod_KEYSIZE = 4; 
		'd180: i_mod_KEYSIZE = 5; 
		'd181: i_mod_KEYSIZE = 6; 
		'd182: i_mod_KEYSIZE = 0; 
		'd183: i_mod_KEYSIZE = 1; 
		'd184: i_mod_KEYSIZE = 2; 
		'd185: i_mod_KEYSIZE = 3; 
		'd186: i_mod_KEYSIZE = 4; 
		'd187: i_mod_KEYSIZE = 5; 
		'd188: i_mod_KEYSIZE = 6; 
		'd189: i_mod_KEYSIZE = 0; 
		'd190: i_mod_KEYSIZE = 1; 
		'd191: i_mod_KEYSIZE = 2; 
		'd192: i_mod_KEYSIZE = 3; 
		'd193: i_mod_KEYSIZE = 4; 
		'd194: i_mod_KEYSIZE = 5; 
		'd195: i_mod_KEYSIZE = 6; 
		'd196: i_mod_KEYSIZE = 0; 
		'd197: i_mod_KEYSIZE = 1; 
		'd198: i_mod_KEYSIZE = 2; 
		'd199: i_mod_KEYSIZE = 3; 
		'd200: i_mod_KEYSIZE = 4; 
		'd201: i_mod_KEYSIZE = 5; 
		'd202: i_mod_KEYSIZE = 6; 
		'd203: i_mod_KEYSIZE = 0; 
		'd204: i_mod_KEYSIZE = 1; 
		'd205: i_mod_KEYSIZE = 2; 
		'd206: i_mod_KEYSIZE = 3; 
		'd207: i_mod_KEYSIZE = 4; 
		'd208: i_mod_KEYSIZE = 5; 
		'd209: i_mod_KEYSIZE = 6; 
		'd210: i_mod_KEYSIZE = 0; 
		'd211: i_mod_KEYSIZE = 1; 
		'd212: i_mod_KEYSIZE = 2; 
		'd213: i_mod_KEYSIZE = 3; 
		'd214: i_mod_KEYSIZE = 4; 
		'd215: i_mod_KEYSIZE = 5; 
		'd216: i_mod_KEYSIZE = 6; 
		'd217: i_mod_KEYSIZE = 0; 
		'd218: i_mod_KEYSIZE = 1; 
		'd219: i_mod_KEYSIZE = 2; 
		'd220: i_mod_KEYSIZE = 3; 
		'd221: i_mod_KEYSIZE = 4; 
		'd222: i_mod_KEYSIZE = 5; 
		'd223: i_mod_KEYSIZE = 6; 
		'd224: i_mod_KEYSIZE = 0; 
		'd225: i_mod_KEYSIZE = 1; 
		'd226: i_mod_KEYSIZE = 2; 
		'd227: i_mod_KEYSIZE = 3; 
		'd228: i_mod_KEYSIZE = 4; 
		'd229: i_mod_KEYSIZE = 5; 
		'd230: i_mod_KEYSIZE = 6; 
		'd231: i_mod_KEYSIZE = 0; 
		'd232: i_mod_KEYSIZE = 1; 
		'd233: i_mod_KEYSIZE = 2; 
		'd234: i_mod_KEYSIZE = 3; 
		'd235: i_mod_KEYSIZE = 4; 
		'd236: i_mod_KEYSIZE = 5; 
		'd237: i_mod_KEYSIZE = 6; 
		'd238: i_mod_KEYSIZE = 0; 
		'd239: i_mod_KEYSIZE = 1; 
		'd240: i_mod_KEYSIZE = 2; 
		'd241: i_mod_KEYSIZE = 3; 
		'd242: i_mod_KEYSIZE = 4; 
		'd243: i_mod_KEYSIZE = 5; 
		'd244: i_mod_KEYSIZE = 6; 
		'd245: i_mod_KEYSIZE = 0; 
		'd246: i_mod_KEYSIZE = 1; 
		'd247: i_mod_KEYSIZE = 2; 
		'd248: i_mod_KEYSIZE = 3; 
		'd249: i_mod_KEYSIZE = 4; 
		'd250: i_mod_KEYSIZE = 5; 
		'd251: i_mod_KEYSIZE = 6; 
		'd252: i_mod_KEYSIZE = 0; 
		'd253: i_mod_KEYSIZE = 1; 
		'd254: i_mod_KEYSIZE = 2; 
		'd255: i_mod_KEYSIZE = 3; 
	endcase
end

assign S_of_i_plus_S_of_j = S_of_i + S_of_j;

always @ (posedge clk or posedge rst) begin
	if (rst) begin
		i <= 8'h0;
		KSState <= 4'h0;
		output_ready <= 0;
		j <= 0;
	end else begin
		prev_i <= i;
		prev_S_of_j <= S_of_j;
		case (KSState)
			4'h0: begin // KSS_KEYREAD state: Read key from input
				if (i == 7) begin
					KSState <= 4'h1;
					i<=8'h00;
				end else begin
					i <= i+1;
					// in place of:
					// key[i] <= password_input;
					case (i) 
		'd0:key_0 <= password_input; 
		'd1:key_1 <= password_input; 
		'd2:key_2 <= password_input; 
		'd3:key_3 <= password_input; 
		'd4:key_4 <= password_input; 
		'd5:key_5 <= password_input; 
		default:key_6 <= password_input; 
	endcase
					// $display ("rc4: key[%d] = %08X",i,password_input);
				end
			end

	// for i from 0 to 255
	//     S[i] := i
	// endfor

			4'h1: begin // KSS_KEYSCHED1: Increment counter for S initialization
				// in place of S[i] <= i;
				case (i) 
		'd0:S_0 <= i; 
		'd1:S_1 <= i; 
		'd2:S_2 <= i; 
		'd3:S_3 <= i; 
		'd4:S_4 <= i; 
		'd5:S_5 <= i; 
		'd6:S_6 <= i; 
		'd7:S_7 <= i; 
		'd8:S_8 <= i; 
		'd9:S_9 <= i; 
		'd10:S_10 <= i; 
		'd11:S_11 <= i; 
		'd12:S_12 <= i; 
		'd13:S_13 <= i; 
		'd14:S_14 <= i; 
		'd15:S_15 <= i; 
		'd16:S_16 <= i; 
		'd17:S_17 <= i; 
		'd18:S_18 <= i; 
		'd19:S_19 <= i; 
		'd20:S_20 <= i; 
		'd21:S_21 <= i; 
		'd22:S_22 <= i; 
		'd23:S_23 <= i; 
		'd24:S_24 <= i; 
		'd25:S_25 <= i; 
		'd26:S_26 <= i; 
		'd27:S_27 <= i; 
		'd28:S_28 <= i; 
		'd29:S_29 <= i; 
		'd30:S_30 <= i; 
		'd31:S_31 <= i; 
		'd32:S_32 <= i; 
		'd33:S_33 <= i; 
		'd34:S_34 <= i; 
		'd35:S_35 <= i; 
		'd36:S_36 <= i; 
		'd37:S_37 <= i; 
		'd38:S_38 <= i; 
		'd39:S_39 <= i; 
		'd40:S_40 <= i; 
		'd41:S_41 <= i; 
		'd42:S_42 <= i; 
		'd43:S_43 <= i; 
		'd44:S_44 <= i; 
		'd45:S_45 <= i; 
		'd46:S_46 <= i; 
		'd47:S_47 <= i; 
		'd48:S_48 <= i; 
		'd49:S_49 <= i; 
		'd50:S_50 <= i; 
		'd51:S_51 <= i; 
		'd52:S_52 <= i; 
		'd53:S_53 <= i; 
		'd54:S_54 <= i; 
		'd55:S_55 <= i; 
		'd56:S_56 <= i; 
		'd57:S_57 <= i; 
		'd58:S_58 <= i; 
		'd59:S_59 <= i; 
		'd60:S_60 <= i; 
		'd61:S_61 <= i; 
		'd62:S_62 <= i; 
		'd63:S_63 <= i; 
		'd64:S_64 <= i; 
		'd65:S_65 <= i; 
		'd66:S_66 <= i; 
		'd67:S_67 <= i; 
		'd68:S_68 <= i; 
		'd69:S_69 <= i; 
		'd70:S_70 <= i; 
		'd71:S_71 <= i; 
		'd72:S_72 <= i; 
		'd73:S_73 <= i; 
		'd74:S_74 <= i; 
		'd75:S_75 <= i; 
		'd76:S_76 <= i; 
		'd77:S_77 <= i; 
		'd78:S_78 <= i; 
		'd79:S_79 <= i; 
		'd80:S_80 <= i; 
		'd81:S_81 <= i; 
		'd82:S_82 <= i; 
		'd83:S_83 <= i; 
		'd84:S_84 <= i; 
		'd85:S_85 <= i; 
		'd86:S_86 <= i; 
		'd87:S_87 <= i; 
		'd88:S_88 <= i; 
		'd89:S_89 <= i; 
		'd90:S_90 <= i; 
		'd91:S_91 <= i; 
		'd92:S_92 <= i; 
		'd93:S_93 <= i; 
		'd94:S_94 <= i; 
		'd95:S_95 <= i; 
		'd96:S_96 <= i; 
		'd97:S_97 <= i; 
		'd98:S_98 <= i; 
		'd99:S_99 <= i; 
		'd100:S_100 <= i; 
		'd101:S_101 <= i; 
		'd102:S_102 <= i; 
		'd103:S_103 <= i; 
		'd104:S_104 <= i; 
		'd105:S_105 <= i; 
		'd106:S_106 <= i; 
		'd107:S_107 <= i; 
		'd108:S_108 <= i; 
		'd109:S_109 <= i; 
		'd110:S_110 <= i; 
		'd111:S_111 <= i; 
		'd112:S_112 <= i; 
		'd113:S_113 <= i; 
		'd114:S_114 <= i; 
		'd115:S_115 <= i; 
		'd116:S_116 <= i; 
		'd117:S_117 <= i; 
		'd118:S_118 <= i; 
		'd119:S_119 <= i; 
		'd120:S_120 <= i; 
		'd121:S_121 <= i; 
		'd122:S_122 <= i; 
		'd123:S_123 <= i; 
		'd124:S_124 <= i; 
		'd125:S_125 <= i; 
		'd126:S_126 <= i; 
		'd127:S_127 <= i; 
		'd128:S_128 <= i; 
		'd129:S_129 <= i; 
		'd130:S_130 <= i; 
		'd131:S_131 <= i; 
		'd132:S_132 <= i; 
		'd133:S_133 <= i; 
		'd134:S_134 <= i; 
		'd135:S_135 <= i; 
		'd136:S_136 <= i; 
		'd137:S_137 <= i; 
		'd138:S_138 <= i; 
		'd139:S_139 <= i; 
		'd140:S_140 <= i; 
		'd141:S_141 <= i; 
		'd142:S_142 <= i; 
		'd143:S_143 <= i; 
		'd144:S_144 <= i; 
		'd145:S_145 <= i; 
		'd146:S_146 <= i; 
		'd147:S_147 <= i; 
		'd148:S_148 <= i; 
		'd149:S_149 <= i; 
		'd150:S_150 <= i; 
		'd151:S_151 <= i; 
		'd152:S_152 <= i; 
		'd153:S_153 <= i; 
		'd154:S_154 <= i; 
		'd155:S_155 <= i; 
		'd156:S_156 <= i; 
		'd157:S_157 <= i; 
		'd158:S_158 <= i; 
		'd159:S_159 <= i; 
		'd160:S_160 <= i; 
		'd161:S_161 <= i; 
		'd162:S_162 <= i; 
		'd163:S_163 <= i; 
		'd164:S_164 <= i; 
		'd165:S_165 <= i; 
		'd166:S_166 <= i; 
		'd167:S_167 <= i; 
		'd168:S_168 <= i; 
		'd169:S_169 <= i; 
		'd170:S_170 <= i; 
		'd171:S_171 <= i; 
		'd172:S_172 <= i; 
		'd173:S_173 <= i; 
		'd174:S_174 <= i; 
		'd175:S_175 <= i; 
		'd176:S_176 <= i; 
		'd177:S_177 <= i; 
		'd178:S_178 <= i; 
		'd179:S_179 <= i; 
		'd180:S_180 <= i; 
		'd181:S_181 <= i; 
		'd182:S_182 <= i; 
		'd183:S_183 <= i; 
		'd184:S_184 <= i; 
		'd185:S_185 <= i; 
		'd186:S_186 <= i; 
		'd187:S_187 <= i; 
		'd188:S_188 <= i; 
		'd189:S_189 <= i; 
		'd190:S_190 <= i; 
		'd191:S_191 <= i; 
		'd192:S_192 <= i; 
		'd193:S_193 <= i; 
		'd194:S_194 <= i; 
		'd195:S_195 <= i; 
		'd196:S_196 <= i; 
		'd197:S_197 <= i; 
		'd198:S_198 <= i; 
		'd199:S_199 <= i; 
		'd200:S_200 <= i; 
		'd201:S_201 <= i; 
		'd202:S_202 <= i; 
		'd203:S_203 <= i; 
		'd204:S_204 <= i; 
		'd205:S_205 <= i; 
		'd206:S_206 <= i; 
		'd207:S_207 <= i; 
		'd208:S_208 <= i; 
		'd209:S_209 <= i; 
		'd210:S_210 <= i; 
		'd211:S_211 <= i; 
		'd212:S_212 <= i; 
		'd213:S_213 <= i; 
		'd214:S_214 <= i; 
		'd215:S_215 <= i; 
		'd216:S_216 <= i; 
		'd217:S_217 <= i; 
		'd218:S_218 <= i; 
		'd219:S_219 <= i; 
		'd220:S_220 <= i; 
		'd221:S_221 <= i; 
		'd222:S_222 <= i; 
		'd223:S_223 <= i; 
		'd224:S_224 <= i; 
		'd225:S_225 <= i; 
		'd226:S_226 <= i; 
		'd227:S_227 <= i; 
		'd228:S_228 <= i; 
		'd229:S_229 <= i; 
		'd230:S_230 <= i; 
		'd231:S_231 <= i; 
		'd232:S_232 <= i; 
		'd233:S_233 <= i; 
		'd234:S_234 <= i; 
		'd235:S_235 <= i; 
		'd236:S_236 <= i; 
		'd237:S_237 <= i; 
		'd238:S_238 <= i; 
		'd239:S_239 <= i; 
		'd240:S_240 <= i; 
		'd241:S_241 <= i; 
		'd242:S_242 <= i; 
		'd243:S_243 <= i; 
		'd244:S_244 <= i; 
		'd245:S_245 <= i; 
		'd246:S_246 <= i; 
		'd247:S_247 <= i; 
		'd248:S_248 <= i; 
		'd249:S_249 <= i; 
		'd250:S_250 <= i; 
		'd251:S_251 <= i; 
		'd252:S_252 <= i; 
		'd253:S_253 <= i; 
		'd254:S_254 <= i; 
		'd255:S_255 <= i; 
		default:S_256 <= i; 
	endcase
				if (i == 8'hFF) begin
					KSState <= 4'h2;
					i <= 8'h00;
				end else begin
					i <= i +1;
				end
			end

	// j := 0
	// for i from 0 to 255
	//     j := (j + S[i] + key[i mod keylength]) mod 256
	//     swap values of S[i] and S[j]
	// endfor

			4'h2: begin // KSS_KEYSCHED2: Initialize S array
				// in place of:
				// j <= (j + S[i] + key[i % `KEY_SIZE]);
				j <= (j + S_of_i + key_of_i_mod_KEYSIZE);
				KSState <= 4'h3;
			end

			4'h3: begin // KSS_KEYSCHED3: S array permutation
				// in place of:
				// S[i]<=S[j]; , see KSS_SWAP_REGS*
				// in place of:
				// S[j]<=S[i];
				case (j) 
		'd0:S_0 <= S_of_i; 
		'd1:S_1 <= S_of_i; 
		'd2:S_2 <= S_of_i; 
		'd3:S_3 <= S_of_i; 
		'd4:S_4 <= S_of_i; 
		'd5:S_5 <= S_of_i; 
		'd6:S_6 <= S_of_i; 
		'd7:S_7 <= S_of_i; 
		'd8:S_8 <= S_of_i; 
		'd9:S_9 <= S_of_i; 
		'd10:S_10 <= S_of_i; 
		'd11:S_11 <= S_of_i; 
		'd12:S_12 <= S_of_i; 
		'd13:S_13 <= S_of_i; 
		'd14:S_14 <= S_of_i; 
		'd15:S_15 <= S_of_i; 
		'd16:S_16 <= S_of_i; 
		'd17:S_17 <= S_of_i; 
		'd18:S_18 <= S_of_i; 
		'd19:S_19 <= S_of_i; 
		'd20:S_20 <= S_of_i; 
		'd21:S_21 <= S_of_i; 
		'd22:S_22 <= S_of_i; 
		'd23:S_23 <= S_of_i; 
		'd24:S_24 <= S_of_i; 
		'd25:S_25 <= S_of_i; 
		'd26:S_26 <= S_of_i; 
		'd27:S_27 <= S_of_i; 
		'd28:S_28 <= S_of_i; 
		'd29:S_29 <= S_of_i; 
		'd30:S_30 <= S_of_i; 
		'd31:S_31 <= S_of_i; 
		'd32:S_32 <= S_of_i; 
		'd33:S_33 <= S_of_i; 
		'd34:S_34 <= S_of_i; 
		'd35:S_35 <= S_of_i; 
		'd36:S_36 <= S_of_i; 
		'd37:S_37 <= S_of_i; 
		'd38:S_38 <= S_of_i; 
		'd39:S_39 <= S_of_i; 
		'd40:S_40 <= S_of_i; 
		'd41:S_41 <= S_of_i; 
		'd42:S_42 <= S_of_i; 
		'd43:S_43 <= S_of_i; 
		'd44:S_44 <= S_of_i; 
		'd45:S_45 <= S_of_i; 
		'd46:S_46 <= S_of_i; 
		'd47:S_47 <= S_of_i; 
		'd48:S_48 <= S_of_i; 
		'd49:S_49 <= S_of_i; 
		'd50:S_50 <= S_of_i; 
		'd51:S_51 <= S_of_i; 
		'd52:S_52 <= S_of_i; 
		'd53:S_53 <= S_of_i; 
		'd54:S_54 <= S_of_i; 
		'd55:S_55 <= S_of_i; 
		'd56:S_56 <= S_of_i; 
		'd57:S_57 <= S_of_i; 
		'd58:S_58 <= S_of_i; 
		'd59:S_59 <= S_of_i; 
		'd60:S_60 <= S_of_i; 
		'd61:S_61 <= S_of_i; 
		'd62:S_62 <= S_of_i; 
		'd63:S_63 <= S_of_i; 
		'd64:S_64 <= S_of_i; 
		'd65:S_65 <= S_of_i; 
		'd66:S_66 <= S_of_i; 
		'd67:S_67 <= S_of_i; 
		'd68:S_68 <= S_of_i; 
		'd69:S_69 <= S_of_i; 
		'd70:S_70 <= S_of_i; 
		'd71:S_71 <= S_of_i; 
		'd72:S_72 <= S_of_i; 
		'd73:S_73 <= S_of_i; 
		'd74:S_74 <= S_of_i; 
		'd75:S_75 <= S_of_i; 
		'd76:S_76 <= S_of_i; 
		'd77:S_77 <= S_of_i; 
		'd78:S_78 <= S_of_i; 
		'd79:S_79 <= S_of_i; 
		'd80:S_80 <= S_of_i; 
		'd81:S_81 <= S_of_i; 
		'd82:S_82 <= S_of_i; 
		'd83:S_83 <= S_of_i; 
		'd84:S_84 <= S_of_i; 
		'd85:S_85 <= S_of_i; 
		'd86:S_86 <= S_of_i; 
		'd87:S_87 <= S_of_i; 
		'd88:S_88 <= S_of_i; 
		'd89:S_89 <= S_of_i; 
		'd90:S_90 <= S_of_i; 
		'd91:S_91 <= S_of_i; 
		'd92:S_92 <= S_of_i; 
		'd93:S_93 <= S_of_i; 
		'd94:S_94 <= S_of_i; 
		'd95:S_95 <= S_of_i; 
		'd96:S_96 <= S_of_i; 
		'd97:S_97 <= S_of_i; 
		'd98:S_98 <= S_of_i; 
		'd99:S_99 <= S_of_i; 
		'd100:S_100 <= S_of_i; 
		'd101:S_101 <= S_of_i; 
		'd102:S_102 <= S_of_i; 
		'd103:S_103 <= S_of_i; 
		'd104:S_104 <= S_of_i; 
		'd105:S_105 <= S_of_i; 
		'd106:S_106 <= S_of_i; 
		'd107:S_107 <= S_of_i; 
		'd108:S_108 <= S_of_i; 
		'd109:S_109 <= S_of_i; 
		'd110:S_110 <= S_of_i; 
		'd111:S_111 <= S_of_i; 
		'd112:S_112 <= S_of_i; 
		'd113:S_113 <= S_of_i; 
		'd114:S_114 <= S_of_i; 
		'd115:S_115 <= S_of_i; 
		'd116:S_116 <= S_of_i; 
		'd117:S_117 <= S_of_i; 
		'd118:S_118 <= S_of_i; 
		'd119:S_119 <= S_of_i; 
		'd120:S_120 <= S_of_i; 
		'd121:S_121 <= S_of_i; 
		'd122:S_122 <= S_of_i; 
		'd123:S_123 <= S_of_i; 
		'd124:S_124 <= S_of_i; 
		'd125:S_125 <= S_of_i; 
		'd126:S_126 <= S_of_i; 
		'd127:S_127 <= S_of_i; 
		'd128:S_128 <= S_of_i; 
		'd129:S_129 <= S_of_i; 
		'd130:S_130 <= S_of_i; 
		'd131:S_131 <= S_of_i; 
		'd132:S_132 <= S_of_i; 
		'd133:S_133 <= S_of_i; 
		'd134:S_134 <= S_of_i; 
		'd135:S_135 <= S_of_i; 
		'd136:S_136 <= S_of_i; 
		'd137:S_137 <= S_of_i; 
		'd138:S_138 <= S_of_i; 
		'd139:S_139 <= S_of_i; 
		'd140:S_140 <= S_of_i; 
		'd141:S_141 <= S_of_i; 
		'd142:S_142 <= S_of_i; 
		'd143:S_143 <= S_of_i; 
		'd144:S_144 <= S_of_i; 
		'd145:S_145 <= S_of_i; 
		'd146:S_146 <= S_of_i; 
		'd147:S_147 <= S_of_i; 
		'd148:S_148 <= S_of_i; 
		'd149:S_149 <= S_of_i; 
		'd150:S_150 <= S_of_i; 
		'd151:S_151 <= S_of_i; 
		'd152:S_152 <= S_of_i; 
		'd153:S_153 <= S_of_i; 
		'd154:S_154 <= S_of_i; 
		'd155:S_155 <= S_of_i; 
		'd156:S_156 <= S_of_i; 
		'd157:S_157 <= S_of_i; 
		'd158:S_158 <= S_of_i; 
		'd159:S_159 <= S_of_i; 
		'd160:S_160 <= S_of_i; 
		'd161:S_161 <= S_of_i; 
		'd162:S_162 <= S_of_i; 
		'd163:S_163 <= S_of_i; 
		'd164:S_164 <= S_of_i; 
		'd165:S_165 <= S_of_i; 
		'd166:S_166 <= S_of_i; 
		'd167:S_167 <= S_of_i; 
		'd168:S_168 <= S_of_i; 
		'd169:S_169 <= S_of_i; 
		'd170:S_170 <= S_of_i; 
		'd171:S_171 <= S_of_i; 
		'd172:S_172 <= S_of_i; 
		'd173:S_173 <= S_of_i; 
		'd174:S_174 <= S_of_i; 
		'd175:S_175 <= S_of_i; 
		'd176:S_176 <= S_of_i; 
		'd177:S_177 <= S_of_i; 
		'd178:S_178 <= S_of_i; 
		'd179:S_179 <= S_of_i; 
		'd180:S_180 <= S_of_i; 
		'd181:S_181 <= S_of_i; 
		'd182:S_182 <= S_of_i; 
		'd183:S_183 <= S_of_i; 
		'd184:S_184 <= S_of_i; 
		'd185:S_185 <= S_of_i; 
		'd186:S_186 <= S_of_i; 
		'd187:S_187 <= S_of_i; 
		'd188:S_188 <= S_of_i; 
		'd189:S_189 <= S_of_i; 
		'd190:S_190 <= S_of_i; 
		'd191:S_191 <= S_of_i; 
		'd192:S_192 <= S_of_i; 
		'd193:S_193 <= S_of_i; 
		'd194:S_194 <= S_of_i; 
		'd195:S_195 <= S_of_i; 
		'd196:S_196 <= S_of_i; 
		'd197:S_197 <= S_of_i; 
		'd198:S_198 <= S_of_i; 
		'd199:S_199 <= S_of_i; 
		'd200:S_200 <= S_of_i; 
		'd201:S_201 <= S_of_i; 
		'd202:S_202 <= S_of_i; 
		'd203:S_203 <= S_of_i; 
		'd204:S_204 <= S_of_i; 
		'd205:S_205 <= S_of_i; 
		'd206:S_206 <= S_of_i; 
		'd207:S_207 <= S_of_i; 
		'd208:S_208 <= S_of_i; 
		'd209:S_209 <= S_of_i; 
		'd210:S_210 <= S_of_i; 
		'd211:S_211 <= S_of_i; 
		'd212:S_212 <= S_of_i; 
		'd213:S_213 <= S_of_i; 
		'd214:S_214 <= S_of_i; 
		'd215:S_215 <= S_of_i; 
		'd216:S_216 <= S_of_i; 
		'd217:S_217 <= S_of_i; 
		'd218:S_218 <= S_of_i; 
		'd219:S_219 <= S_of_i; 
		'd220:S_220 <= S_of_i; 
		'd221:S_221 <= S_of_i; 
		'd222:S_222 <= S_of_i; 
		'd223:S_223 <= S_of_i; 
		'd224:S_224 <= S_of_i; 
		'd225:S_225 <= S_of_i; 
		'd226:S_226 <= S_of_i; 
		'd227:S_227 <= S_of_i; 
		'd228:S_228 <= S_of_i; 
		'd229:S_229 <= S_of_i; 
		'd230:S_230 <= S_of_i; 
		'd231:S_231 <= S_of_i; 
		'd232:S_232 <= S_of_i; 
		'd233:S_233 <= S_of_i; 
		'd234:S_234 <= S_of_i; 
		'd235:S_235 <= S_of_i; 
		'd236:S_236 <= S_of_i; 
		'd237:S_237 <= S_of_i; 
		'd238:S_238 <= S_of_i; 
		'd239:S_239 <= S_of_i; 
		'd240:S_240 <= S_of_i; 
		'd241:S_241 <= S_of_i; 
		'd242:S_242 <= S_of_i; 
		'd243:S_243 <= S_of_i; 
		'd244:S_244 <= S_of_i; 
		'd245:S_245 <= S_of_i; 
		'd246:S_246 <= S_of_i; 
		'd247:S_247 <= S_of_i; 
		'd248:S_248 <= S_of_i; 
		'd249:S_249 <= S_of_i; 
		'd250:S_250 <= S_of_i; 
		'd251:S_251 <= S_of_i; 
		'd252:S_252 <= S_of_i; 
		'd253:S_253 <= S_of_i; 
		'd254:S_254 <= S_of_i; 
		'd255:S_255 <= S_of_i; 
		default:S_256 <= S_of_i; 
	endcase
				if (i == 8'hFF) begin
					KSState <= 4'h7;
					i <= 8'h01;
					j <= S_1;
					discardCount <= 11'h0;
					output_ready <= 0; // K not valid yet
				end else begin
					i <= i + 1;
					KSState <= 4'h5;
				end
			end

	// i := 0
	// j := 0
	// while GeneratingOutput:
	//     i := (i + 1) mod 256
	//     j := (j + S[i]) mod 256
	//     swap values of S[i] and S[j]
	//     K := S[(S[i] + S[j]) mod 256]
	//     output K
	// endwhile

			4'h4: begin
				// in place of:
				// S[i] <= S[j], see KSS_SWAP_REGS*
				// in place of:
				// S[j] <= S[i]; // We can do this because of verilog.
				case (j) 
		'd0:S_0 <= S_of_i; 
		'd1:S_1 <= S_of_i; 
		'd2:S_2 <= S_of_i; 
		'd3:S_3 <= S_of_i; 
		'd4:S_4 <= S_of_i; 
		'd5:S_5 <= S_of_i; 
		'd6:S_6 <= S_of_i; 
		'd7:S_7 <= S_of_i; 
		'd8:S_8 <= S_of_i; 
		'd9:S_9 <= S_of_i; 
		'd10:S_10 <= S_of_i; 
		'd11:S_11 <= S_of_i; 
		'd12:S_12 <= S_of_i; 
		'd13:S_13 <= S_of_i; 
		'd14:S_14 <= S_of_i; 
		'd15:S_15 <= S_of_i; 
		'd16:S_16 <= S_of_i; 
		'd17:S_17 <= S_of_i; 
		'd18:S_18 <= S_of_i; 
		'd19:S_19 <= S_of_i; 
		'd20:S_20 <= S_of_i; 
		'd21:S_21 <= S_of_i; 
		'd22:S_22 <= S_of_i; 
		'd23:S_23 <= S_of_i; 
		'd24:S_24 <= S_of_i; 
		'd25:S_25 <= S_of_i; 
		'd26:S_26 <= S_of_i; 
		'd27:S_27 <= S_of_i; 
		'd28:S_28 <= S_of_i; 
		'd29:S_29 <= S_of_i; 
		'd30:S_30 <= S_of_i; 
		'd31:S_31 <= S_of_i; 
		'd32:S_32 <= S_of_i; 
		'd33:S_33 <= S_of_i; 
		'd34:S_34 <= S_of_i; 
		'd35:S_35 <= S_of_i; 
		'd36:S_36 <= S_of_i; 
		'd37:S_37 <= S_of_i; 
		'd38:S_38 <= S_of_i; 
		'd39:S_39 <= S_of_i; 
		'd40:S_40 <= S_of_i; 
		'd41:S_41 <= S_of_i; 
		'd42:S_42 <= S_of_i; 
		'd43:S_43 <= S_of_i; 
		'd44:S_44 <= S_of_i; 
		'd45:S_45 <= S_of_i; 
		'd46:S_46 <= S_of_i; 
		'd47:S_47 <= S_of_i; 
		'd48:S_48 <= S_of_i; 
		'd49:S_49 <= S_of_i; 
		'd50:S_50 <= S_of_i; 
		'd51:S_51 <= S_of_i; 
		'd52:S_52 <= S_of_i; 
		'd53:S_53 <= S_of_i; 
		'd54:S_54 <= S_of_i; 
		'd55:S_55 <= S_of_i; 
		'd56:S_56 <= S_of_i; 
		'd57:S_57 <= S_of_i; 
		'd58:S_58 <= S_of_i; 
		'd59:S_59 <= S_of_i; 
		'd60:S_60 <= S_of_i; 
		'd61:S_61 <= S_of_i; 
		'd62:S_62 <= S_of_i; 
		'd63:S_63 <= S_of_i; 
		'd64:S_64 <= S_of_i; 
		'd65:S_65 <= S_of_i; 
		'd66:S_66 <= S_of_i; 
		'd67:S_67 <= S_of_i; 
		'd68:S_68 <= S_of_i; 
		'd69:S_69 <= S_of_i; 
		'd70:S_70 <= S_of_i; 
		'd71:S_71 <= S_of_i; 
		'd72:S_72 <= S_of_i; 
		'd73:S_73 <= S_of_i; 
		'd74:S_74 <= S_of_i; 
		'd75:S_75 <= S_of_i; 
		'd76:S_76 <= S_of_i; 
		'd77:S_77 <= S_of_i; 
		'd78:S_78 <= S_of_i; 
		'd79:S_79 <= S_of_i; 
		'd80:S_80 <= S_of_i; 
		'd81:S_81 <= S_of_i; 
		'd82:S_82 <= S_of_i; 
		'd83:S_83 <= S_of_i; 
		'd84:S_84 <= S_of_i; 
		'd85:S_85 <= S_of_i; 
		'd86:S_86 <= S_of_i; 
		'd87:S_87 <= S_of_i; 
		'd88:S_88 <= S_of_i; 
		'd89:S_89 <= S_of_i; 
		'd90:S_90 <= S_of_i; 
		'd91:S_91 <= S_of_i; 
		'd92:S_92 <= S_of_i; 
		'd93:S_93 <= S_of_i; 
		'd94:S_94 <= S_of_i; 
		'd95:S_95 <= S_of_i; 
		'd96:S_96 <= S_of_i; 
		'd97:S_97 <= S_of_i; 
		'd98:S_98 <= S_of_i; 
		'd99:S_99 <= S_of_i; 
		'd100:S_100 <= S_of_i; 
		'd101:S_101 <= S_of_i; 
		'd102:S_102 <= S_of_i; 
		'd103:S_103 <= S_of_i; 
		'd104:S_104 <= S_of_i; 
		'd105:S_105 <= S_of_i; 
		'd106:S_106 <= S_of_i; 
		'd107:S_107 <= S_of_i; 
		'd108:S_108 <= S_of_i; 
		'd109:S_109 <= S_of_i; 
		'd110:S_110 <= S_of_i; 
		'd111:S_111 <= S_of_i; 
		'd112:S_112 <= S_of_i; 
		'd113:S_113 <= S_of_i; 
		'd114:S_114 <= S_of_i; 
		'd115:S_115 <= S_of_i; 
		'd116:S_116 <= S_of_i; 
		'd117:S_117 <= S_of_i; 
		'd118:S_118 <= S_of_i; 
		'd119:S_119 <= S_of_i; 
		'd120:S_120 <= S_of_i; 
		'd121:S_121 <= S_of_i; 
		'd122:S_122 <= S_of_i; 
		'd123:S_123 <= S_of_i; 
		'd124:S_124 <= S_of_i; 
		'd125:S_125 <= S_of_i; 
		'd126:S_126 <= S_of_i; 
		'd127:S_127 <= S_of_i; 
		'd128:S_128 <= S_of_i; 
		'd129:S_129 <= S_of_i; 
		'd130:S_130 <= S_of_i; 
		'd131:S_131 <= S_of_i; 
		'd132:S_132 <= S_of_i; 
		'd133:S_133 <= S_of_i; 
		'd134:S_134 <= S_of_i; 
		'd135:S_135 <= S_of_i; 
		'd136:S_136 <= S_of_i; 
		'd137:S_137 <= S_of_i; 
		'd138:S_138 <= S_of_i; 
		'd139:S_139 <= S_of_i; 
		'd140:S_140 <= S_of_i; 
		'd141:S_141 <= S_of_i; 
		'd142:S_142 <= S_of_i; 
		'd143:S_143 <= S_of_i; 
		'd144:S_144 <= S_of_i; 
		'd145:S_145 <= S_of_i; 
		'd146:S_146 <= S_of_i; 
		'd147:S_147 <= S_of_i; 
		'd148:S_148 <= S_of_i; 
		'd149:S_149 <= S_of_i; 
		'd150:S_150 <= S_of_i; 
		'd151:S_151 <= S_of_i; 
		'd152:S_152 <= S_of_i; 
		'd153:S_153 <= S_of_i; 
		'd154:S_154 <= S_of_i; 
		'd155:S_155 <= S_of_i; 
		'd156:S_156 <= S_of_i; 
		'd157:S_157 <= S_of_i; 
		'd158:S_158 <= S_of_i; 
		'd159:S_159 <= S_of_i; 
		'd160:S_160 <= S_of_i; 
		'd161:S_161 <= S_of_i; 
		'd162:S_162 <= S_of_i; 
		'd163:S_163 <= S_of_i; 
		'd164:S_164 <= S_of_i; 
		'd165:S_165 <= S_of_i; 
		'd166:S_166 <= S_of_i; 
		'd167:S_167 <= S_of_i; 
		'd168:S_168 <= S_of_i; 
		'd169:S_169 <= S_of_i; 
		'd170:S_170 <= S_of_i; 
		'd171:S_171 <= S_of_i; 
		'd172:S_172 <= S_of_i; 
		'd173:S_173 <= S_of_i; 
		'd174:S_174 <= S_of_i; 
		'd175:S_175 <= S_of_i; 
		'd176:S_176 <= S_of_i; 
		'd177:S_177 <= S_of_i; 
		'd178:S_178 <= S_of_i; 
		'd179:S_179 <= S_of_i; 
		'd180:S_180 <= S_of_i; 
		'd181:S_181 <= S_of_i; 
		'd182:S_182 <= S_of_i; 
		'd183:S_183 <= S_of_i; 
		'd184:S_184 <= S_of_i; 
		'd185:S_185 <= S_of_i; 
		'd186:S_186 <= S_of_i; 
		'd187:S_187 <= S_of_i; 
		'd188:S_188 <= S_of_i; 
		'd189:S_189 <= S_of_i; 
		'd190:S_190 <= S_of_i; 
		'd191:S_191 <= S_of_i; 
		'd192:S_192 <= S_of_i; 
		'd193:S_193 <= S_of_i; 
		'd194:S_194 <= S_of_i; 
		'd195:S_195 <= S_of_i; 
		'd196:S_196 <= S_of_i; 
		'd197:S_197 <= S_of_i; 
		'd198:S_198 <= S_of_i; 
		'd199:S_199 <= S_of_i; 
		'd200:S_200 <= S_of_i; 
		'd201:S_201 <= S_of_i; 
		'd202:S_202 <= S_of_i; 
		'd203:S_203 <= S_of_i; 
		'd204:S_204 <= S_of_i; 
		'd205:S_205 <= S_of_i; 
		'd206:S_206 <= S_of_i; 
		'd207:S_207 <= S_of_i; 
		'd208:S_208 <= S_of_i; 
		'd209:S_209 <= S_of_i; 
		'd210:S_210 <= S_of_i; 
		'd211:S_211 <= S_of_i; 
		'd212:S_212 <= S_of_i; 
		'd213:S_213 <= S_of_i; 
		'd214:S_214 <= S_of_i; 
		'd215:S_215 <= S_of_i; 
		'd216:S_216 <= S_of_i; 
		'd217:S_217 <= S_of_i; 
		'd218:S_218 <= S_of_i; 
		'd219:S_219 <= S_of_i; 
		'd220:S_220 <= S_of_i; 
		'd221:S_221 <= S_of_i; 
		'd222:S_222 <= S_of_i; 
		'd223:S_223 <= S_of_i; 
		'd224:S_224 <= S_of_i; 
		'd225:S_225 <= S_of_i; 
		'd226:S_226 <= S_of_i; 
		'd227:S_227 <= S_of_i; 
		'd228:S_228 <= S_of_i; 
		'd229:S_229 <= S_of_i; 
		'd230:S_230 <= S_of_i; 
		'd231:S_231 <= S_of_i; 
		'd232:S_232 <= S_of_i; 
		'd233:S_233 <= S_of_i; 
		'd234:S_234 <= S_of_i; 
		'd235:S_235 <= S_of_i; 
		'd236:S_236 <= S_of_i; 
		'd237:S_237 <= S_of_i; 
		'd238:S_238 <= S_of_i; 
		'd239:S_239 <= S_of_i; 
		'd240:S_240 <= S_of_i; 
		'd241:S_241 <= S_of_i; 
		'd242:S_242 <= S_of_i; 
		'd243:S_243 <= S_of_i; 
		'd244:S_244 <= S_of_i; 
		'd245:S_245 <= S_of_i; 
		'd246:S_246 <= S_of_i; 
		'd247:S_247 <= S_of_i; 
		'd248:S_248 <= S_of_i; 
		'd249:S_249 <= S_of_i; 
		'd250:S_250 <= S_of_i; 
		'd251:S_251 <= S_of_i; 
		'd252:S_252 <= S_of_i; 
		'd253:S_253 <= S_of_i; 
		'd254:S_254 <= S_of_i; 
		'd255:S_255 <= S_of_i; 
		default:S_256 <= S_of_i; 
	endcase
				// in place of:
				// K <= S[ S[i]+S[j] ];
				case (S_of_i_plus_S_of_j) 
		'd0:K <= S_0; 
		'd1:K <= S_1; 
		'd2:K <= S_2; 
		'd3:K <= S_3; 
		'd4:K <= S_4; 
		'd5:K <= S_5; 
		'd6:K <= S_6; 
		'd7:K <= S_7; 
		'd8:K <= S_8; 
		'd9:K <= S_9; 
		'd10:K <= S_10; 
		'd11:K <= S_11; 
		'd12:K <= S_12; 
		'd13:K <= S_13; 
		'd14:K <= S_14; 
		'd15:K <= S_15; 
		'd16:K <= S_16; 
		'd17:K <= S_17; 
		'd18:K <= S_18; 
		'd19:K <= S_19; 
		'd20:K <= S_20; 
		'd21:K <= S_21; 
		'd22:K <= S_22; 
		'd23:K <= S_23; 
		'd24:K <= S_24; 
		'd25:K <= S_25; 
		'd26:K <= S_26; 
		'd27:K <= S_27; 
		'd28:K <= S_28; 
		'd29:K <= S_29; 
		'd30:K <= S_30; 
		'd31:K <= S_31; 
		'd32:K <= S_32; 
		'd33:K <= S_33; 
		'd34:K <= S_34; 
		'd35:K <= S_35; 
		'd36:K <= S_36; 
		'd37:K <= S_37; 
		'd38:K <= S_38; 
		'd39:K <= S_39; 
		'd40:K <= S_40; 
		'd41:K <= S_41; 
		'd42:K <= S_42; 
		'd43:K <= S_43; 
		'd44:K <= S_44; 
		'd45:K <= S_45; 
		'd46:K <= S_46; 
		'd47:K <= S_47; 
		'd48:K <= S_48; 
		'd49:K <= S_49; 
		'd50:K <= S_50; 
		'd51:K <= S_51; 
		'd52:K <= S_52; 
		'd53:K <= S_53; 
		'd54:K <= S_54; 
		'd55:K <= S_55; 
		'd56:K <= S_56; 
		'd57:K <= S_57; 
		'd58:K <= S_58; 
		'd59:K <= S_59; 
		'd60:K <= S_60; 
		'd61:K <= S_61; 
		'd62:K <= S_62; 
		'd63:K <= S_63; 
		'd64:K <= S_64; 
		'd65:K <= S_65; 
		'd66:K <= S_66; 
		'd67:K <= S_67; 
		'd68:K <= S_68; 
		'd69:K <= S_69; 
		'd70:K <= S_70; 
		'd71:K <= S_71; 
		'd72:K <= S_72; 
		'd73:K <= S_73; 
		'd74:K <= S_74; 
		'd75:K <= S_75; 
		'd76:K <= S_76; 
		'd77:K <= S_77; 
		'd78:K <= S_78; 
		'd79:K <= S_79; 
		'd80:K <= S_80; 
		'd81:K <= S_81; 
		'd82:K <= S_82; 
		'd83:K <= S_83; 
		'd84:K <= S_84; 
		'd85:K <= S_85; 
		'd86:K <= S_86; 
		'd87:K <= S_87; 
		'd88:K <= S_88; 
		'd89:K <= S_89; 
		'd90:K <= S_90; 
		'd91:K <= S_91; 
		'd92:K <= S_92; 
		'd93:K <= S_93; 
		'd94:K <= S_94; 
		'd95:K <= S_95; 
		'd96:K <= S_96; 
		'd97:K <= S_97; 
		'd98:K <= S_98; 
		'd99:K <= S_99; 
		'd100:K <= S_100; 
		'd101:K <= S_101; 
		'd102:K <= S_102; 
		'd103:K <= S_103; 
		'd104:K <= S_104; 
		'd105:K <= S_105; 
		'd106:K <= S_106; 
		'd107:K <= S_107; 
		'd108:K <= S_108; 
		'd109:K <= S_109; 
		'd110:K <= S_110; 
		'd111:K <= S_111; 
		'd112:K <= S_112; 
		'd113:K <= S_113; 
		'd114:K <= S_114; 
		'd115:K <= S_115; 
		'd116:K <= S_116; 
		'd117:K <= S_117; 
		'd118:K <= S_118; 
		'd119:K <= S_119; 
		'd120:K <= S_120; 
		'd121:K <= S_121; 
		'd122:K <= S_122; 
		'd123:K <= S_123; 
		'd124:K <= S_124; 
		'd125:K <= S_125; 
		'd126:K <= S_126; 
		'd127:K <= S_127; 
		'd128:K <= S_128; 
		'd129:K <= S_129; 
		'd130:K <= S_130; 
		'd131:K <= S_131; 
		'd132:K <= S_132; 
		'd133:K <= S_133; 
		'd134:K <= S_134; 
		'd135:K <= S_135; 
		'd136:K <= S_136; 
		'd137:K <= S_137; 
		'd138:K <= S_138; 
		'd139:K <= S_139; 
		'd140:K <= S_140; 
		'd141:K <= S_141; 
		'd142:K <= S_142; 
		'd143:K <= S_143; 
		'd144:K <= S_144; 
		'd145:K <= S_145; 
		'd146:K <= S_146; 
		'd147:K <= S_147; 
		'd148:K <= S_148; 
		'd149:K <= S_149; 
		'd150:K <= S_150; 
		'd151:K <= S_151; 
		'd152:K <= S_152; 
		'd153:K <= S_153; 
		'd154:K <= S_154; 
		'd155:K <= S_155; 
		'd156:K <= S_156; 
		'd157:K <= S_157; 
		'd158:K <= S_158; 
		'd159:K <= S_159; 
		'd160:K <= S_160; 
		'd161:K <= S_161; 
		'd162:K <= S_162; 
		'd163:K <= S_163; 
		'd164:K <= S_164; 
		'd165:K <= S_165; 
		'd166:K <= S_166; 
		'd167:K <= S_167; 
		'd168:K <= S_168; 
		'd169:K <= S_169; 
		'd170:K <= S_170; 
		'd171:K <= S_171; 
		'd172:K <= S_172; 
		'd173:K <= S_173; 
		'd174:K <= S_174; 
		'd175:K <= S_175; 
		'd176:K <= S_176; 
		'd177:K <= S_177; 
		'd178:K <= S_178; 
		'd179:K <= S_179; 
		'd180:K <= S_180; 
		'd181:K <= S_181; 
		'd182:K <= S_182; 
		'd183:K <= S_183; 
		'd184:K <= S_184; 
		'd185:K <= S_185; 
		'd186:K <= S_186; 
		'd187:K <= S_187; 
		'd188:K <= S_188; 
		'd189:K <= S_189; 
		'd190:K <= S_190; 
		'd191:K <= S_191; 
		'd192:K <= S_192; 
		'd193:K <= S_193; 
		'd194:K <= S_194; 
		'd195:K <= S_195; 
		'd196:K <= S_196; 
		'd197:K <= S_197; 
		'd198:K <= S_198; 
		'd199:K <= S_199; 
		'd200:K <= S_200; 
		'd201:K <= S_201; 
		'd202:K <= S_202; 
		'd203:K <= S_203; 
		'd204:K <= S_204; 
		'd205:K <= S_205; 
		'd206:K <= S_206; 
		'd207:K <= S_207; 
		'd208:K <= S_208; 
		'd209:K <= S_209; 
		'd210:K <= S_210; 
		'd211:K <= S_211; 
		'd212:K <= S_212; 
		'd213:K <= S_213; 
		'd214:K <= S_214; 
		'd215:K <= S_215; 
		'd216:K <= S_216; 
		'd217:K <= S_217; 
		'd218:K <= S_218; 
		'd219:K <= S_219; 
		'd220:K <= S_220; 
		'd221:K <= S_221; 
		'd222:K <= S_222; 
		'd223:K <= S_223; 
		'd224:K <= S_224; 
		'd225:K <= S_225; 
		'd226:K <= S_226; 
		'd227:K <= S_227; 
		'd228:K <= S_228; 
		'd229:K <= S_229; 
		'd230:K <= S_230; 
		'd231:K <= S_231; 
		'd232:K <= S_232; 
		'd233:K <= S_233; 
		'd234:K <= S_234; 
		'd235:K <= S_235; 
		'd236:K <= S_236; 
		'd237:K <= S_237; 
		'd238:K <= S_238; 
		'd239:K <= S_239; 
		'd240:K <= S_240; 
		'd241:K <= S_241; 
		'd242:K <= S_242; 
		'd243:K <= S_243; 
		'd244:K <= S_244; 
		'd245:K <= S_245; 
		'd246:K <= S_246; 
		'd247:K <= S_247; 
		'd248:K <= S_248; 
		'd249:K <= S_249; 
		'd250:K <= S_250; 
		'd251:K <= S_251; 
		'd252:K <= S_252; 
		'd253:K <= S_253; 
		'd254:K <= S_254; 
		'd255:K <= S_255; 
		default:K <= S_256; 
	endcase
				if (discardCount<11'h600) begin // discard first 1536 values / RFC 4345
					discardCount<=discardCount+1;
				end else begin
					output_ready <= 1; // Valid K at output
				end

				i <= i+1;
				// Here is the secret of 1-clock: we develop all possible values of j in the future
				if (j==i+1) begin
				     // j <= (j + S[i]);
				     j <= (j + S_of_i);
				end else begin
					if (i==255) begin
						j <= (j + S_0);
					end else begin
						// in place of:
						// j <= (j + S[i+1]);
						j <= (j + S_of_i_plus_1);
					end
				end
				//$display ("rc4: output = %08X",K);
			end

			default: begin
				case (prev_i) 
		'd0:S_0 <= prev_S_of_j; 
		'd1:S_1 <= prev_S_of_j; 
		'd2:S_2 <= prev_S_of_j; 
		'd3:S_3 <= prev_S_of_j; 
		'd4:S_4 <= prev_S_of_j; 
		'd5:S_5 <= prev_S_of_j; 
		'd6:S_6 <= prev_S_of_j; 
		'd7:S_7 <= prev_S_of_j; 
		'd8:S_8 <= prev_S_of_j; 
		'd9:S_9 <= prev_S_of_j; 
		'd10:S_10 <= prev_S_of_j; 
		'd11:S_11 <= prev_S_of_j; 
		'd12:S_12 <= prev_S_of_j; 
		'd13:S_13 <= prev_S_of_j; 
		'd14:S_14 <= prev_S_of_j; 
		'd15:S_15 <= prev_S_of_j; 
		'd16:S_16 <= prev_S_of_j; 
		'd17:S_17 <= prev_S_of_j; 
		'd18:S_18 <= prev_S_of_j; 
		'd19:S_19 <= prev_S_of_j; 
		'd20:S_20 <= prev_S_of_j; 
		'd21:S_21 <= prev_S_of_j; 
		'd22:S_22 <= prev_S_of_j; 
		'd23:S_23 <= prev_S_of_j; 
		'd24:S_24 <= prev_S_of_j; 
		'd25:S_25 <= prev_S_of_j; 
		'd26:S_26 <= prev_S_of_j; 
		'd27:S_27 <= prev_S_of_j; 
		'd28:S_28 <= prev_S_of_j; 
		'd29:S_29 <= prev_S_of_j; 
		'd30:S_30 <= prev_S_of_j; 
		'd31:S_31 <= prev_S_of_j; 
		'd32:S_32 <= prev_S_of_j; 
		'd33:S_33 <= prev_S_of_j; 
		'd34:S_34 <= prev_S_of_j; 
		'd35:S_35 <= prev_S_of_j; 
		'd36:S_36 <= prev_S_of_j; 
		'd37:S_37 <= prev_S_of_j; 
		'd38:S_38 <= prev_S_of_j; 
		'd39:S_39 <= prev_S_of_j; 
		'd40:S_40 <= prev_S_of_j; 
		'd41:S_41 <= prev_S_of_j; 
		'd42:S_42 <= prev_S_of_j; 
		'd43:S_43 <= prev_S_of_j; 
		'd44:S_44 <= prev_S_of_j; 
		'd45:S_45 <= prev_S_of_j; 
		'd46:S_46 <= prev_S_of_j; 
		'd47:S_47 <= prev_S_of_j; 
		'd48:S_48 <= prev_S_of_j; 
		'd49:S_49 <= prev_S_of_j; 
		'd50:S_50 <= prev_S_of_j; 
		'd51:S_51 <= prev_S_of_j; 
		'd52:S_52 <= prev_S_of_j; 
		'd53:S_53 <= prev_S_of_j; 
		'd54:S_54 <= prev_S_of_j; 
		'd55:S_55 <= prev_S_of_j; 
		'd56:S_56 <= prev_S_of_j; 
		'd57:S_57 <= prev_S_of_j; 
		'd58:S_58 <= prev_S_of_j; 
		'd59:S_59 <= prev_S_of_j; 
		'd60:S_60 <= prev_S_of_j; 
		'd61:S_61 <= prev_S_of_j; 
		'd62:S_62 <= prev_S_of_j; 
		'd63:S_63 <= prev_S_of_j; 
		'd64:S_64 <= prev_S_of_j; 
		'd65:S_65 <= prev_S_of_j; 
		'd66:S_66 <= prev_S_of_j; 
		'd67:S_67 <= prev_S_of_j; 
		'd68:S_68 <= prev_S_of_j; 
		'd69:S_69 <= prev_S_of_j; 
		'd70:S_70 <= prev_S_of_j; 
		'd71:S_71 <= prev_S_of_j; 
		'd72:S_72 <= prev_S_of_j; 
		'd73:S_73 <= prev_S_of_j; 
		'd74:S_74 <= prev_S_of_j; 
		'd75:S_75 <= prev_S_of_j; 
		'd76:S_76 <= prev_S_of_j; 
		'd77:S_77 <= prev_S_of_j; 
		'd78:S_78 <= prev_S_of_j; 
		'd79:S_79 <= prev_S_of_j; 
		'd80:S_80 <= prev_S_of_j; 
		'd81:S_81 <= prev_S_of_j; 
		'd82:S_82 <= prev_S_of_j; 
		'd83:S_83 <= prev_S_of_j; 
		'd84:S_84 <= prev_S_of_j; 
		'd85:S_85 <= prev_S_of_j; 
		'd86:S_86 <= prev_S_of_j; 
		'd87:S_87 <= prev_S_of_j; 
		'd88:S_88 <= prev_S_of_j; 
		'd89:S_89 <= prev_S_of_j; 
		'd90:S_90 <= prev_S_of_j; 
		'd91:S_91 <= prev_S_of_j; 
		'd92:S_92 <= prev_S_of_j; 
		'd93:S_93 <= prev_S_of_j; 
		'd94:S_94 <= prev_S_of_j; 
		'd95:S_95 <= prev_S_of_j; 
		'd96:S_96 <= prev_S_of_j; 
		'd97:S_97 <= prev_S_of_j; 
		'd98:S_98 <= prev_S_of_j; 
		'd99:S_99 <= prev_S_of_j; 
		'd100:S_100 <= prev_S_of_j; 
		'd101:S_101 <= prev_S_of_j; 
		'd102:S_102 <= prev_S_of_j; 
		'd103:S_103 <= prev_S_of_j; 
		'd104:S_104 <= prev_S_of_j; 
		'd105:S_105 <= prev_S_of_j; 
		'd106:S_106 <= prev_S_of_j; 
		'd107:S_107 <= prev_S_of_j; 
		'd108:S_108 <= prev_S_of_j; 
		'd109:S_109 <= prev_S_of_j; 
		'd110:S_110 <= prev_S_of_j; 
		'd111:S_111 <= prev_S_of_j; 
		'd112:S_112 <= prev_S_of_j; 
		'd113:S_113 <= prev_S_of_j; 
		'd114:S_114 <= prev_S_of_j; 
		'd115:S_115 <= prev_S_of_j; 
		'd116:S_116 <= prev_S_of_j; 
		'd117:S_117 <= prev_S_of_j; 
		'd118:S_118 <= prev_S_of_j; 
		'd119:S_119 <= prev_S_of_j; 
		'd120:S_120 <= prev_S_of_j; 
		'd121:S_121 <= prev_S_of_j; 
		'd122:S_122 <= prev_S_of_j; 
		'd123:S_123 <= prev_S_of_j; 
		'd124:S_124 <= prev_S_of_j; 
		'd125:S_125 <= prev_S_of_j; 
		'd126:S_126 <= prev_S_of_j; 
		'd127:S_127 <= prev_S_of_j; 
		'd128:S_128 <= prev_S_of_j; 
		'd129:S_129 <= prev_S_of_j; 
		'd130:S_130 <= prev_S_of_j; 
		'd131:S_131 <= prev_S_of_j; 
		'd132:S_132 <= prev_S_of_j; 
		'd133:S_133 <= prev_S_of_j; 
		'd134:S_134 <= prev_S_of_j; 
		'd135:S_135 <= prev_S_of_j; 
		'd136:S_136 <= prev_S_of_j; 
		'd137:S_137 <= prev_S_of_j; 
		'd138:S_138 <= prev_S_of_j; 
		'd139:S_139 <= prev_S_of_j; 
		'd140:S_140 <= prev_S_of_j; 
		'd141:S_141 <= prev_S_of_j; 
		'd142:S_142 <= prev_S_of_j; 
		'd143:S_143 <= prev_S_of_j; 
		'd144:S_144 <= prev_S_of_j; 
		'd145:S_145 <= prev_S_of_j; 
		'd146:S_146 <= prev_S_of_j; 
		'd147:S_147 <= prev_S_of_j; 
		'd148:S_148 <= prev_S_of_j; 
		'd149:S_149 <= prev_S_of_j; 
		'd150:S_150 <= prev_S_of_j; 
		'd151:S_151 <= prev_S_of_j; 
		'd152:S_152 <= prev_S_of_j; 
		'd153:S_153 <= prev_S_of_j; 
		'd154:S_154 <= prev_S_of_j; 
		'd155:S_155 <= prev_S_of_j; 
		'd156:S_156 <= prev_S_of_j; 
		'd157:S_157 <= prev_S_of_j; 
		'd158:S_158 <= prev_S_of_j; 
		'd159:S_159 <= prev_S_of_j; 
		'd160:S_160 <= prev_S_of_j; 
		'd161:S_161 <= prev_S_of_j; 
		'd162:S_162 <= prev_S_of_j; 
		'd163:S_163 <= prev_S_of_j; 
		'd164:S_164 <= prev_S_of_j; 
		'd165:S_165 <= prev_S_of_j; 
		'd166:S_166 <= prev_S_of_j; 
		'd167:S_167 <= prev_S_of_j; 
		'd168:S_168 <= prev_S_of_j; 
		'd169:S_169 <= prev_S_of_j; 
		'd170:S_170 <= prev_S_of_j; 
		'd171:S_171 <= prev_S_of_j; 
		'd172:S_172 <= prev_S_of_j; 
		'd173:S_173 <= prev_S_of_j; 
		'd174:S_174 <= prev_S_of_j; 
		'd175:S_175 <= prev_S_of_j; 
		'd176:S_176 <= prev_S_of_j; 
		'd177:S_177 <= prev_S_of_j; 
		'd178:S_178 <= prev_S_of_j; 
		'd179:S_179 <= prev_S_of_j; 
		'd180:S_180 <= prev_S_of_j; 
		'd181:S_181 <= prev_S_of_j; 
		'd182:S_182 <= prev_S_of_j; 
		'd183:S_183 <= prev_S_of_j; 
		'd184:S_184 <= prev_S_of_j; 
		'd185:S_185 <= prev_S_of_j; 
		'd186:S_186 <= prev_S_of_j; 
		'd187:S_187 <= prev_S_of_j; 
		'd188:S_188 <= prev_S_of_j; 
		'd189:S_189 <= prev_S_of_j; 
		'd190:S_190 <= prev_S_of_j; 
		'd191:S_191 <= prev_S_of_j; 
		'd192:S_192 <= prev_S_of_j; 
		'd193:S_193 <= prev_S_of_j; 
		'd194:S_194 <= prev_S_of_j; 
		'd195:S_195 <= prev_S_of_j; 
		'd196:S_196 <= prev_S_of_j; 
		'd197:S_197 <= prev_S_of_j; 
		'd198:S_198 <= prev_S_of_j; 
		'd199:S_199 <= prev_S_of_j; 
		'd200:S_200 <= prev_S_of_j; 
		'd201:S_201 <= prev_S_of_j; 
		'd202:S_202 <= prev_S_of_j; 
		'd203:S_203 <= prev_S_of_j; 
		'd204:S_204 <= prev_S_of_j; 
		'd205:S_205 <= prev_S_of_j; 
		'd206:S_206 <= prev_S_of_j; 
		'd207:S_207 <= prev_S_of_j; 
		'd208:S_208 <= prev_S_of_j; 
		'd209:S_209 <= prev_S_of_j; 
		'd210:S_210 <= prev_S_of_j; 
		'd211:S_211 <= prev_S_of_j; 
		'd212:S_212 <= prev_S_of_j; 
		'd213:S_213 <= prev_S_of_j; 
		'd214:S_214 <= prev_S_of_j; 
		'd215:S_215 <= prev_S_of_j; 
		'd216:S_216 <= prev_S_of_j; 
		'd217:S_217 <= prev_S_of_j; 
		'd218:S_218 <= prev_S_of_j; 
		'd219:S_219 <= prev_S_of_j; 
		'd220:S_220 <= prev_S_of_j; 
		'd221:S_221 <= prev_S_of_j; 
		'd222:S_222 <= prev_S_of_j; 
		'd223:S_223 <= prev_S_of_j; 
		'd224:S_224 <= prev_S_of_j; 
		'd225:S_225 <= prev_S_of_j; 
		'd226:S_226 <= prev_S_of_j; 
		'd227:S_227 <= prev_S_of_j; 
		'd228:S_228 <= prev_S_of_j; 
		'd229:S_229 <= prev_S_of_j; 
		'd230:S_230 <= prev_S_of_j; 
		'd231:S_231 <= prev_S_of_j; 
		'd232:S_232 <= prev_S_of_j; 
		'd233:S_233 <= prev_S_of_j; 
		'd234:S_234 <= prev_S_of_j; 
		'd235:S_235 <= prev_S_of_j; 
		'd236:S_236 <= prev_S_of_j; 
		'd237:S_237 <= prev_S_of_j; 
		'd238:S_238 <= prev_S_of_j; 
		'd239:S_239 <= prev_S_of_j; 
		'd240:S_240 <= prev_S_of_j; 
		'd241:S_241 <= prev_S_of_j; 
		'd242:S_242 <= prev_S_of_j; 
		'd243:S_243 <= prev_S_of_j; 
		'd244:S_244 <= prev_S_of_j; 
		'd245:S_245 <= prev_S_of_j; 
		'd246:S_246 <= prev_S_of_j; 
		'd247:S_247 <= prev_S_of_j; 
		'd248:S_248 <= prev_S_of_j; 
		'd249:S_249 <= prev_S_of_j; 
		'd250:S_250 <= prev_S_of_j; 
		'd251:S_251 <= prev_S_of_j; 
		'd252:S_252 <= prev_S_of_j; 
		'd253:S_253 <= prev_S_of_j; 
		'd254:S_254 <= prev_S_of_j; 
		'd255:S_255 <= prev_S_of_j; 
		default:S_256 <= prev_S_of_j; 
	endcase
				case (KSState)
					4'h5:    KSState <= 4'h2;
					4'h6:    KSState <= 4'h3;
					4'h7: KSState <= 4'h4;
				endcase
			end
		endcase
	end
end

endmodule

