
// Copyright (C) 2014 John Leitch (johnleitch@outlook.com)

// This program is free software: you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation, either version 3 of the License, or
// (at your option) any later version.

// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.

// You should have received a copy of the GNU General Public License
// along with this program.  If not, see <http://www.gnu.org/licenses/>.




module Md5Core ( clk,
 wb,
 a0,
 b0,
 c0,
 d0,
 a64,
 b64,
 c64,
 d64);
input clk;
input [511:0] wb;
input [31:0] a0;
input [31:0] b0;
input [31:0] c0;
input [31:0] d0;
output [31:0] a64;
reg    [31:0] a64;
output [31:0] b64;
reg    [31:0] b64;
output [31:0] c64;
reg    [31:0] c64;
output [31:0] d64;
reg    [31:0] d64;



  wire [31:0] w0_0;
wire [31:0] w0_1;
wire [31:0] w0_2;
wire [31:0] w0_3;
wire [31:0] w0_4;
wire [31:0] w0_5;
wire [31:0] w0_6;
wire [31:0] w0_7;
wire [31:0] w0_8;
wire [31:0] w0_9;
wire [31:0] w0_10;
wire [31:0] w0_11;
wire [31:0] w0_12;
wire [31:0] w0_13;
wire [31:0] w0_14;
wire [31:0] w0_15;

  assign w0_0 = wb[31:0];
  assign w0_1 = wb[63:32];
  assign w0_2 = wb[95:64];
  assign w0_3 = wb[127:96];
  assign w0_4 = wb[159:128];
  assign w0_5 = wb[191:160];
  assign w0_6 = wb[223:192];
  assign w0_7 = wb[255:224];
  assign w0_8 = wb[287:256];
  assign w0_9 = wb[319:288];
  assign w0_10 = wb[351:320];
  assign w0_11 = wb[383:352];
  assign w0_12 = wb[415:384];
  assign w0_13 = wb[447:416];
  assign w0_14 = wb[479:448];
  assign w0_15 = wb[511:480];

  reg [31:0]
  a1, b1, c1, d1,
  a2, b2, c2, d2,
  a3, b3, c3, d3,
  a4, b4, c4, d4,
  a5, b5, c5, d5,
  a6, b6, c6, d6,
  a7, b7, c7, d7,
  a8, b8, c8, d8,
  a9, b9, c9, d9,
  a10, b10, c10, d10,
  a11, b11, c11, d11,
  a12, b12, c12, d12,
  a13, b13, c13, d13,
  a14, b14, c14, d14,
  a15, b15, c15, d15,
  a16, b16, c16, d16,
  a17, b17, c17, d17,
  a18, b18, c18, d18,
  a19, b19, c19, d19,
  a20, b20, c20, d20,
  a21, b21, c21, d21,
  a22, b22, c22, d22,
  a23, b23, c23, d23,
  a24, b24, c24, d24,
  a25, b25, c25, d25,
  a26, b26, c26, d26,
  a27, b27, c27, d27,
  a28, b28, c28, d28,
  a29, b29, c29, d29,
  a30, b30, c30, d30,
  a31, b31, c31, d31,
  a32, b32, c32, d32,
  a33, b33, c33, d33,
  a34, b34, c34, d34,
  a35, b35, c35, d35,
  a36, b36, c36, d36,
  a37, b37, c37, d37,
  a38, b38, c38, d38,
  a39, b39, c39, d39,
  a40, b40, c40, d40,
  a41, b41, c41, d41,
  a42, b42, c42, d42,
  a43, b43, c43, d43,
  a44, b44, c44, d44,
  a45, b45, c45, d45,
  a46, b46, c46, d46,
  a47, b47, c47, d47,
  a48, b48, c48, d48,
  a49, b49, c49, d49,
  a50, b50, c50, d50,
  a51, b51, c51, d51,
  a52, b52, c52, d52,
  a53, b53, c53, d53,
  a54, b54, c54, d54,
  a55, b55, c55, d55,
  a56, b56, c56, d56,
  a57, b57, c57, d57,
  a58, b58, c58, d58,
  a59, b59, c59, d59,
  a60, b60, c60, d60,
  a61, b61, c61, d61,
  a62, b62, c62, d62,
  a63, b63, c63, d63;

  reg [31:0] w1_0;
reg [31:0] w1_1;
reg [31:0] w1_2;
reg [31:0] w1_3;
reg [31:0] w1_4;
reg [31:0] w1_5;
reg [31:0] w1_6;
reg [31:0] w1_7;
reg [31:0] w1_8;
reg [31:0] w1_9;
reg [31:0] w1_10;
reg [31:0] w1_11;
reg [31:0] w1_12;
reg [31:0] w1_13;
reg [31:0] w1_14;
reg [31:0] w1_15;

  reg [31:0] w2_0;
reg [31:0] w2_1;
reg [31:0] w2_2;
reg [31:0] w2_3;
reg [31:0] w2_4;
reg [31:0] w2_5;
reg [31:0] w2_6;
reg [31:0] w2_7;
reg [31:0] w2_8;
reg [31:0] w2_9;
reg [31:0] w2_10;
reg [31:0] w2_11;
reg [31:0] w2_12;
reg [31:0] w2_13;
reg [31:0] w2_14;
reg [31:0] w2_15;

  reg [31:0] w3_0;
reg [31:0] w3_1;
reg [31:0] w3_2;
reg [31:0] w3_3;
reg [31:0] w3_4;
reg [31:0] w3_5;
reg [31:0] w3_6;
reg [31:0] w3_7;
reg [31:0] w3_8;
reg [31:0] w3_9;
reg [31:0] w3_10;
reg [31:0] w3_11;
reg [31:0] w3_12;
reg [31:0] w3_13;
reg [31:0] w3_14;
reg [31:0] w3_15;

  reg [31:0] w4_0;
reg [31:0] w4_1;
reg [31:0] w4_2;
reg [31:0] w4_3;
reg [31:0] w4_4;
reg [31:0] w4_5;
reg [31:0] w4_6;
reg [31:0] w4_7;
reg [31:0] w4_8;
reg [31:0] w4_9;
reg [31:0] w4_10;
reg [31:0] w4_11;
reg [31:0] w4_12;
reg [31:0] w4_13;
reg [31:0] w4_14;
reg [31:0] w4_15;

  reg [31:0] w5_0;
reg [31:0] w5_1;
reg [31:0] w5_2;
reg [31:0] w5_3;
reg [31:0] w5_4;
reg [31:0] w5_5;
reg [31:0] w5_6;
reg [31:0] w5_7;
reg [31:0] w5_8;
reg [31:0] w5_9;
reg [31:0] w5_10;
reg [31:0] w5_11;
reg [31:0] w5_12;
reg [31:0] w5_13;
reg [31:0] w5_14;
reg [31:0] w5_15;

  reg [31:0] w6_0;
reg [31:0] w6_1;
reg [31:0] w6_2;
reg [31:0] w6_3;
reg [31:0] w6_4;
reg [31:0] w6_5;
reg [31:0] w6_6;
reg [31:0] w6_7;
reg [31:0] w6_8;
reg [31:0] w6_9;
reg [31:0] w6_10;
reg [31:0] w6_11;
reg [31:0] w6_12;
reg [31:0] w6_13;
reg [31:0] w6_14;
reg [31:0] w6_15;

  reg [31:0] w7_0;
reg [31:0] w7_1;
reg [31:0] w7_2;
reg [31:0] w7_3;
reg [31:0] w7_4;
reg [31:0] w7_5;
reg [31:0] w7_6;
reg [31:0] w7_7;
reg [31:0] w7_8;
reg [31:0] w7_9;
reg [31:0] w7_10;
reg [31:0] w7_11;
reg [31:0] w7_12;
reg [31:0] w7_13;
reg [31:0] w7_14;
reg [31:0] w7_15;

  reg [31:0] w8_0;
reg [31:0] w8_1;
reg [31:0] w8_2;
reg [31:0] w8_3;
reg [31:0] w8_4;
reg [31:0] w8_5;
reg [31:0] w8_6;
reg [31:0] w8_7;
reg [31:0] w8_8;
reg [31:0] w8_9;
reg [31:0] w8_10;
reg [31:0] w8_11;
reg [31:0] w8_12;
reg [31:0] w8_13;
reg [31:0] w8_14;
reg [31:0] w8_15;

  reg [31:0] w9_0;
reg [31:0] w9_1;
reg [31:0] w9_2;
reg [31:0] w9_3;
reg [31:0] w9_4;
reg [31:0] w9_5;
reg [31:0] w9_6;
reg [31:0] w9_7;
reg [31:0] w9_8;
reg [31:0] w9_9;
reg [31:0] w9_10;
reg [31:0] w9_11;
reg [31:0] w9_12;
reg [31:0] w9_13;
reg [31:0] w9_14;
reg [31:0] w9_15;

  reg [31:0] w10_0;
reg [31:0] w10_1;
reg [31:0] w10_2;
reg [31:0] w10_3;
reg [31:0] w10_4;
reg [31:0] w10_5;
reg [31:0] w10_6;
reg [31:0] w10_7;
reg [31:0] w10_8;
reg [31:0] w10_9;
reg [31:0] w10_10;
reg [31:0] w10_11;
reg [31:0] w10_12;
reg [31:0] w10_13;
reg [31:0] w10_14;
reg [31:0] w10_15;

  reg [31:0] w11_0;
reg [31:0] w11_1;
reg [31:0] w11_2;
reg [31:0] w11_3;
reg [31:0] w11_4;
reg [31:0] w11_5;
reg [31:0] w11_6;
reg [31:0] w11_7;
reg [31:0] w11_8;
reg [31:0] w11_9;
reg [31:0] w11_10;
reg [31:0] w11_11;
reg [31:0] w11_12;
reg [31:0] w11_13;
reg [31:0] w11_14;
reg [31:0] w11_15;

  reg [31:0] w12_0;
reg [31:0] w12_1;
reg [31:0] w12_2;
reg [31:0] w12_3;
reg [31:0] w12_4;
reg [31:0] w12_5;
reg [31:0] w12_6;
reg [31:0] w12_7;
reg [31:0] w12_8;
reg [31:0] w12_9;
reg [31:0] w12_10;
reg [31:0] w12_11;
reg [31:0] w12_12;
reg [31:0] w12_13;
reg [31:0] w12_14;
reg [31:0] w12_15;

  reg [31:0] w13_0;
reg [31:0] w13_1;
reg [31:0] w13_2;
reg [31:0] w13_3;
reg [31:0] w13_4;
reg [31:0] w13_5;
reg [31:0] w13_6;
reg [31:0] w13_7;
reg [31:0] w13_8;
reg [31:0] w13_9;
reg [31:0] w13_10;
reg [31:0] w13_11;
reg [31:0] w13_12;
reg [31:0] w13_13;
reg [31:0] w13_14;
reg [31:0] w13_15;

  reg [31:0] w14_0;
reg [31:0] w14_1;
reg [31:0] w14_2;
reg [31:0] w14_3;
reg [31:0] w14_4;
reg [31:0] w14_5;
reg [31:0] w14_6;
reg [31:0] w14_7;
reg [31:0] w14_8;
reg [31:0] w14_9;
reg [31:0] w14_10;
reg [31:0] w14_11;
reg [31:0] w14_12;
reg [31:0] w14_13;
reg [31:0] w14_14;
reg [31:0] w14_15;

  reg [31:0] w15_0;
reg [31:0] w15_1;
reg [31:0] w15_2;
reg [31:0] w15_3;
reg [31:0] w15_4;
reg [31:0] w15_5;
reg [31:0] w15_6;
reg [31:0] w15_7;
reg [31:0] w15_8;
reg [31:0] w15_9;
reg [31:0] w15_10;
reg [31:0] w15_11;
reg [31:0] w15_12;
reg [31:0] w15_13;
reg [31:0] w15_14;
reg [31:0] w15_15;

  reg [31:0] w16_0;
reg [31:0] w16_1;
reg [31:0] w16_2;
reg [31:0] w16_3;
reg [31:0] w16_4;
reg [31:0] w16_5;
reg [31:0] w16_6;
reg [31:0] w16_7;
reg [31:0] w16_8;
reg [31:0] w16_9;
reg [31:0] w16_10;
reg [31:0] w16_11;
reg [31:0] w16_12;
reg [31:0] w16_13;
reg [31:0] w16_14;
reg [31:0] w16_15;

  reg [31:0] w17_0;
reg [31:0] w17_1;
reg [31:0] w17_2;
reg [31:0] w17_3;
reg [31:0] w17_4;
reg [31:0] w17_5;
reg [31:0] w17_6;
reg [31:0] w17_7;
reg [31:0] w17_8;
reg [31:0] w17_9;
reg [31:0] w17_10;
reg [31:0] w17_11;
reg [31:0] w17_12;
reg [31:0] w17_13;
reg [31:0] w17_14;
reg [31:0] w17_15;

  reg [31:0] w18_0;
reg [31:0] w18_1;
reg [31:0] w18_2;
reg [31:0] w18_3;
reg [31:0] w18_4;
reg [31:0] w18_5;
reg [31:0] w18_6;
reg [31:0] w18_7;
reg [31:0] w18_8;
reg [31:0] w18_9;
reg [31:0] w18_10;
reg [31:0] w18_11;
reg [31:0] w18_12;
reg [31:0] w18_13;
reg [31:0] w18_14;
reg [31:0] w18_15;

  reg [31:0] w19_0;
reg [31:0] w19_1;
reg [31:0] w19_2;
reg [31:0] w19_3;
reg [31:0] w19_4;
reg [31:0] w19_5;
reg [31:0] w19_6;
reg [31:0] w19_7;
reg [31:0] w19_8;
reg [31:0] w19_9;
reg [31:0] w19_10;
reg [31:0] w19_11;
reg [31:0] w19_12;
reg [31:0] w19_13;
reg [31:0] w19_14;
reg [31:0] w19_15;

  reg [31:0] w20_0;
reg [31:0] w20_1;
reg [31:0] w20_2;
reg [31:0] w20_3;
reg [31:0] w20_4;
reg [31:0] w20_5;
reg [31:0] w20_6;
reg [31:0] w20_7;
reg [31:0] w20_8;
reg [31:0] w20_9;
reg [31:0] w20_10;
reg [31:0] w20_11;
reg [31:0] w20_12;
reg [31:0] w20_13;
reg [31:0] w20_14;
reg [31:0] w20_15;

  reg [31:0] w21_0;
reg [31:0] w21_1;
reg [31:0] w21_2;
reg [31:0] w21_3;
reg [31:0] w21_4;
reg [31:0] w21_5;
reg [31:0] w21_6;
reg [31:0] w21_7;
reg [31:0] w21_8;
reg [31:0] w21_9;
reg [31:0] w21_10;
reg [31:0] w21_11;
reg [31:0] w21_12;
reg [31:0] w21_13;
reg [31:0] w21_14;
reg [31:0] w21_15;

  reg [31:0] w22_0;
reg [31:0] w22_1;
reg [31:0] w22_2;
reg [31:0] w22_3;
reg [31:0] w22_4;
reg [31:0] w22_5;
reg [31:0] w22_6;
reg [31:0] w22_7;
reg [31:0] w22_8;
reg [31:0] w22_9;
reg [31:0] w22_10;
reg [31:0] w22_11;
reg [31:0] w22_12;
reg [31:0] w22_13;
reg [31:0] w22_14;
reg [31:0] w22_15;

  reg [31:0] w23_0;
reg [31:0] w23_1;
reg [31:0] w23_2;
reg [31:0] w23_3;
reg [31:0] w23_4;
reg [31:0] w23_5;
reg [31:0] w23_6;
reg [31:0] w23_7;
reg [31:0] w23_8;
reg [31:0] w23_9;
reg [31:0] w23_10;
reg [31:0] w23_11;
reg [31:0] w23_12;
reg [31:0] w23_13;
reg [31:0] w23_14;
reg [31:0] w23_15;

  reg [31:0] w24_0;
reg [31:0] w24_1;
reg [31:0] w24_2;
reg [31:0] w24_3;
reg [31:0] w24_4;
reg [31:0] w24_5;
reg [31:0] w24_6;
reg [31:0] w24_7;
reg [31:0] w24_8;
reg [31:0] w24_9;
reg [31:0] w24_10;
reg [31:0] w24_11;
reg [31:0] w24_12;
reg [31:0] w24_13;
reg [31:0] w24_14;
reg [31:0] w24_15;

  reg [31:0] w25_0;
reg [31:0] w25_1;
reg [31:0] w25_2;
reg [31:0] w25_3;
reg [31:0] w25_4;
reg [31:0] w25_5;
reg [31:0] w25_6;
reg [31:0] w25_7;
reg [31:0] w25_8;
reg [31:0] w25_9;
reg [31:0] w25_10;
reg [31:0] w25_11;
reg [31:0] w25_12;
reg [31:0] w25_13;
reg [31:0] w25_14;
reg [31:0] w25_15;

  reg [31:0] w26_0;
reg [31:0] w26_1;
reg [31:0] w26_2;
reg [31:0] w26_3;
reg [31:0] w26_4;
reg [31:0] w26_5;
reg [31:0] w26_6;
reg [31:0] w26_7;
reg [31:0] w26_8;
reg [31:0] w26_9;
reg [31:0] w26_10;
reg [31:0] w26_11;
reg [31:0] w26_12;
reg [31:0] w26_13;
reg [31:0] w26_14;
reg [31:0] w26_15;

  reg [31:0] w27_0;
reg [31:0] w27_1;
reg [31:0] w27_2;
reg [31:0] w27_3;
reg [31:0] w27_4;
reg [31:0] w27_5;
reg [31:0] w27_6;
reg [31:0] w27_7;
reg [31:0] w27_8;
reg [31:0] w27_9;
reg [31:0] w27_10;
reg [31:0] w27_11;
reg [31:0] w27_12;
reg [31:0] w27_13;
reg [31:0] w27_14;
reg [31:0] w27_15;

  reg [31:0] w28_0;
reg [31:0] w28_1;
reg [31:0] w28_2;
reg [31:0] w28_3;
reg [31:0] w28_4;
reg [31:0] w28_5;
reg [31:0] w28_6;
reg [31:0] w28_7;
reg [31:0] w28_8;
reg [31:0] w28_9;
reg [31:0] w28_10;
reg [31:0] w28_11;
reg [31:0] w28_12;
reg [31:0] w28_13;
reg [31:0] w28_14;
reg [31:0] w28_15;

  reg [31:0] w29_0;
reg [31:0] w29_1;
reg [31:0] w29_2;
reg [31:0] w29_3;
reg [31:0] w29_4;
reg [31:0] w29_5;
reg [31:0] w29_6;
reg [31:0] w29_7;
reg [31:0] w29_8;
reg [31:0] w29_9;
reg [31:0] w29_10;
reg [31:0] w29_11;
reg [31:0] w29_12;
reg [31:0] w29_13;
reg [31:0] w29_14;
reg [31:0] w29_15;

  reg [31:0] w30_0;
reg [31:0] w30_1;
reg [31:0] w30_2;
reg [31:0] w30_3;
reg [31:0] w30_4;
reg [31:0] w30_5;
reg [31:0] w30_6;
reg [31:0] w30_7;
reg [31:0] w30_8;
reg [31:0] w30_9;
reg [31:0] w30_10;
reg [31:0] w30_11;
reg [31:0] w30_12;
reg [31:0] w30_13;
reg [31:0] w30_14;
reg [31:0] w30_15;

  reg [31:0] w31_0;
reg [31:0] w31_1;
reg [31:0] w31_2;
reg [31:0] w31_3;
reg [31:0] w31_4;
reg [31:0] w31_5;
reg [31:0] w31_6;
reg [31:0] w31_7;
reg [31:0] w31_8;
reg [31:0] w31_9;
reg [31:0] w31_10;
reg [31:0] w31_11;
reg [31:0] w31_12;
reg [31:0] w31_13;
reg [31:0] w31_14;
reg [31:0] w31_15;

  reg [31:0] w32_0;
reg [31:0] w32_1;
reg [31:0] w32_2;
reg [31:0] w32_3;
reg [31:0] w32_4;
reg [31:0] w32_5;
reg [31:0] w32_6;
reg [31:0] w32_7;
reg [31:0] w32_8;
reg [31:0] w32_9;
reg [31:0] w32_10;
reg [31:0] w32_11;
reg [31:0] w32_12;
reg [31:0] w32_13;
reg [31:0] w32_14;
reg [31:0] w32_15;

  reg [31:0] w33_0;
reg [31:0] w33_1;
reg [31:0] w33_2;
reg [31:0] w33_3;
reg [31:0] w33_4;
reg [31:0] w33_5;
reg [31:0] w33_6;
reg [31:0] w33_7;
reg [31:0] w33_8;
reg [31:0] w33_9;
reg [31:0] w33_10;
reg [31:0] w33_11;
reg [31:0] w33_12;
reg [31:0] w33_13;
reg [31:0] w33_14;
reg [31:0] w33_15;

  reg [31:0] w34_0;
reg [31:0] w34_1;
reg [31:0] w34_2;
reg [31:0] w34_3;
reg [31:0] w34_4;
reg [31:0] w34_5;
reg [31:0] w34_6;
reg [31:0] w34_7;
reg [31:0] w34_8;
reg [31:0] w34_9;
reg [31:0] w34_10;
reg [31:0] w34_11;
reg [31:0] w34_12;
reg [31:0] w34_13;
reg [31:0] w34_14;
reg [31:0] w34_15;

  reg [31:0] w35_0;
reg [31:0] w35_1;
reg [31:0] w35_2;
reg [31:0] w35_3;
reg [31:0] w35_4;
reg [31:0] w35_5;
reg [31:0] w35_6;
reg [31:0] w35_7;
reg [31:0] w35_8;
reg [31:0] w35_9;
reg [31:0] w35_10;
reg [31:0] w35_11;
reg [31:0] w35_12;
reg [31:0] w35_13;
reg [31:0] w35_14;
reg [31:0] w35_15;

  reg [31:0] w36_0;
reg [31:0] w36_1;
reg [31:0] w36_2;
reg [31:0] w36_3;
reg [31:0] w36_4;
reg [31:0] w36_5;
reg [31:0] w36_6;
reg [31:0] w36_7;
reg [31:0] w36_8;
reg [31:0] w36_9;
reg [31:0] w36_10;
reg [31:0] w36_11;
reg [31:0] w36_12;
reg [31:0] w36_13;
reg [31:0] w36_14;
reg [31:0] w36_15;

  reg [31:0] w37_0;
reg [31:0] w37_1;
reg [31:0] w37_2;
reg [31:0] w37_3;
reg [31:0] w37_4;
reg [31:0] w37_5;
reg [31:0] w37_6;
reg [31:0] w37_7;
reg [31:0] w37_8;
reg [31:0] w37_9;
reg [31:0] w37_10;
reg [31:0] w37_11;
reg [31:0] w37_12;
reg [31:0] w37_13;
reg [31:0] w37_14;
reg [31:0] w37_15;

  reg [31:0] w38_0;
reg [31:0] w38_1;
reg [31:0] w38_2;
reg [31:0] w38_3;
reg [31:0] w38_4;
reg [31:0] w38_5;
reg [31:0] w38_6;
reg [31:0] w38_7;
reg [31:0] w38_8;
reg [31:0] w38_9;
reg [31:0] w38_10;
reg [31:0] w38_11;
reg [31:0] w38_12;
reg [31:0] w38_13;
reg [31:0] w38_14;
reg [31:0] w38_15;

  reg [31:0] w39_0;
reg [31:0] w39_1;
reg [31:0] w39_2;
reg [31:0] w39_3;
reg [31:0] w39_4;
reg [31:0] w39_5;
reg [31:0] w39_6;
reg [31:0] w39_7;
reg [31:0] w39_8;
reg [31:0] w39_9;
reg [31:0] w39_10;
reg [31:0] w39_11;
reg [31:0] w39_12;
reg [31:0] w39_13;
reg [31:0] w39_14;
reg [31:0] w39_15;

  reg [31:0] w40_0;
reg [31:0] w40_1;
reg [31:0] w40_2;
reg [31:0] w40_3;
reg [31:0] w40_4;
reg [31:0] w40_5;
reg [31:0] w40_6;
reg [31:0] w40_7;
reg [31:0] w40_8;
reg [31:0] w40_9;
reg [31:0] w40_10;
reg [31:0] w40_11;
reg [31:0] w40_12;
reg [31:0] w40_13;
reg [31:0] w40_14;
reg [31:0] w40_15;

  reg [31:0] w41_0;
reg [31:0] w41_1;
reg [31:0] w41_2;
reg [31:0] w41_3;
reg [31:0] w41_4;
reg [31:0] w41_5;
reg [31:0] w41_6;
reg [31:0] w41_7;
reg [31:0] w41_8;
reg [31:0] w41_9;
reg [31:0] w41_10;
reg [31:0] w41_11;
reg [31:0] w41_12;
reg [31:0] w41_13;
reg [31:0] w41_14;
reg [31:0] w41_15;

  reg [31:0] w42_0;
reg [31:0] w42_1;
reg [31:0] w42_2;
reg [31:0] w42_3;
reg [31:0] w42_4;
reg [31:0] w42_5;
reg [31:0] w42_6;
reg [31:0] w42_7;
reg [31:0] w42_8;
reg [31:0] w42_9;
reg [31:0] w42_10;
reg [31:0] w42_11;
reg [31:0] w42_12;
reg [31:0] w42_13;
reg [31:0] w42_14;
reg [31:0] w42_15;

  reg [31:0] w43_0;
reg [31:0] w43_1;
reg [31:0] w43_2;
reg [31:0] w43_3;
reg [31:0] w43_4;
reg [31:0] w43_5;
reg [31:0] w43_6;
reg [31:0] w43_7;
reg [31:0] w43_8;
reg [31:0] w43_9;
reg [31:0] w43_10;
reg [31:0] w43_11;
reg [31:0] w43_12;
reg [31:0] w43_13;
reg [31:0] w43_14;
reg [31:0] w43_15;

  reg [31:0] w44_0;
reg [31:0] w44_1;
reg [31:0] w44_2;
reg [31:0] w44_3;
reg [31:0] w44_4;
reg [31:0] w44_5;
reg [31:0] w44_6;
reg [31:0] w44_7;
reg [31:0] w44_8;
reg [31:0] w44_9;
reg [31:0] w44_10;
reg [31:0] w44_11;
reg [31:0] w44_12;
reg [31:0] w44_13;
reg [31:0] w44_14;
reg [31:0] w44_15;

  reg [31:0] w45_0;
reg [31:0] w45_1;
reg [31:0] w45_2;
reg [31:0] w45_3;
reg [31:0] w45_4;
reg [31:0] w45_5;
reg [31:0] w45_6;
reg [31:0] w45_7;
reg [31:0] w45_8;
reg [31:0] w45_9;
reg [31:0] w45_10;
reg [31:0] w45_11;
reg [31:0] w45_12;
reg [31:0] w45_13;
reg [31:0] w45_14;
reg [31:0] w45_15;

  reg [31:0] w46_0;
reg [31:0] w46_1;
reg [31:0] w46_2;
reg [31:0] w46_3;
reg [31:0] w46_4;
reg [31:0] w46_5;
reg [31:0] w46_6;
reg [31:0] w46_7;
reg [31:0] w46_8;
reg [31:0] w46_9;
reg [31:0] w46_10;
reg [31:0] w46_11;
reg [31:0] w46_12;
reg [31:0] w46_13;
reg [31:0] w46_14;
reg [31:0] w46_15;

  reg [31:0] w47_0;
reg [31:0] w47_1;
reg [31:0] w47_2;
reg [31:0] w47_3;
reg [31:0] w47_4;
reg [31:0] w47_5;
reg [31:0] w47_6;
reg [31:0] w47_7;
reg [31:0] w47_8;
reg [31:0] w47_9;
reg [31:0] w47_10;
reg [31:0] w47_11;
reg [31:0] w47_12;
reg [31:0] w47_13;
reg [31:0] w47_14;
reg [31:0] w47_15;

  reg [31:0] w48_0;
reg [31:0] w48_1;
reg [31:0] w48_2;
reg [31:0] w48_3;
reg [31:0] w48_4;
reg [31:0] w48_5;
reg [31:0] w48_6;
reg [31:0] w48_7;
reg [31:0] w48_8;
reg [31:0] w48_9;
reg [31:0] w48_10;
reg [31:0] w48_11;
reg [31:0] w48_12;
reg [31:0] w48_13;
reg [31:0] w48_14;
reg [31:0] w48_15;

  reg [31:0] w49_0;
reg [31:0] w49_1;
reg [31:0] w49_2;
reg [31:0] w49_3;
reg [31:0] w49_4;
reg [31:0] w49_5;
reg [31:0] w49_6;
reg [31:0] w49_7;
reg [31:0] w49_8;
reg [31:0] w49_9;
reg [31:0] w49_10;
reg [31:0] w49_11;
reg [31:0] w49_12;
reg [31:0] w49_13;
reg [31:0] w49_14;
reg [31:0] w49_15;

  reg [31:0] w50_0;
reg [31:0] w50_1;
reg [31:0] w50_2;
reg [31:0] w50_3;
reg [31:0] w50_4;
reg [31:0] w50_5;
reg [31:0] w50_6;
reg [31:0] w50_7;
reg [31:0] w50_8;
reg [31:0] w50_9;
reg [31:0] w50_10;
reg [31:0] w50_11;
reg [31:0] w50_12;
reg [31:0] w50_13;
reg [31:0] w50_14;
reg [31:0] w50_15;

  reg [31:0] w51_0;
reg [31:0] w51_1;
reg [31:0] w51_2;
reg [31:0] w51_3;
reg [31:0] w51_4;
reg [31:0] w51_5;
reg [31:0] w51_6;
reg [31:0] w51_7;
reg [31:0] w51_8;
reg [31:0] w51_9;
reg [31:0] w51_10;
reg [31:0] w51_11;
reg [31:0] w51_12;
reg [31:0] w51_13;
reg [31:0] w51_14;
reg [31:0] w51_15;

  reg [31:0] w52_0;
reg [31:0] w52_1;
reg [31:0] w52_2;
reg [31:0] w52_3;
reg [31:0] w52_4;
reg [31:0] w52_5;
reg [31:0] w52_6;
reg [31:0] w52_7;
reg [31:0] w52_8;
reg [31:0] w52_9;
reg [31:0] w52_10;
reg [31:0] w52_11;
reg [31:0] w52_12;
reg [31:0] w52_13;
reg [31:0] w52_14;
reg [31:0] w52_15;

  reg [31:0] w53_0;
reg [31:0] w53_1;
reg [31:0] w53_2;
reg [31:0] w53_3;
reg [31:0] w53_4;
reg [31:0] w53_5;
reg [31:0] w53_6;
reg [31:0] w53_7;
reg [31:0] w53_8;
reg [31:0] w53_9;
reg [31:0] w53_10;
reg [31:0] w53_11;
reg [31:0] w53_12;
reg [31:0] w53_13;
reg [31:0] w53_14;
reg [31:0] w53_15;

  reg [31:0] w54_0;
reg [31:0] w54_1;
reg [31:0] w54_2;
reg [31:0] w54_3;
reg [31:0] w54_4;
reg [31:0] w54_5;
reg [31:0] w54_6;
reg [31:0] w54_7;
reg [31:0] w54_8;
reg [31:0] w54_9;
reg [31:0] w54_10;
reg [31:0] w54_11;
reg [31:0] w54_12;
reg [31:0] w54_13;
reg [31:0] w54_14;
reg [31:0] w54_15;

  reg [31:0] w55_0;
reg [31:0] w55_1;
reg [31:0] w55_2;
reg [31:0] w55_3;
reg [31:0] w55_4;
reg [31:0] w55_5;
reg [31:0] w55_6;
reg [31:0] w55_7;
reg [31:0] w55_8;
reg [31:0] w55_9;
reg [31:0] w55_10;
reg [31:0] w55_11;
reg [31:0] w55_12;
reg [31:0] w55_13;
reg [31:0] w55_14;
reg [31:0] w55_15;

  reg [31:0] w56_0;
reg [31:0] w56_1;
reg [31:0] w56_2;
reg [31:0] w56_3;
reg [31:0] w56_4;
reg [31:0] w56_5;
reg [31:0] w56_6;
reg [31:0] w56_7;
reg [31:0] w56_8;
reg [31:0] w56_9;
reg [31:0] w56_10;
reg [31:0] w56_11;
reg [31:0] w56_12;
reg [31:0] w56_13;
reg [31:0] w56_14;
reg [31:0] w56_15;

  reg [31:0] w57_0;
reg [31:0] w57_1;
reg [31:0] w57_2;
reg [31:0] w57_3;
reg [31:0] w57_4;
reg [31:0] w57_5;
reg [31:0] w57_6;
reg [31:0] w57_7;
reg [31:0] w57_8;
reg [31:0] w57_9;
reg [31:0] w57_10;
reg [31:0] w57_11;
reg [31:0] w57_12;
reg [31:0] w57_13;
reg [31:0] w57_14;
reg [31:0] w57_15;

  reg [31:0] w58_0;
reg [31:0] w58_1;
reg [31:0] w58_2;
reg [31:0] w58_3;
reg [31:0] w58_4;
reg [31:0] w58_5;
reg [31:0] w58_6;
reg [31:0] w58_7;
reg [31:0] w58_8;
reg [31:0] w58_9;
reg [31:0] w58_10;
reg [31:0] w58_11;
reg [31:0] w58_12;
reg [31:0] w58_13;
reg [31:0] w58_14;
reg [31:0] w58_15;

  reg [31:0] w59_0;
reg [31:0] w59_1;
reg [31:0] w59_2;
reg [31:0] w59_3;
reg [31:0] w59_4;
reg [31:0] w59_5;
reg [31:0] w59_6;
reg [31:0] w59_7;
reg [31:0] w59_8;
reg [31:0] w59_9;
reg [31:0] w59_10;
reg [31:0] w59_11;
reg [31:0] w59_12;
reg [31:0] w59_13;
reg [31:0] w59_14;
reg [31:0] w59_15;

  reg [31:0] w60_0;
reg [31:0] w60_1;
reg [31:0] w60_2;
reg [31:0] w60_3;
reg [31:0] w60_4;
reg [31:0] w60_5;
reg [31:0] w60_6;
reg [31:0] w60_7;
reg [31:0] w60_8;
reg [31:0] w60_9;
reg [31:0] w60_10;
reg [31:0] w60_11;
reg [31:0] w60_12;
reg [31:0] w60_13;
reg [31:0] w60_14;
reg [31:0] w60_15;

  reg [31:0] w61_0;
reg [31:0] w61_1;
reg [31:0] w61_2;
reg [31:0] w61_3;
reg [31:0] w61_4;
reg [31:0] w61_5;
reg [31:0] w61_6;
reg [31:0] w61_7;
reg [31:0] w61_8;
reg [31:0] w61_9;
reg [31:0] w61_10;
reg [31:0] w61_11;
reg [31:0] w61_12;
reg [31:0] w61_13;
reg [31:0] w61_14;
reg [31:0] w61_15;

  reg [31:0] w62_0;
reg [31:0] w62_1;
reg [31:0] w62_2;
reg [31:0] w62_3;
reg [31:0] w62_4;
reg [31:0] w62_5;
reg [31:0] w62_6;
reg [31:0] w62_7;
reg [31:0] w62_8;
reg [31:0] w62_9;
reg [31:0] w62_10;
reg [31:0] w62_11;
reg [31:0] w62_12;
reg [31:0] w62_13;
reg [31:0] w62_14;
reg [31:0] w62_15;

  reg [31:0] w63_0;
reg [31:0] w63_1;
reg [31:0] w63_2;
reg [31:0] w63_3;
reg [31:0] w63_4;
reg [31:0] w63_5;
reg [31:0] w63_6;
reg [31:0] w63_7;
reg [31:0] w63_8;
reg [31:0] w63_9;
reg [31:0] w63_10;
reg [31:0] w63_11;
reg [31:0] w63_12;
reg [31:0] w63_13;
reg [31:0] w63_14;
reg [31:0] w63_15;


  always @(posedge clk)
    begin
      a1 <= d0;                                                     
  d1 <= c0;                                                     
  c1 <= b0;
      b1 <= b0 + ((((a0 + ((b0 & c0) | ((~b0) & d0)) + 'hd76aa478 + w0_0) << 7) | ((a0 + ((b0 & c0) | ((~b0) & d0)) + 'hd76aa478 + w0_0) >> (32 - 7))));
      w1_0 <= w0_0;         
  w1_1 <= w0_1;         
  w1_2 <= w0_2;         
  w1_3 <= w0_3;         
  w1_4 <= w0_4;         
  w1_5 <= w0_5;         
  w1_6 <= w0_6;         
  w1_7 <= w0_7;         
  w1_8 <= w0_8;         
  w1_9 <= w0_9;         
  w1_10 <= w0_10;       
  w1_11 <= w0_11;       
  w1_12 <= w0_12;       
  w1_13 <= w0_13;       
  w1_14 <= w0_14;       
  w1_15 <= w0_15;

      a2 <= d1;                                                     
  d2 <= c1;                                                     
  c2 <= b1;
      b2 <= b1 + (((a1 + ((b1 & c1) | ((~b1) & d1)) + 'he8c7b756 + w1_1) << 12) | ((a1 + ((b1 & c1) | ((~b1) & d1)) + 'he8c7b756 + w1_1) >> (32 - 12)));
      w2_0 <= w1_0;         
  w2_1 <= w1_1;         
  w2_2 <= w1_2;         
  w2_3 <= w1_3;         
  w2_4 <= w1_4;         
  w2_5 <= w1_5;         
  w2_6 <= w1_6;         
  w2_7 <= w1_7;         
  w2_8 <= w1_8;         
  w2_9 <= w1_9;         
  w2_10 <= w1_10;       
  w2_11 <= w1_11;       
  w2_12 <= w1_12;       
  w2_13 <= w1_13;       
  w2_14 <= w1_14;       
  w2_15 <= w1_15;

      a3 <= d2;                                                     
  d3 <= c2;                                                     
  c3 <= b2;
      b3 <= b2 + (((a2 + ((b2 & c2) | ((~b2) & d2)) + 'h242070db + w2_2) << 17) | ((a2 + ((b2 & c2) | ((~b2) & d2)) + 'h242070db + w2_2) >> (32 - 17)));
      w3_0 <= w2_0;         
  w3_1 <= w2_1;         
  w3_2 <= w2_2;         
  w3_3 <= w2_3;         
  w3_4 <= w2_4;         
  w3_5 <= w2_5;         
  w3_6 <= w2_6;         
  w3_7 <= w2_7;         
  w3_8 <= w2_8;         
  w3_9 <= w2_9;         
  w3_10 <= w2_10;       
  w3_11 <= w2_11;       
  w3_12 <= w2_12;       
  w3_13 <= w2_13;       
  w3_14 <= w2_14;       
  w3_15 <= w2_15;

      a4 <= d3;                                                     
  d4 <= c3;                                                     
  c4 <= b3;
      b4 <= b3 + (((a3 + ((b3 & c3) | ((~b3) & d3)) + 'hc1bdceee + w3_3) << 22) | ((a3 + ((b3 & c3) | ((~b3) & d3)) + 'hc1bdceee + w3_3) >> (32 - 22)));
      w4_0 <= w3_0;         
  w4_1 <= w3_1;         
  w4_2 <= w3_2;         
  w4_3 <= w3_3;         
  w4_4 <= w3_4;         
  w4_5 <= w3_5;         
  w4_6 <= w3_6;         
  w4_7 <= w3_7;         
  w4_8 <= w3_8;         
  w4_9 <= w3_9;         
  w4_10 <= w3_10;       
  w4_11 <= w3_11;       
  w4_12 <= w3_12;       
  w4_13 <= w3_13;       
  w4_14 <= w3_14;       
  w4_15 <= w3_15;

      a5 <= d4;                                                     
  d5 <= c4;                                                     
  c5 <= b4;
      b5 <= b4 + (((a4 + ((b4 & c4) | ((~b4) & d4)) + 'hf57c0faf + w4_4) << 7) | ((a4 + ((b4 & c4) | ((~b4) & d4)) + 'hf57c0faf + w4_4) >> (32 - 7)));
      w5_0 <= w4_0;         
  w5_1 <= w4_1;         
  w5_2 <= w4_2;         
  w5_3 <= w4_3;         
  w5_4 <= w4_4;         
  w5_5 <= w4_5;         
  w5_6 <= w4_6;         
  w5_7 <= w4_7;         
  w5_8 <= w4_8;         
  w5_9 <= w4_9;         
  w5_10 <= w4_10;       
  w5_11 <= w4_11;       
  w5_12 <= w4_12;       
  w5_13 <= w4_13;       
  w5_14 <= w4_14;       
  w5_15 <= w4_15;

      a6 <= d5;                                                     
  d6 <= c5;                                                     
  c6 <= b5;
      b6 <= b5 + (((a5 + ((b5 & c5) | ((~b5) & d5)) + 'h4787c62a + w5_5) << 12) | ((a5 + ((b5 & c5) | ((~b5) & d5)) + 'h4787c62a + w5_5) >> (32 - 12)));
      w6_0 <= w5_0;         
  w6_1 <= w5_1;         
  w6_2 <= w5_2;         
  w6_3 <= w5_3;         
  w6_4 <= w5_4;         
  w6_5 <= w5_5;         
  w6_6 <= w5_6;         
  w6_7 <= w5_7;         
  w6_8 <= w5_8;         
  w6_9 <= w5_9;         
  w6_10 <= w5_10;       
  w6_11 <= w5_11;       
  w6_12 <= w5_12;       
  w6_13 <= w5_13;       
  w6_14 <= w5_14;       
  w6_15 <= w5_15;

      a7 <= d6;                                                     
  d7 <= c6;                                                     
  c7 <= b6;
      b7 <= b6 + (((a6 + ((b6 & c6) | ((~b6) & d6)) + 'ha8304613 + w6_6) << 17) | ((a6 + ((b6 & c6) | ((~b6) & d6)) + 'ha8304613 + w6_6) >> (32 - 17)));
      w7_0 <= w6_0;         
  w7_1 <= w6_1;         
  w7_2 <= w6_2;         
  w7_3 <= w6_3;         
  w7_4 <= w6_4;         
  w7_5 <= w6_5;         
  w7_6 <= w6_6;         
  w7_7 <= w6_7;         
  w7_8 <= w6_8;         
  w7_9 <= w6_9;         
  w7_10 <= w6_10;       
  w7_11 <= w6_11;       
  w7_12 <= w6_12;       
  w7_13 <= w6_13;       
  w7_14 <= w6_14;       
  w7_15 <= w6_15;

      a8 <= d7;                                                     
  d8 <= c7;                                                     
  c8 <= b7;
      b8 <= b7 + (((a7 + ((b7 & c7) | ((~b7) & d7)) + 'hfd469501 + w7_7) << 22) | ((a7 + ((b7 & c7) | ((~b7) & d7)) + 'hfd469501 + w7_7) >> (32 - 22)));
      w8_0 <= w7_0;         
  w8_1 <= w7_1;         
  w8_2 <= w7_2;         
  w8_3 <= w7_3;         
  w8_4 <= w7_4;         
  w8_5 <= w7_5;         
  w8_6 <= w7_6;         
  w8_7 <= w7_7;         
  w8_8 <= w7_8;         
  w8_9 <= w7_9;         
  w8_10 <= w7_10;       
  w8_11 <= w7_11;       
  w8_12 <= w7_12;       
  w8_13 <= w7_13;       
  w8_14 <= w7_14;       
  w8_15 <= w7_15;

      a9 <= d8;                                                     
  d9 <= c8;                                                     
  c9 <= b8;
      b9 <= b8 + (((a8 + ((b8 & c8) | ((~b8) & d8)) + 'h698098d8 + w8_8) << 7) | ((a8 + ((b8 & c8) | ((~b8) & d8)) + 'h698098d8 + w8_8) >> (32 - 7)));
      w9_0 <= w8_0;         
  w9_1 <= w8_1;         
  w9_2 <= w8_2;         
  w9_3 <= w8_3;         
  w9_4 <= w8_4;         
  w9_5 <= w8_5;         
  w9_6 <= w8_6;         
  w9_7 <= w8_7;         
  w9_8 <= w8_8;         
  w9_9 <= w8_9;         
  w9_10 <= w8_10;       
  w9_11 <= w8_11;       
  w9_12 <= w8_12;       
  w9_13 <= w8_13;       
  w9_14 <= w8_14;       
  w9_15 <= w8_15;

      a10 <= d9;                                                     
  d10 <= c9;                                                     
  c10 <= b9;
      b10 <= b9 + (((a9 + ((b9 & c9) | ((~b9) & d9)) + 'h8b44f7af + w9_9) << 12) | ((a9 + ((b9 & c9) | ((~b9) & d9)) + 'h8b44f7af + w9_9) >> (32 - 12)));
      w10_0 <= w9_0;         
  w10_1 <= w9_1;         
  w10_2 <= w9_2;         
  w10_3 <= w9_3;         
  w10_4 <= w9_4;         
  w10_5 <= w9_5;         
  w10_6 <= w9_6;         
  w10_7 <= w9_7;         
  w10_8 <= w9_8;         
  w10_9 <= w9_9;         
  w10_10 <= w9_10;       
  w10_11 <= w9_11;       
  w10_12 <= w9_12;       
  w10_13 <= w9_13;       
  w10_14 <= w9_14;       
  w10_15 <= w9_15;

      a11 <= d10;                                                     
  d11 <= c10;                                                     
  c11 <= b10;
      b11 <= b10 + (((a10 + ((b10 & c10) | ((~b10) & d10)) + 'hffff5bb1 + w10_10) << 17) | ((a10 + ((b10 & c10) | ((~b10) & d10)) + 'hffff5bb1 + w10_10) >> (32 - 17)));
      w11_0 <= w10_0;         
  w11_1 <= w10_1;         
  w11_2 <= w10_2;         
  w11_3 <= w10_3;         
  w11_4 <= w10_4;         
  w11_5 <= w10_5;         
  w11_6 <= w10_6;         
  w11_7 <= w10_7;         
  w11_8 <= w10_8;         
  w11_9 <= w10_9;         
  w11_10 <= w10_10;       
  w11_11 <= w10_11;       
  w11_12 <= w10_12;       
  w11_13 <= w10_13;       
  w11_14 <= w10_14;       
  w11_15 <= w10_15;

      a12 <= d11;                                                     
  d12 <= c11;                                                     
  c12 <= b11;
      b12 <= b11 + (((a11 + ((b11 & c11) | ((~b11) & d11)) + 'h895cd7be + w11_11) << 22) | ((a11 + ((b11 & c11) | ((~b11) & d11)) + 'h895cd7be + w11_11) >> (32 - 22)));
      w12_0 <= w11_0;         
  w12_1 <= w11_1;         
  w12_2 <= w11_2;         
  w12_3 <= w11_3;         
  w12_4 <= w11_4;         
  w12_5 <= w11_5;         
  w12_6 <= w11_6;         
  w12_7 <= w11_7;         
  w12_8 <= w11_8;         
  w12_9 <= w11_9;         
  w12_10 <= w11_10;       
  w12_11 <= w11_11;       
  w12_12 <= w11_12;       
  w12_13 <= w11_13;       
  w12_14 <= w11_14;       
  w12_15 <= w11_15;

      a13 <= d12;                                                     
  d13 <= c12;                                                     
  c13 <= b12;
      b13 <= b12 + (((a12 + ((b12 & c12) | ((~b12) & d12)) + 'h6b901122 + w12_12) << 7) | ((a12 + ((b12 & c12) | ((~b12) & d12)) + 'h6b901122 + w12_12) >> (32 - 7)));
      w13_0 <= w12_0;         
  w13_1 <= w12_1;         
  w13_2 <= w12_2;         
  w13_3 <= w12_3;         
  w13_4 <= w12_4;         
  w13_5 <= w12_5;         
  w13_6 <= w12_6;         
  w13_7 <= w12_7;         
  w13_8 <= w12_8;         
  w13_9 <= w12_9;         
  w13_10 <= w12_10;       
  w13_11 <= w12_11;       
  w13_12 <= w12_12;       
  w13_13 <= w12_13;       
  w13_14 <= w12_14;       
  w13_15 <= w12_15;

      a14 <= d13;                                                     
  d14 <= c13;                                                     
  c14 <= b13;
      b14 <= b13 + (((a13 + ((b13 & c13) | ((~b13) & d13)) + 'hfd987193 + w13_13) << 12) | ((a13 + ((b13 & c13) | ((~b13) & d13)) + 'hfd987193 + w13_13) >> (32 - 12)));
      w14_0 <= w13_0;         
  w14_1 <= w13_1;         
  w14_2 <= w13_2;         
  w14_3 <= w13_3;         
  w14_4 <= w13_4;         
  w14_5 <= w13_5;         
  w14_6 <= w13_6;         
  w14_7 <= w13_7;         
  w14_8 <= w13_8;         
  w14_9 <= w13_9;         
  w14_10 <= w13_10;       
  w14_11 <= w13_11;       
  w14_12 <= w13_12;       
  w14_13 <= w13_13;       
  w14_14 <= w13_14;       
  w14_15 <= w13_15;

      a15 <= d14;                                                     
  d15 <= c14;                                                     
  c15 <= b14;
      b15 <= b14 + (((a14 + ((b14 & c14) | ((~b14) & d14)) + 'ha679438e + w14_14) << 17) | ((a14 + ((b14 & c14) | ((~b14) & d14)) + 'ha679438e + w14_14) >> (32 - 17)));
      w15_0 <= w14_0;         
  w15_1 <= w14_1;         
  w15_2 <= w14_2;         
  w15_3 <= w14_3;         
  w15_4 <= w14_4;         
  w15_5 <= w14_5;         
  w15_6 <= w14_6;         
  w15_7 <= w14_7;         
  w15_8 <= w14_8;         
  w15_9 <= w14_9;         
  w15_10 <= w14_10;       
  w15_11 <= w14_11;       
  w15_12 <= w14_12;       
  w15_13 <= w14_13;       
  w15_14 <= w14_14;       
  w15_15 <= w14_15;

      a16 <= d15;                                                     
  d16 <= c15;                                                     
  c16 <= b15;
      b16 <= b15 + (((a15 + ((b15 & c15) | ((~b15) & d15)) + 'h49b40821 + w15_15) << 22) | ((a15 + ((b15 & c15) | ((~b15) & d15)) + 'h49b40821 + w15_15) >> (32 - 22)));
      w16_0 <= w15_0;         
  w16_1 <= w15_1;         
  w16_2 <= w15_2;         
  w16_3 <= w15_3;         
  w16_4 <= w15_4;         
  w16_5 <= w15_5;         
  w16_6 <= w15_6;         
  w16_7 <= w15_7;         
  w16_8 <= w15_8;         
  w16_9 <= w15_9;         
  w16_10 <= w15_10;       
  w16_11 <= w15_11;       
  w16_12 <= w15_12;       
  w16_13 <= w15_13;       
  w16_14 <= w15_14;       
  w16_15 <= w15_15;

      a17 <= d16;                                                     
  d17 <= c16;                                                     
  c17 <= b16;
      b17 <= b16 + (((a16 + ((d16 & b16) | ((~d16) & c16)) + 'hf61e2562 + w16_1) << 5) | ((a16 + ((d16 & b16) | ((~d16) & c16)) + 'hf61e2562 + w16_1) >> (32 - 5)));
      w17_0 <= w16_0;         
  w17_1 <= w16_1;         
  w17_2 <= w16_2;         
  w17_3 <= w16_3;         
  w17_4 <= w16_4;         
  w17_5 <= w16_5;         
  w17_6 <= w16_6;         
  w17_7 <= w16_7;         
  w17_8 <= w16_8;         
  w17_9 <= w16_9;         
  w17_10 <= w16_10;       
  w17_11 <= w16_11;       
  w17_12 <= w16_12;       
  w17_13 <= w16_13;       
  w17_14 <= w16_14;       
  w17_15 <= w16_15;

      a18 <= d17;                                                     
  d18 <= c17;                                                     
  c18 <= b17;
      b18 <= b17 + (((a17 + ((d17 & b17) | ((~d17) & c17)) + 'hc040b340 + w17_6) << 9) | ((a17 + ((d17 & b17) | ((~d17) & c17)) + 'hc040b340 + w17_6) >> (32 - 9)));
      w18_0 <= w17_0;         
  w18_1 <= w17_1;         
  w18_2 <= w17_2;         
  w18_3 <= w17_3;         
  w18_4 <= w17_4;         
  w18_5 <= w17_5;         
  w18_6 <= w17_6;         
  w18_7 <= w17_7;         
  w18_8 <= w17_8;         
  w18_9 <= w17_9;         
  w18_10 <= w17_10;       
  w18_11 <= w17_11;       
  w18_12 <= w17_12;       
  w18_13 <= w17_13;       
  w18_14 <= w17_14;       
  w18_15 <= w17_15;

      a19 <= d18;                                                     
  d19 <= c18;                                                     
  c19 <= b18;
      b19 <= b18 + (((a18 + ((d18 & b18) | ((~d18) & c18)) + 'h265e5a51 + w18_11) << 14) | ((a18 + ((d18 & b18) | ((~d18) & c18)) + 'h265e5a51 + w18_11) >> (32 - 14)));
      w19_0 <= w18_0;         
  w19_1 <= w18_1;         
  w19_2 <= w18_2;         
  w19_3 <= w18_3;         
  w19_4 <= w18_4;         
  w19_5 <= w18_5;         
  w19_6 <= w18_6;         
  w19_7 <= w18_7;         
  w19_8 <= w18_8;         
  w19_9 <= w18_9;         
  w19_10 <= w18_10;       
  w19_11 <= w18_11;       
  w19_12 <= w18_12;       
  w19_13 <= w18_13;       
  w19_14 <= w18_14;       
  w19_15 <= w18_15;

      a20 <= d19;                                                     
  d20 <= c19;                                                     
  c20 <= b19;
      b20 <= b19 + (((a19 + ((d19 & b19) | ((~d19) & c19)) + 'he9b6c7aa + w19_0) << 20) | ((a19 + ((d19 & b19) | ((~d19) & c19)) + 'he9b6c7aa + w19_0) >> (32 - 20)));
      w20_0 <= w19_0;         
  w20_1 <= w19_1;         
  w20_2 <= w19_2;         
  w20_3 <= w19_3;         
  w20_4 <= w19_4;         
  w20_5 <= w19_5;         
  w20_6 <= w19_6;         
  w20_7 <= w19_7;         
  w20_8 <= w19_8;         
  w20_9 <= w19_9;         
  w20_10 <= w19_10;       
  w20_11 <= w19_11;       
  w20_12 <= w19_12;       
  w20_13 <= w19_13;       
  w20_14 <= w19_14;       
  w20_15 <= w19_15;

      a21 <= d20;                                                     
  d21 <= c20;                                                     
  c21 <= b20;
      b21 <= b20 + (((a20 + ((d20 & b20) | ((~d20) & c20)) + 'hd62f105d + w20_5) << 5) | ((a20 + ((d20 & b20) | ((~d20) & c20)) + 'hd62f105d + w20_5) >> (32 - 5)));
      w21_0 <= w20_0;         
  w21_1 <= w20_1;         
  w21_2 <= w20_2;         
  w21_3 <= w20_3;         
  w21_4 <= w20_4;         
  w21_5 <= w20_5;         
  w21_6 <= w20_6;         
  w21_7 <= w20_7;         
  w21_8 <= w20_8;         
  w21_9 <= w20_9;         
  w21_10 <= w20_10;       
  w21_11 <= w20_11;       
  w21_12 <= w20_12;       
  w21_13 <= w20_13;       
  w21_14 <= w20_14;       
  w21_15 <= w20_15;

      a22 <= d21;                                                     
  d22 <= c21;                                                     
  c22 <= b21;
      b22 <= b21 + (((a21 + ((d21 & b21) | ((~d21) & c21)) + 'h02441453 + w21_10) << 9) | ((a21 + ((d21 & b21) | ((~d21) & c21)) + 'h02441453 + w21_10) >> (32 - 9)));
      w22_0 <= w21_0;         
  w22_1 <= w21_1;         
  w22_2 <= w21_2;         
  w22_3 <= w21_3;         
  w22_4 <= w21_4;         
  w22_5 <= w21_5;         
  w22_6 <= w21_6;         
  w22_7 <= w21_7;         
  w22_8 <= w21_8;         
  w22_9 <= w21_9;         
  w22_10 <= w21_10;       
  w22_11 <= w21_11;       
  w22_12 <= w21_12;       
  w22_13 <= w21_13;       
  w22_14 <= w21_14;       
  w22_15 <= w21_15;

      a23 <= d22;                                                     
  d23 <= c22;                                                     
  c23 <= b22;
      b23 <= b22 + (((a22 + ((d22 & b22) | ((~d22) & c22)) + 'hd8a1e681 + w22_15) << 14) | ((a22 + ((d22 & b22) | ((~d22) & c22)) + 'hd8a1e681 + w22_15) >> (32 - 14)));
      w23_0 <= w22_0;         
  w23_1 <= w22_1;         
  w23_2 <= w22_2;         
  w23_3 <= w22_3;         
  w23_4 <= w22_4;         
  w23_5 <= w22_5;         
  w23_6 <= w22_6;         
  w23_7 <= w22_7;         
  w23_8 <= w22_8;         
  w23_9 <= w22_9;         
  w23_10 <= w22_10;       
  w23_11 <= w22_11;       
  w23_12 <= w22_12;       
  w23_13 <= w22_13;       
  w23_14 <= w22_14;       
  w23_15 <= w22_15;

      a24 <= d23;                                                     
  d24 <= c23;                                                     
  c24 <= b23;
      b24 <= b23 + (((a23 + ((d23 & b23) | ((~d23) & c23)) + 'he7d3fbc8 + w23_4) << 20) | ((a23 + ((d23 & b23) | ((~d23) & c23)) + 'he7d3fbc8 + w23_4) >> (32 - 20)));
      w24_0 <= w23_0;         
  w24_1 <= w23_1;         
  w24_2 <= w23_2;         
  w24_3 <= w23_3;         
  w24_4 <= w23_4;         
  w24_5 <= w23_5;         
  w24_6 <= w23_6;         
  w24_7 <= w23_7;         
  w24_8 <= w23_8;         
  w24_9 <= w23_9;         
  w24_10 <= w23_10;       
  w24_11 <= w23_11;       
  w24_12 <= w23_12;       
  w24_13 <= w23_13;       
  w24_14 <= w23_14;       
  w24_15 <= w23_15;

      a25 <= d24;                                                     
  d25 <= c24;                                                     
  c25 <= b24;
      b25 <= b24 + (((a24 + ((d24 & b24) | ((~d24) & c24)) + 'h21e1cde6 + w24_9) << 5) | ((a24 + ((d24 & b24) | ((~d24) & c24)) + 'h21e1cde6 + w24_9) >> (32 - 5)));
      w25_0 <= w24_0;         
  w25_1 <= w24_1;         
  w25_2 <= w24_2;         
  w25_3 <= w24_3;         
  w25_4 <= w24_4;         
  w25_5 <= w24_5;         
  w25_6 <= w24_6;         
  w25_7 <= w24_7;         
  w25_8 <= w24_8;         
  w25_9 <= w24_9;         
  w25_10 <= w24_10;       
  w25_11 <= w24_11;       
  w25_12 <= w24_12;       
  w25_13 <= w24_13;       
  w25_14 <= w24_14;       
  w25_15 <= w24_15;

      a26 <= d25;                                                     
  d26 <= c25;                                                     
  c26 <= b25;
      b26 <= b25 + (((a25 + ((d25 & b25) | ((~d25) & c25)) + 'hc33707d6 + w25_14) << 9) | ((a25 + ((d25 & b25) | ((~d25) & c25)) + 'hc33707d6 + w25_14) >> (32 - 9)));
      w26_0 <= w25_0;         
  w26_1 <= w25_1;         
  w26_2 <= w25_2;         
  w26_3 <= w25_3;         
  w26_4 <= w25_4;         
  w26_5 <= w25_5;         
  w26_6 <= w25_6;         
  w26_7 <= w25_7;         
  w26_8 <= w25_8;         
  w26_9 <= w25_9;         
  w26_10 <= w25_10;       
  w26_11 <= w25_11;       
  w26_12 <= w25_12;       
  w26_13 <= w25_13;       
  w26_14 <= w25_14;       
  w26_15 <= w25_15;

      a27 <= d26;                                                     
  d27 <= c26;                                                     
  c27 <= b26;
      b27 <= b26 + (((a26 + ((d26 & b26) | ((~d26) & c26)) + 'hf4d50d87 + w26_3) << 14) | ((a26 + ((d26 & b26) | ((~d26) & c26)) + 'hf4d50d87 + w26_3) >> (32 - 14)));
      w27_0 <= w26_0;         
  w27_1 <= w26_1;         
  w27_2 <= w26_2;         
  w27_3 <= w26_3;         
  w27_4 <= w26_4;         
  w27_5 <= w26_5;         
  w27_6 <= w26_6;         
  w27_7 <= w26_7;         
  w27_8 <= w26_8;         
  w27_9 <= w26_9;         
  w27_10 <= w26_10;       
  w27_11 <= w26_11;       
  w27_12 <= w26_12;       
  w27_13 <= w26_13;       
  w27_14 <= w26_14;       
  w27_15 <= w26_15;

      a28 <= d27;                                                     
  d28 <= c27;                                                     
  c28 <= b27;
      b28 <= b27 + (((a27 + ((d27 & b27) | ((~d27) & c27)) + 'h455a14ed + w27_8) << 20) | ((a27 + ((d27 & b27) | ((~d27) & c27)) + 'h455a14ed + w27_8) >> (32 - 20)));
      w28_0 <= w27_0;         
  w28_1 <= w27_1;         
  w28_2 <= w27_2;         
  w28_3 <= w27_3;         
  w28_4 <= w27_4;         
  w28_5 <= w27_5;         
  w28_6 <= w27_6;         
  w28_7 <= w27_7;         
  w28_8 <= w27_8;         
  w28_9 <= w27_9;         
  w28_10 <= w27_10;       
  w28_11 <= w27_11;       
  w28_12 <= w27_12;       
  w28_13 <= w27_13;       
  w28_14 <= w27_14;       
  w28_15 <= w27_15;

      a29 <= d28;                                                     
  d29 <= c28;                                                     
  c29 <= b28;
      b29 <= b28 + (((a28 + ((d28 & b28) | ((~d28) & c28)) + 'ha9e3e905 + w28_13) << 5) | ((a28 + ((d28 & b28) | ((~d28) & c28)) + 'ha9e3e905 + w28_13) >> (32 - 5)));
      w29_0 <= w28_0;         
  w29_1 <= w28_1;         
  w29_2 <= w28_2;         
  w29_3 <= w28_3;         
  w29_4 <= w28_4;         
  w29_5 <= w28_5;         
  w29_6 <= w28_6;         
  w29_7 <= w28_7;         
  w29_8 <= w28_8;         
  w29_9 <= w28_9;         
  w29_10 <= w28_10;       
  w29_11 <= w28_11;       
  w29_12 <= w28_12;       
  w29_13 <= w28_13;       
  w29_14 <= w28_14;       
  w29_15 <= w28_15;

      a30 <= d29;                                                     
  d30 <= c29;                                                     
  c30 <= b29;
      b30 <= b29 + (((a29 + ((d29 & b29) | ((~d29) & c29)) + 'hfcefa3f8 + w29_2) << 9) | ((a29 + ((d29 & b29) | ((~d29) & c29)) + 'hfcefa3f8 + w29_2) >> (32 - 9)));
      w30_0 <= w29_0;         
  w30_1 <= w29_1;         
  w30_2 <= w29_2;         
  w30_3 <= w29_3;         
  w30_4 <= w29_4;         
  w30_5 <= w29_5;         
  w30_6 <= w29_6;         
  w30_7 <= w29_7;         
  w30_8 <= w29_8;         
  w30_9 <= w29_9;         
  w30_10 <= w29_10;       
  w30_11 <= w29_11;       
  w30_12 <= w29_12;       
  w30_13 <= w29_13;       
  w30_14 <= w29_14;       
  w30_15 <= w29_15;

      a31 <= d30;                                                     
  d31 <= c30;                                                     
  c31 <= b30;
      b31 <= b30 + (((a30 + ((d30 & b30) | ((~d30) & c30)) + 'h676f02d9 + w30_7) << 14) | ((a30 + ((d30 & b30) | ((~d30) & c30)) + 'h676f02d9 + w30_7) >> (32 - 14)));
      w31_0 <= w30_0;         
  w31_1 <= w30_1;         
  w31_2 <= w30_2;         
  w31_3 <= w30_3;         
  w31_4 <= w30_4;         
  w31_5 <= w30_5;         
  w31_6 <= w30_6;         
  w31_7 <= w30_7;         
  w31_8 <= w30_8;         
  w31_9 <= w30_9;         
  w31_10 <= w30_10;       
  w31_11 <= w30_11;       
  w31_12 <= w30_12;       
  w31_13 <= w30_13;       
  w31_14 <= w30_14;       
  w31_15 <= w30_15;

      a32 <= d31;                                                     
  d32 <= c31;                                                     
  c32 <= b31;
      b32 <= b31 + (((a31 + ((d31 & b31) | ((~d31) & c31)) + 'h8d2a4c8a + w31_12) << 20) | ((a31 + ((d31 & b31) | ((~d31) & c31)) + 'h8d2a4c8a + w31_12) >> (32 - 20)));
      w32_0 <= w31_0;         
  w32_1 <= w31_1;         
  w32_2 <= w31_2;         
  w32_3 <= w31_3;         
  w32_4 <= w31_4;         
  w32_5 <= w31_5;         
  w32_6 <= w31_6;         
  w32_7 <= w31_7;         
  w32_8 <= w31_8;         
  w32_9 <= w31_9;         
  w32_10 <= w31_10;       
  w32_11 <= w31_11;       
  w32_12 <= w31_12;       
  w32_13 <= w31_13;       
  w32_14 <= w31_14;       
  w32_15 <= w31_15;

      a33 <= d32;                                                     
  d33 <= c32;                                                     
  c33 <= b32;
      b33 <= b32 + (((a32 + (b32 ^ c32 ^ d32) + 'hfffa3942 + w32_5) << 4) | ((a32 + (b32 ^ c32 ^ d32) + 'hfffa3942 + w32_5) >> (32 - 4)));
      w33_0 <= w32_0;         
  w33_1 <= w32_1;         
  w33_2 <= w32_2;         
  w33_3 <= w32_3;         
  w33_4 <= w32_4;         
  w33_5 <= w32_5;         
  w33_6 <= w32_6;         
  w33_7 <= w32_7;         
  w33_8 <= w32_8;         
  w33_9 <= w32_9;         
  w33_10 <= w32_10;       
  w33_11 <= w32_11;       
  w33_12 <= w32_12;       
  w33_13 <= w32_13;       
  w33_14 <= w32_14;       
  w33_15 <= w32_15;

      a34 <= d33;                                                     
  d34 <= c33;                                                     
  c34 <= b33;
      b34 <= b33 + (((a33 + (b33 ^ c33 ^ d33) + 'h8771f681 + w33_8) << 11) | ((a33 + (b33 ^ c33 ^ d33) + 'h8771f681 + w33_8) >> (32 - 11)));
      w34_0 <= w33_0;         
  w34_1 <= w33_1;         
  w34_2 <= w33_2;         
  w34_3 <= w33_3;         
  w34_4 <= w33_4;         
  w34_5 <= w33_5;         
  w34_6 <= w33_6;         
  w34_7 <= w33_7;         
  w34_8 <= w33_8;         
  w34_9 <= w33_9;         
  w34_10 <= w33_10;       
  w34_11 <= w33_11;       
  w34_12 <= w33_12;       
  w34_13 <= w33_13;       
  w34_14 <= w33_14;       
  w34_15 <= w33_15;

      a35 <= d34;                                                     
  d35 <= c34;                                                     
  c35 <= b34;
      b35 <= b34 + (((a34 + (b34 ^ c34 ^ d34) + 'h6d9d6122 + w34_11) << 16) | ((a34 + (b34 ^ c34 ^ d34) + 'h6d9d6122 + w34_11) >> (32 - 16)));
      w35_0 <= w34_0;         
  w35_1 <= w34_1;         
  w35_2 <= w34_2;         
  w35_3 <= w34_3;         
  w35_4 <= w34_4;         
  w35_5 <= w34_5;         
  w35_6 <= w34_6;         
  w35_7 <= w34_7;         
  w35_8 <= w34_8;         
  w35_9 <= w34_9;         
  w35_10 <= w34_10;       
  w35_11 <= w34_11;       
  w35_12 <= w34_12;       
  w35_13 <= w34_13;       
  w35_14 <= w34_14;       
  w35_15 <= w34_15;

      a36 <= d35;                                                     
  d36 <= c35;                                                     
  c36 <= b35;
      b36 <= b35 + (((a35 + (b35 ^ c35 ^ d35) + 'hfde5380c + w35_14) << 23) | ((a35 + (b35 ^ c35 ^ d35) + 'hfde5380c + w35_14) >> (32 - 23)));
      w36_0 <= w35_0;         
  w36_1 <= w35_1;         
  w36_2 <= w35_2;         
  w36_3 <= w35_3;         
  w36_4 <= w35_4;         
  w36_5 <= w35_5;         
  w36_6 <= w35_6;         
  w36_7 <= w35_7;         
  w36_8 <= w35_8;         
  w36_9 <= w35_9;         
  w36_10 <= w35_10;       
  w36_11 <= w35_11;       
  w36_12 <= w35_12;       
  w36_13 <= w35_13;       
  w36_14 <= w35_14;       
  w36_15 <= w35_15;

      a37 <= d36;                                                     
  d37 <= c36;                                                     
  c37 <= b36;
      b37 <= b36 + (((a36 + (b36 ^ c36 ^ d36) + 'ha4beea44 + w36_1) << 4) | ((a36 + (b36 ^ c36 ^ d36) + 'ha4beea44 + w36_1) >> (32 - 4)));
      w37_0 <= w36_0;         
  w37_1 <= w36_1;         
  w37_2 <= w36_2;         
  w37_3 <= w36_3;         
  w37_4 <= w36_4;         
  w37_5 <= w36_5;         
  w37_6 <= w36_6;         
  w37_7 <= w36_7;         
  w37_8 <= w36_8;         
  w37_9 <= w36_9;         
  w37_10 <= w36_10;       
  w37_11 <= w36_11;       
  w37_12 <= w36_12;       
  w37_13 <= w36_13;       
  w37_14 <= w36_14;       
  w37_15 <= w36_15;

      a38 <= d37;                                                     
  d38 <= c37;                                                     
  c38 <= b37;
      b38 <= b37 + (((a37 + (b37 ^ c37 ^ d37) + 'h4bdecfa9 + w37_4) << 11) | ((a37 + (b37 ^ c37 ^ d37) + 'h4bdecfa9 + w37_4) >> (32 - 11)));
      w38_0 <= w37_0;         
  w38_1 <= w37_1;         
  w38_2 <= w37_2;         
  w38_3 <= w37_3;         
  w38_4 <= w37_4;         
  w38_5 <= w37_5;         
  w38_6 <= w37_6;         
  w38_7 <= w37_7;         
  w38_8 <= w37_8;         
  w38_9 <= w37_9;         
  w38_10 <= w37_10;       
  w38_11 <= w37_11;       
  w38_12 <= w37_12;       
  w38_13 <= w37_13;       
  w38_14 <= w37_14;       
  w38_15 <= w37_15;

      a39 <= d38;                                                     
  d39 <= c38;                                                     
  c39 <= b38;
      b39 <= b38 + (((a38 + (b38 ^ c38 ^ d38) + 'hf6bb4b60 + w38_7) << 16) | ((a38 + (b38 ^ c38 ^ d38) + 'hf6bb4b60 + w38_7) >> (32 - 16)));
      w39_0 <= w38_0;         
  w39_1 <= w38_1;         
  w39_2 <= w38_2;         
  w39_3 <= w38_3;         
  w39_4 <= w38_4;         
  w39_5 <= w38_5;         
  w39_6 <= w38_6;         
  w39_7 <= w38_7;         
  w39_8 <= w38_8;         
  w39_9 <= w38_9;         
  w39_10 <= w38_10;       
  w39_11 <= w38_11;       
  w39_12 <= w38_12;       
  w39_13 <= w38_13;       
  w39_14 <= w38_14;       
  w39_15 <= w38_15;

      a40 <= d39;                                                     
  d40 <= c39;                                                     
  c40 <= b39;
      b40 <= b39 + (((a39 + (b39 ^ c39 ^ d39) + 'hbebfbc70 + w39_10) << 23) | ((a39 + (b39 ^ c39 ^ d39) + 'hbebfbc70 + w39_10) >> (32 - 23)));
      w40_0 <= w39_0;         
  w40_1 <= w39_1;         
  w40_2 <= w39_2;         
  w40_3 <= w39_3;         
  w40_4 <= w39_4;         
  w40_5 <= w39_5;         
  w40_6 <= w39_6;         
  w40_7 <= w39_7;         
  w40_8 <= w39_8;         
  w40_9 <= w39_9;         
  w40_10 <= w39_10;       
  w40_11 <= w39_11;       
  w40_12 <= w39_12;       
  w40_13 <= w39_13;       
  w40_14 <= w39_14;       
  w40_15 <= w39_15;

      a41 <= d40;                                                     
  d41 <= c40;                                                     
  c41 <= b40;
      b41 <= b40 + (((a40 + (b40 ^ c40 ^ d40) + 'h289b7ec6 + w40_13) << 4) | ((a40 + (b40 ^ c40 ^ d40) + 'h289b7ec6 + w40_13) >> (32 - 4)));
      w41_0 <= w40_0;         
  w41_1 <= w40_1;         
  w41_2 <= w40_2;         
  w41_3 <= w40_3;         
  w41_4 <= w40_4;         
  w41_5 <= w40_5;         
  w41_6 <= w40_6;         
  w41_7 <= w40_7;         
  w41_8 <= w40_8;         
  w41_9 <= w40_9;         
  w41_10 <= w40_10;       
  w41_11 <= w40_11;       
  w41_12 <= w40_12;       
  w41_13 <= w40_13;       
  w41_14 <= w40_14;       
  w41_15 <= w40_15;

      a42 <= d41;                                                     
  d42 <= c41;                                                     
  c42 <= b41;
      b42 <= b41 + (((a41 + (b41 ^ c41 ^ d41) + 'heaa127fa + w41_0) << 11) | ((a41 + (b41 ^ c41 ^ d41) + 'heaa127fa + w41_0) >> (32 - 11)));
      w42_0 <= w41_0;         
  w42_1 <= w41_1;         
  w42_2 <= w41_2;         
  w42_3 <= w41_3;         
  w42_4 <= w41_4;         
  w42_5 <= w41_5;         
  w42_6 <= w41_6;         
  w42_7 <= w41_7;         
  w42_8 <= w41_8;         
  w42_9 <= w41_9;         
  w42_10 <= w41_10;       
  w42_11 <= w41_11;       
  w42_12 <= w41_12;       
  w42_13 <= w41_13;       
  w42_14 <= w41_14;       
  w42_15 <= w41_15;

      a43 <= d42;                                                     
  d43 <= c42;                                                     
  c43 <= b42;
      b43 <= b42 + (((a42 + (b42 ^ c42 ^ d42) + 'hd4ef3085 + w42_3) << 16) | ((a42 + (b42 ^ c42 ^ d42) + 'hd4ef3085 + w42_3) >> (32 - 16)));
      w43_0 <= w42_0;         
  w43_1 <= w42_1;         
  w43_2 <= w42_2;         
  w43_3 <= w42_3;         
  w43_4 <= w42_4;         
  w43_5 <= w42_5;         
  w43_6 <= w42_6;         
  w43_7 <= w42_7;         
  w43_8 <= w42_8;         
  w43_9 <= w42_9;         
  w43_10 <= w42_10;       
  w43_11 <= w42_11;       
  w43_12 <= w42_12;       
  w43_13 <= w42_13;       
  w43_14 <= w42_14;       
  w43_15 <= w42_15;

      a44 <= d43;                                                     
  d44 <= c43;                                                     
  c44 <= b43;
      b44 <= b43 + (((a43 + (b43 ^ c43 ^ d43) + 'h04881d05 + w43_6) << 23) | ((a43 + (b43 ^ c43 ^ d43) + 'h04881d05 + w43_6) >> (32 - 23)));
      w44_0 <= w43_0;         
  w44_1 <= w43_1;         
  w44_2 <= w43_2;         
  w44_3 <= w43_3;         
  w44_4 <= w43_4;         
  w44_5 <= w43_5;         
  w44_6 <= w43_6;         
  w44_7 <= w43_7;         
  w44_8 <= w43_8;         
  w44_9 <= w43_9;         
  w44_10 <= w43_10;       
  w44_11 <= w43_11;       
  w44_12 <= w43_12;       
  w44_13 <= w43_13;       
  w44_14 <= w43_14;       
  w44_15 <= w43_15;

      a45 <= d44;                                                     
  d45 <= c44;                                                     
  c45 <= b44;
      b45 <= b44 + (((a44 + (b44 ^ c44 ^ d44) + 'hd9d4d039 + w44_9) << 4) | ((a44 + (b44 ^ c44 ^ d44) + 'hd9d4d039 + w44_9) >> (32 - 4)));
      w45_0 <= w44_0;         
  w45_1 <= w44_1;         
  w45_2 <= w44_2;         
  w45_3 <= w44_3;         
  w45_4 <= w44_4;         
  w45_5 <= w44_5;         
  w45_6 <= w44_6;         
  w45_7 <= w44_7;         
  w45_8 <= w44_8;         
  w45_9 <= w44_9;         
  w45_10 <= w44_10;       
  w45_11 <= w44_11;       
  w45_12 <= w44_12;       
  w45_13 <= w44_13;       
  w45_14 <= w44_14;       
  w45_15 <= w44_15;

      a46 <= d45;                                                     
  d46 <= c45;                                                     
  c46 <= b45;
      b46 <= b45 + (((a45 + (b45 ^ c45 ^ d45) + 'he6db99e5 + w45_12) << 11) | ((a45 + (b45 ^ c45 ^ d45) + 'he6db99e5 + w45_12) >> (32 - 11)));
      w46_0 <= w45_0;         
  w46_1 <= w45_1;         
  w46_2 <= w45_2;         
  w46_3 <= w45_3;         
  w46_4 <= w45_4;         
  w46_5 <= w45_5;         
  w46_6 <= w45_6;         
  w46_7 <= w45_7;         
  w46_8 <= w45_8;         
  w46_9 <= w45_9;         
  w46_10 <= w45_10;       
  w46_11 <= w45_11;       
  w46_12 <= w45_12;       
  w46_13 <= w45_13;       
  w46_14 <= w45_14;       
  w46_15 <= w45_15;

      a47 <= d46;                                                     
  d47 <= c46;                                                     
  c47 <= b46;
      b47 <= b46 + (((a46 + (b46 ^ c46 ^ d46) + 'h1fa27cf8 + w46_15) << 16) | ((a46 + (b46 ^ c46 ^ d46) + 'h1fa27cf8 + w46_15) >> (32 - 16)));
      w47_0 <= w46_0;         
  w47_1 <= w46_1;         
  w47_2 <= w46_2;         
  w47_3 <= w46_3;         
  w47_4 <= w46_4;         
  w47_5 <= w46_5;         
  w47_6 <= w46_6;         
  w47_7 <= w46_7;         
  w47_8 <= w46_8;         
  w47_9 <= w46_9;         
  w47_10 <= w46_10;       
  w47_11 <= w46_11;       
  w47_12 <= w46_12;       
  w47_13 <= w46_13;       
  w47_14 <= w46_14;       
  w47_15 <= w46_15;

      a48 <= d47;                                                     
  d48 <= c47;                                                     
  c48 <= b47;
      b48 <= b47 + (((a47 + (b47 ^ c47 ^ d47) + 'hc4ac5665 + w47_2) << 23) | ((a47 + (b47 ^ c47 ^ d47) + 'hc4ac5665 + w47_2) >> (32 - 23)));
      w48_0 <= w47_0;         
  w48_1 <= w47_1;         
  w48_2 <= w47_2;         
  w48_3 <= w47_3;         
  w48_4 <= w47_4;         
  w48_5 <= w47_5;         
  w48_6 <= w47_6;         
  w48_7 <= w47_7;         
  w48_8 <= w47_8;         
  w48_9 <= w47_9;         
  w48_10 <= w47_10;       
  w48_11 <= w47_11;       
  w48_12 <= w47_12;       
  w48_13 <= w47_13;       
  w48_14 <= w47_14;       
  w48_15 <= w47_15;

      a49 <= d48;                                                     
  d49 <= c48;                                                     
  c49 <= b48;
      b49 <= b48 + (((a48 + (c48 ^ (b48 | (~d48))) + 'hf4292244 + w48_0) << 6) | ((a48 + (c48 ^ (b48 | (~d48))) + 'hf4292244 + w48_0) >> (32 - 6)));
      w49_0 <= w48_0;         
  w49_1 <= w48_1;         
  w49_2 <= w48_2;         
  w49_3 <= w48_3;         
  w49_4 <= w48_4;         
  w49_5 <= w48_5;         
  w49_6 <= w48_6;         
  w49_7 <= w48_7;         
  w49_8 <= w48_8;         
  w49_9 <= w48_9;         
  w49_10 <= w48_10;       
  w49_11 <= w48_11;       
  w49_12 <= w48_12;       
  w49_13 <= w48_13;       
  w49_14 <= w48_14;       
  w49_15 <= w48_15;

      a50 <= d49;                                                     
  d50 <= c49;                                                     
  c50 <= b49;
      b50 <= b49 + (((a49 + (c49 ^ (b49 | (~d49))) + 'h432aff97 + w49_7) << 10) | ((a49 + (c49 ^ (b49 | (~d49))) + 'h432aff97 + w49_7) >> (32 - 10)));
      w50_0 <= w49_0;         
  w50_1 <= w49_1;         
  w50_2 <= w49_2;         
  w50_3 <= w49_3;         
  w50_4 <= w49_4;         
  w50_5 <= w49_5;         
  w50_6 <= w49_6;         
  w50_7 <= w49_7;         
  w50_8 <= w49_8;         
  w50_9 <= w49_9;         
  w50_10 <= w49_10;       
  w50_11 <= w49_11;       
  w50_12 <= w49_12;       
  w50_13 <= w49_13;       
  w50_14 <= w49_14;       
  w50_15 <= w49_15;

      a51 <= d50;                                                     
  d51 <= c50;                                                     
  c51 <= b50;
      b51 <= b50 + (((a50 + (c50 ^ (b50 | (~d50))) + 'hab9423a7 + w50_14) << 15) | ((a50 + (c50 ^ (b50 | (~d50))) + 'hab9423a7 + w50_14) >> (32 - 15)));
      w51_0 <= w50_0;         
  w51_1 <= w50_1;         
  w51_2 <= w50_2;         
  w51_3 <= w50_3;         
  w51_4 <= w50_4;         
  w51_5 <= w50_5;         
  w51_6 <= w50_6;         
  w51_7 <= w50_7;         
  w51_8 <= w50_8;         
  w51_9 <= w50_9;         
  w51_10 <= w50_10;       
  w51_11 <= w50_11;       
  w51_12 <= w50_12;       
  w51_13 <= w50_13;       
  w51_14 <= w50_14;       
  w51_15 <= w50_15;

      a52 <= d51;                                                     
  d52 <= c51;                                                     
  c52 <= b51;
      b52 <= b51 + (((a51 + (c51 ^ (b51 | (~d51))) + 'hfc93a039 + w51_5) << 21) | ((a51 + (c51 ^ (b51 | (~d51))) + 'hfc93a039 + w51_5) >> (32 - 21)));
      w52_0 <= w51_0;         
  w52_1 <= w51_1;         
  w52_2 <= w51_2;         
  w52_3 <= w51_3;         
  w52_4 <= w51_4;         
  w52_5 <= w51_5;         
  w52_6 <= w51_6;         
  w52_7 <= w51_7;         
  w52_8 <= w51_8;         
  w52_9 <= w51_9;         
  w52_10 <= w51_10;       
  w52_11 <= w51_11;       
  w52_12 <= w51_12;       
  w52_13 <= w51_13;       
  w52_14 <= w51_14;       
  w52_15 <= w51_15;

      a53 <= d52;                                                     
  d53 <= c52;                                                     
  c53 <= b52;
      b53 <= b52 + (((a52 + (c52 ^ (b52 | (~d52))) + 'h655b59c3 + w52_12) << 6) | ((a52 + (c52 ^ (b52 | (~d52))) + 'h655b59c3 + w52_12) >> (32 - 6)));
      w53_0 <= w52_0;         
  w53_1 <= w52_1;         
  w53_2 <= w52_2;         
  w53_3 <= w52_3;         
  w53_4 <= w52_4;         
  w53_5 <= w52_5;         
  w53_6 <= w52_6;         
  w53_7 <= w52_7;         
  w53_8 <= w52_8;         
  w53_9 <= w52_9;         
  w53_10 <= w52_10;       
  w53_11 <= w52_11;       
  w53_12 <= w52_12;       
  w53_13 <= w52_13;       
  w53_14 <= w52_14;       
  w53_15 <= w52_15;

      a54 <= d53;                                                     
  d54 <= c53;                                                     
  c54 <= b53;
      b54 <= b53 + (((a53 + (c53 ^ (b53 | (~d53))) + 'h8f0ccc92 + w53_3) << 10) | ((a53 + (c53 ^ (b53 | (~d53))) + 'h8f0ccc92 + w53_3) >> (32 - 10)));
      w54_0 <= w53_0;         
  w54_1 <= w53_1;         
  w54_2 <= w53_2;         
  w54_3 <= w53_3;         
  w54_4 <= w53_4;         
  w54_5 <= w53_5;         
  w54_6 <= w53_6;         
  w54_7 <= w53_7;         
  w54_8 <= w53_8;         
  w54_9 <= w53_9;         
  w54_10 <= w53_10;       
  w54_11 <= w53_11;       
  w54_12 <= w53_12;       
  w54_13 <= w53_13;       
  w54_14 <= w53_14;       
  w54_15 <= w53_15;

      a55 <= d54;                                                     
  d55 <= c54;                                                     
  c55 <= b54;
      b55 <= b54 + (((a54 + (c54 ^ (b54 | (~d54))) + 'hffeff47d + w54_10) << 15) | ((a54 + (c54 ^ (b54 | (~d54))) + 'hffeff47d + w54_10) >> (32 - 15)));
      w55_0 <= w54_0;         
  w55_1 <= w54_1;         
  w55_2 <= w54_2;         
  w55_3 <= w54_3;         
  w55_4 <= w54_4;         
  w55_5 <= w54_5;         
  w55_6 <= w54_6;         
  w55_7 <= w54_7;         
  w55_8 <= w54_8;         
  w55_9 <= w54_9;         
  w55_10 <= w54_10;       
  w55_11 <= w54_11;       
  w55_12 <= w54_12;       
  w55_13 <= w54_13;       
  w55_14 <= w54_14;       
  w55_15 <= w54_15;

      a56 <= d55;                                                     
  d56 <= c55;                                                     
  c56 <= b55;
      b56 <= b55 + (((a55 + (c55 ^ (b55 | (~d55))) + 'h85845dd1 + w55_1) << 21) | ((a55 + (c55 ^ (b55 | (~d55))) + 'h85845dd1 + w55_1) >> (32 - 21)));
      w56_0 <= w55_0;         
  w56_1 <= w55_1;         
  w56_2 <= w55_2;         
  w56_3 <= w55_3;         
  w56_4 <= w55_4;         
  w56_5 <= w55_5;         
  w56_6 <= w55_6;         
  w56_7 <= w55_7;         
  w56_8 <= w55_8;         
  w56_9 <= w55_9;         
  w56_10 <= w55_10;       
  w56_11 <= w55_11;       
  w56_12 <= w55_12;       
  w56_13 <= w55_13;       
  w56_14 <= w55_14;       
  w56_15 <= w55_15;

      a57 <= d56;                                                     
  d57 <= c56;                                                     
  c57 <= b56;
      b57 <= b56 + (((a56 + (c56 ^ (b56 | (~d56))) + 'h6fa87e4f + w56_8) << 6) | ((a56 + (c56 ^ (b56 | (~d56))) + 'h6fa87e4f + w56_8) >> (32 - 6)));
      w57_0 <= w56_0;         
  w57_1 <= w56_1;         
  w57_2 <= w56_2;         
  w57_3 <= w56_3;         
  w57_4 <= w56_4;         
  w57_5 <= w56_5;         
  w57_6 <= w56_6;         
  w57_7 <= w56_7;         
  w57_8 <= w56_8;         
  w57_9 <= w56_9;         
  w57_10 <= w56_10;       
  w57_11 <= w56_11;       
  w57_12 <= w56_12;       
  w57_13 <= w56_13;       
  w57_14 <= w56_14;       
  w57_15 <= w56_15;

      a58 <= d57;                                                     
  d58 <= c57;                                                     
  c58 <= b57;
      b58 <= b57 + (((a57 + (c57 ^ (b57 | (~d57))) + 'hfe2ce6e0 + w57_15) << 10) | ((a57 + (c57 ^ (b57 | (~d57))) + 'hfe2ce6e0 + w57_15) >> (32 - 10)));
      w58_0 <= w57_0;         
  w58_1 <= w57_1;         
  w58_2 <= w57_2;         
  w58_3 <= w57_3;         
  w58_4 <= w57_4;         
  w58_5 <= w57_5;         
  w58_6 <= w57_6;         
  w58_7 <= w57_7;         
  w58_8 <= w57_8;         
  w58_9 <= w57_9;         
  w58_10 <= w57_10;       
  w58_11 <= w57_11;       
  w58_12 <= w57_12;       
  w58_13 <= w57_13;       
  w58_14 <= w57_14;       
  w58_15 <= w57_15;

      a59 <= d58;                                                     
  d59 <= c58;                                                     
  c59 <= b58;
      b59 <= b58 + (((a58 + (c58 ^ (b58 | (~d58))) + 'ha3014314 + w58_6) << 15) | ((a58 + (c58 ^ (b58 | (~d58))) + 'ha3014314 + w58_6) >> (32 - 15)));
      w59_0 <= w58_0;         
  w59_1 <= w58_1;         
  w59_2 <= w58_2;         
  w59_3 <= w58_3;         
  w59_4 <= w58_4;         
  w59_5 <= w58_5;         
  w59_6 <= w58_6;         
  w59_7 <= w58_7;         
  w59_8 <= w58_8;         
  w59_9 <= w58_9;         
  w59_10 <= w58_10;       
  w59_11 <= w58_11;       
  w59_12 <= w58_12;       
  w59_13 <= w58_13;       
  w59_14 <= w58_14;       
  w59_15 <= w58_15;

      a60 <= d59;                                                     
  d60 <= c59;                                                     
  c60 <= b59;
      b60 <= b59 + (((a59 + (c59 ^ (b59 | (~d59))) + 'h4e0811a1 + w59_13) << 21) | ((a59 + (c59 ^ (b59 | (~d59))) + 'h4e0811a1 + w59_13) >> (32 - 21)));
      w60_0 <= w59_0;         
  w60_1 <= w59_1;         
  w60_2 <= w59_2;         
  w60_3 <= w59_3;         
  w60_4 <= w59_4;         
  w60_5 <= w59_5;         
  w60_6 <= w59_6;         
  w60_7 <= w59_7;         
  w60_8 <= w59_8;         
  w60_9 <= w59_9;         
  w60_10 <= w59_10;       
  w60_11 <= w59_11;       
  w60_12 <= w59_12;       
  w60_13 <= w59_13;       
  w60_14 <= w59_14;       
  w60_15 <= w59_15;

      a61 <= d60;                                                     
  d61 <= c60;                                                     
  c61 <= b60;
      b61 <= b60 + (((a60 + (c60 ^ (b60 | (~d60))) + 'hf7537e82 + w60_4) << 6) | ((a60 + (c60 ^ (b60 | (~d60))) + 'hf7537e82 + w60_4) >> (32 - 6)));
      w61_0 <= w60_0;         
  w61_1 <= w60_1;         
  w61_2 <= w60_2;         
  w61_3 <= w60_3;         
  w61_4 <= w60_4;         
  w61_5 <= w60_5;         
  w61_6 <= w60_6;         
  w61_7 <= w60_7;         
  w61_8 <= w60_8;         
  w61_9 <= w60_9;         
  w61_10 <= w60_10;       
  w61_11 <= w60_11;       
  w61_12 <= w60_12;       
  w61_13 <= w60_13;       
  w61_14 <= w60_14;       
  w61_15 <= w60_15;

      a62 <= d61;                                                     
  d62 <= c61;                                                     
  c62 <= b61;
      b62 <= b61 + (((a61 + (c61 ^ (b61 | (~d61))) + 'hbd3af235 + w61_11) << 10) | ((a61 + (c61 ^ (b61 | (~d61))) + 'hbd3af235 + w61_11) >> (32 - 10)));
      w62_0 <= w61_0;         
  w62_1 <= w61_1;         
  w62_2 <= w61_2;         
  w62_3 <= w61_3;         
  w62_4 <= w61_4;         
  w62_5 <= w61_5;         
  w62_6 <= w61_6;         
  w62_7 <= w61_7;         
  w62_8 <= w61_8;         
  w62_9 <= w61_9;         
  w62_10 <= w61_10;       
  w62_11 <= w61_11;       
  w62_12 <= w61_12;       
  w62_13 <= w61_13;       
  w62_14 <= w61_14;       
  w62_15 <= w61_15;

      a63 <= d62;                                                     
  d63 <= c62;                                                     
  c63 <= b62;
      b63 <= b62 + (((a62 + (c62 ^ (b62 | (~d62))) + 'h2ad7d2bb + w62_2) << 15) | ((a62 + (c62 ^ (b62 | (~d62))) + 'h2ad7d2bb + w62_2) >> (32 - 15)));
      w63_0 <= w62_0;         
  w63_1 <= w62_1;         
  w63_2 <= w62_2;         
  w63_3 <= w62_3;         
  w63_4 <= w62_4;         
  w63_5 <= w62_5;         
  w63_6 <= w62_6;         
  w63_7 <= w62_7;         
  w63_8 <= w62_8;         
  w63_9 <= w62_9;         
  w63_10 <= w62_10;       
  w63_11 <= w62_11;       
  w63_12 <= w62_12;       
  w63_13 <= w62_13;       
  w63_14 <= w62_14;       
  w63_15 <= w62_15;

      a64 <= d63;                                                     
  d64 <= c63;                                                     
  c64 <= b63;
      b64 <= b63 + (((a63 + (c63 ^ (b63 | (~d63))) + 'heb86d391 + w63_9) << 21) | ((a63 + (c63 ^ (b63 | (~d63))) + 'heb86d391 + w63_9) >> (32 - 21)));
    end
endmodule
