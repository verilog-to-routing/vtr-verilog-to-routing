/*
 * Wide range test
*/

`define WIDTH 3
`define operator nor
`include "replicate_any_width_binary_test.v"