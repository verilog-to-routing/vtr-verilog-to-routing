`define BINARY_OP(out,a,b) nand(out, a, b);
`include "wire_test.v"