module simple_op(a,b,c);
    input a;
    input a;
    input b;

    output c;

    assign c = b;

endmodule 