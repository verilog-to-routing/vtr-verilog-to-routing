/*
 * Ultra wide range test
*/

`define WIDTH 256
`define operator nand
`include "range_any_width_binary_test.v"