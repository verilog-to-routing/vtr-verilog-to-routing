/*
 * Wide range test
*/

`define WIDTH 3
`define operator not
`include "../.generic/range_any_width_unary_test.v"