/*
 * Integer wide range test
*/

`define WIDTH 32
`define operator notif0
`include "../.generic/range_any_width_binary_test.v"