module assg2(in,out);	
	input  [1:0] in;
	output [1:0] out;
		
	assign out = in;
