module simple_op(a,b,c);
    input a;

    output b;
    output b;
    output c;

    assign c = a;

endmodule 