/*
 * Integer wide range test
*/

`define WIDTH 32
`define operator and
`include "range_any_width_binary_test.v"