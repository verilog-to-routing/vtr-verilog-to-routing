`define UNARY_OP(out,a) not(out, a);
`include "wire_test.v"