
`timescale 1ns/10ps

module timescale_syntax (a,b,c);

input a;
input b;
output c;

assign c = a ^ b;

endmodule