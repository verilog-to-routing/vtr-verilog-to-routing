// Content from two_kmeans.v

module top (
    input  wire                        clk,
    input  wire                        rst,

    /*
     * AXI slave interface
     */
    input  wire [7:0]                  s_axi_awid,
    input  wire [7:0]                  s_axi_awaddr,
    input  wire [7:0]                  s_axi_awlen,
    input  wire [2:0]                  s_axi_awsize,
    input  wire [1:0]                  s_axi_awburst,
    input  wire                        s_axi_awlock,
    input  wire [3:0]                  s_axi_awcache,
    input  wire [2:0]                  s_axi_awprot,
    input  wire                        s_axi_awvalid,
    output wire                        s_axi_awready,
    input  wire [31:0]   s_axi_wdata,
    input  wire [3:0]   s_axi_wstrb,
    input  wire                        s_axi_wlast,
    input  wire                        s_axi_wvalid,
    output wire                        s_axi_wready,
    output wire [7:0]     s_axi_bid,
    output wire [1:0]                  s_axi_bresp,
    output wire                        s_axi_bvalid,
    input  wire                        s_axi_bready,
    input  wire [7:0]     s_axi_arid,
    input  wire [7:0]       s_axi_araddr,
    input  wire [7:0]                  s_axi_arlen,
    input  wire [2:0]                  s_axi_arsize,
    input  wire [1:0]                  s_axi_arburst,
    input  wire                        s_axi_arlock,
    input  wire [3:0]                  s_axi_arcache,
    input  wire [2:0]                  s_axi_arprot,
    input  wire                        s_axi_arvalid,
    output wire                        s_axi_arready,
    output wire [7:0]     s_axi_rid,
    output wire [31:0]   s_axi_rdata,
    output wire [1:0]                  s_axi_rresp,
    output wire                        s_axi_rlast,
    output wire                        s_axi_rvalid,
    input  wire                        s_axi_rready,


    /*
     * AXI master interface
     */
    output wire [7:0]      m00_axi_awid,
    output wire [63:0]    m00_axi_awaddr,
    output wire [7:0]               m00_axi_awlen,
    output wire [2:0]               m00_axi_awsize,
    output wire [1:0]               m00_axi_awburst,
    output wire                     m00_axi_awlock,
    output wire [3:0]               m00_axi_awcache,
    output wire [2:0]               m00_axi_awprot,
    output wire [3:0]               m00_axi_awqos,
    output wire [3:0]               m00_axi_awregion,
    output wire [0:0]  m00_axi_awuser,
    output wire                     m00_axi_awvalid,
    input  wire                     m00_axi_awready,
    output wire [63:0]    m00_axi_wdata,
    output wire [7:0]    m00_axi_wstrb,
    output wire                     m00_axi_wlast,
    output wire [0:0]   m00_axi_wuser,
    output wire                     m00_axi_wvalid,
    input  wire                     m00_axi_wready,
    input  wire [7:0]      m00_axi_bid,
    input  wire [1:0]               m00_axi_bresp,
    input  wire [0:0]   m00_axi_buser,
    input  wire                     m00_axi_bvalid,
    output wire                     m00_axi_bready,
    output wire [7:0]      m00_axi_arid,
    output wire [63:0]    m00_axi_araddr,
    output wire [7:0]               m00_axi_arlen,
    output wire [2:0]               m00_axi_arsize,
    output wire [1:0]               m00_axi_arburst,
    output wire                     m00_axi_arlock,
    output wire [3:0]               m00_axi_arcache,
    output wire [2:0]               m00_axi_arprot,
    output wire [3:0]               m00_axi_arqos,
    output wire [3:0]               m00_axi_arregion,
    output wire [0:0]  m00_axi_aruser,
    output wire                     m00_axi_arvalid,
    input  wire                     m00_axi_arready,
    input  wire [7:0]      m00_axi_rid,
    input  wire [63:0]    m00_axi_rdata,
    input  wire [1:0]               m00_axi_rresp,
    input  wire                     m00_axi_rlast,
    input  wire [0:0]   m00_axi_ruser,
    input  wire                     m00_axi_rvalid,
    output wire                     m00_axi_rready

);

    wire ap_clk;
    wire ap_rst_n;

    assign ap_clk = clk;
    assign ap_rst_n = ~rst;
    
    wire axi0_mem_AWVALID;
    wire axi0_mem_AWREADY;
    wire [63:0] axi0_mem_AWADDR;
    wire [0:0] axi0_mem_AWID;
    wire [7:0] axi0_mem_AWLEN;
    wire [2:0] axi0_mem_AWSIZE;
    wire [1:0] axi0_mem_AWBURST;
    wire [1:0] axi0_mem_AWLOCK;
    wire [3:0] axi0_mem_AWCACHE;
    wire [2:0] axi0_mem_AWPROT;
    wire [3:0] axi0_mem_AWQOS;
    wire [3:0] axi0_mem_AWREGION;
    wire [0:0] axi0_mem_AWUSER;
    
    wire axi0_mem_WVALID;
    wire axi0_mem_WREADY;
    wire [63:0] axi0_mem_WDATA;
    wire [7:0] axi0_mem_WSTRB;
    wire axi0_mem_WLAST;
    wire [0:0] axi0_mem_WID;
    wire [0:0] axi0_mem_WUSER;
    
    wire axi0_mem_ARVALID;
    wire axi0_mem_ARREADY;
    wire [63:0] axi0_mem_ARADDR;
    wire [0:0] axi0_mem_ARID;
    wire [7:0] axi0_mem_ARLEN;
    wire [2:0] axi0_mem_ARSIZE;
    wire [1:0] axi0_mem_ARBURST;
    wire [1:0] axi0_mem_ARLOCK;
    wire [3:0] axi0_mem_ARCACHE;
    wire [2:0] axi0_mem_ARPROT;
    wire [3:0] axi0_mem_ARQOS;
    wire [3:0] axi0_mem_ARREGION;
    wire [0:0] axi0_mem_ARUSER;
    
    wire axi0_mem_RVALID;
    wire axi0_mem_RREADY;
    wire [63:0] axi0_mem_RDATA;
    wire axi0_mem_RLAST;
    wire [0:0] axi0_mem_RID;
    wire [0:0] axi0_mem_RUSER;
    wire [1:0] axi0_mem_RRESP;
    
    wire axi0_mem_BVALID;
    wire axi0_mem_BREADY;
    wire [1:0] axi0_mem_BRESP;
    wire [0:0] axi0_mem_BID;
    wire [0:0] axi0_mem_BUSER;
    
    wire axi0_cfg_AWVALID;
    wire axi0_cfg_AWREADY;
    wire [7:0] axi0_cfg_AWADDR;
    wire axi0_cfg_WVALID;
    wire axi0_cfg_WREADY;
    wire [31:0] axi0_cfg_WDATA;
    wire [3:0] axi0_cfg_WSTRB;
    wire axi0_cfg_ARVALID;
    wire axi0_cfg_ARREADY;
    wire [7:0] axi0_cfg_ARADDR;
    
    wire axi0_cfg_RVALID;
    wire axi0_cfg_RREADY;
    wire [31:0] axi0_cfg_RDATA;
    wire [1:0] axi0_cfg_RRESP;
    
    wire axi0_cfg_BVALID;
    wire axi0_cfg_BREADY;
    wire [1:0] axi0_cfg_BRESP;
    wire interrupt0;

    wire axi1_mem_AWVALID;
    wire axi1_mem_AWREADY;
    wire [63:0] axi1_mem_AWADDR;
    wire [0:0] axi1_mem_AWID;
    wire [7:0] axi1_mem_AWLEN;
    wire [2:0] axi1_mem_AWSIZE;
    wire [1:0] axi1_mem_AWBURST;
    wire [1:0] axi1_mem_AWLOCK;
    wire [3:0] axi1_mem_AWCACHE;
    wire [2:0] axi1_mem_AWPROT;
    wire [3:0] axi1_mem_AWQOS;
    wire [3:0] axi1_mem_AWREGION;
    wire [0:0] axi1_mem_AWUSER;

    wire axi1_mem_WVALID;
    wire axi1_mem_WREADY;
    wire [63:0] axi1_mem_WDATA;
    wire [7:0] axi1_mem_WSTRB;
    wire axi1_mem_WLAST;
    wire [0:0] axi1_mem_WID;
    wire [0:0] axi1_mem_WUSER;

    wire axi1_mem_ARVALID;
    wire axi1_mem_ARREADY;
    wire [63:0] axi1_mem_ARADDR;
    wire [0:0] axi1_mem_ARID;
    wire [7:0] axi1_mem_ARLEN;
    wire [2:0] axi1_mem_ARSIZE;
    wire [1:0] axi1_mem_ARBURST;
    wire [1:0] axi1_mem_ARLOCK;
    wire [3:0] axi1_mem_ARCACHE;
    wire [2:0] axi1_mem_ARPROT;
    wire [3:0] axi1_mem_ARQOS;
    wire [3:0] axi1_mem_ARREGION;
    wire [0:0] axi1_mem_ARUSER;

    wire axi1_mem_RVALID;
    wire axi1_mem_RREADY;
    wire [63:0] axi1_mem_RDATA;
    wire axi1_mem_RLAST;
    wire [0:0] axi1_mem_RID;
    wire [0:0] axi1_mem_RUSER;
    wire [1:0] axi1_mem_RRESP;

    wire axi1_mem_BVALID;
    wire axi1_mem_BREADY;
    wire [1:0] axi1_mem_BRESP;
    wire [0:0] axi1_mem_BID;
    wire [0:0] axi1_mem_BUSER;

    wire axi1_cfg_AWVALID;
    wire axi1_cfg_AWREADY;
    wire [7:0] axi1_cfg_AWADDR;
    wire axi1_cfg_WVALID;
    wire axi1_cfg_WREADY;
    wire [31:0] axi1_cfg_WDATA;
    wire [3:0] axi1_cfg_WSTRB;
    wire axi1_cfg_ARVALID;
    wire axi1_cfg_ARREADY;
    wire [7:0] axi1_cfg_ARADDR;

    wire axi1_cfg_RVALID;
    wire axi1_cfg_RREADY;
    wire [31:0] axi1_cfg_RDATA;
    wire [1:0] axi1_cfg_RRESP;

    wire axi1_cfg_BVALID;
    wire axi1_cfg_BREADY;
    wire [1:0] axi1_cfg_BRESP;
    wire interrupt1;

    wire axi_shared_cfg_AWVALID;
    wire axi_shared_cfg_AWREADY;
    wire [7:0] axi_shared_cfg_AWADDR;
    wire axi_shared_cfg_WVALID;
    wire axi_shared_cfg_WREADY;
    wire [31:0] axi_shared_cfg_WDATA;
    wire [3:0] axi_shared_cfg_WSTRB;
    wire axi_shared_cfg_ARVALID;
    wire axi_shared_cfg_ARREADY;
    wire [7:0] axi_shared_cfg_ARADDR;
    wire axi_shared_cfg_RVALID;
    wire axi_shared_cfg_RREADY;
    wire [31:0] axi_shared_cfg_RDATA;
    wire [1:0] axi_shared_cfg_RRESP;
    wire axi_shared_cfg_BVALID;
    wire axi_shared_cfg_BREADY;
    wire [1:0] axi_shared_cfg_BRESP;
    
    kmeans_flat kmeans_inst0 (
        .ap_clk(ap_clk),
        .ap_rst_n(ap_rst_n),

        .m_axi_mem_AWVALID(axi0_mem_AWVALID),
        .m_axi_mem_AWREADY(axi0_mem_AWREADY),
        .m_axi_mem_AWADDR(axi0_mem_AWADDR),
        .m_axi_mem_AWID(axi0_mem_AWID),
        .m_axi_mem_AWLEN(axi0_mem_AWLEN),
        .m_axi_mem_AWSIZE(axi0_mem_AWSIZE),
        .m_axi_mem_AWBURST(axi0_mem_AWBURST),
        .m_axi_mem_AWLOCK(axi0_mem_AWLOCK),
        .m_axi_mem_AWCACHE(axi0_mem_AWCACHE),
        .m_axi_mem_AWPROT(axi0_mem_AWPROT),
        .m_axi_mem_AWQOS(axi0_mem_AWQOS),
        .m_axi_mem_AWREGION(axi0_mem_AWREGION),
        .m_axi_mem_AWUSER(axi0_mem_AWUSER),
        .m_axi_mem_WVALID(axi0_mem_WVALID),
        .m_axi_mem_WREADY(axi0_mem_WREADY),
        .m_axi_mem_WDATA(axi0_mem_WDATA),
        .m_axi_mem_WSTRB(axi0_mem_WSTRB),
        .m_axi_mem_WLAST(axi0_mem_WLAST),
        .m_axi_mem_WID(axi0_mem_WID),
        .m_axi_mem_WUSER(axi0_mem_WUSER),
        .m_axi_mem_ARVALID(axi0_mem_ARVALID),
        .m_axi_mem_ARREADY(axi0_mem_ARREADY),
        .m_axi_mem_ARADDR(axi0_mem_ARADDR),
        .m_axi_mem_ARID(axi0_mem_ARID),
        .m_axi_mem_ARLEN(axi0_mem_ARLEN),
        .m_axi_mem_ARSIZE(axi0_mem_ARSIZE),
        .m_axi_mem_ARBURST(axi0_mem_ARBURST),
        .m_axi_mem_ARLOCK(axi0_mem_ARLOCK),
        .m_axi_mem_ARCACHE(axi0_mem_ARCACHE),
        .m_axi_mem_ARPROT(axi0_mem_ARPROT),
        .m_axi_mem_ARQOS(axi0_mem_ARQOS),
        .m_axi_mem_ARREGION(axi0_mem_ARREGION),
        .m_axi_mem_ARUSER(axi0_mem_ARUSER),
        .m_axi_mem_RVALID(axi0_mem_RVALID),
        .m_axi_mem_RREADY(axi0_mem_RREADY),
        .m_axi_mem_RDATA(axi0_mem_RDATA),
        .m_axi_mem_RLAST(axi0_mem_RLAST),
        .m_axi_mem_RID(axi0_mem_RID),
        .m_axi_mem_RUSER(axi0_mem_RUSER),
        .m_axi_mem_RRESP(axi0_mem_RRESP),
        .m_axi_mem_BVALID(axi0_mem_BVALID),
        .m_axi_mem_BREADY(axi0_mem_BREADY),
        .m_axi_mem_BRESP(axi0_mem_BRESP),
        .m_axi_mem_BID(axi0_mem_BID),
        .m_axi_mem_BUSER(axi0_mem_BUSER),

        .s_axi_cfg_AWVALID(axi0_cfg_AWVALID),
        .s_axi_cfg_AWREADY(axi0_cfg_AWREADY),
        .s_axi_cfg_AWADDR(axi0_cfg_AWADDR),
        .s_axi_cfg_WVALID(axi0_cfg_WVALID),
        .s_axi_cfg_WREADY(axi0_cfg_WREADY),
        .s_axi_cfg_WDATA(axi0_cfg_WDATA),
        .s_axi_cfg_WSTRB(axi0_cfg_WSTRB),
        .s_axi_cfg_ARVALID(axi0_cfg_ARVALID),
        .s_axi_cfg_ARREADY(axi0_cfg_ARREADY),
        .s_axi_cfg_ARADDR(axi0_cfg_ARADDR),
        .s_axi_cfg_RVALID(axi0_cfg_RVALID),
        .s_axi_cfg_RREADY(axi0_cfg_RREADY),
        .s_axi_cfg_RDATA(axi0_cfg_RDATA),
        .s_axi_cfg_RRESP(axi0_cfg_RRESP),
        .s_axi_cfg_BVALID(axi0_cfg_BVALID),
        .s_axi_cfg_BREADY(axi0_cfg_BREADY),
        .s_axi_cfg_BRESP(axi0_cfg_BRESP),
        .interrupt(interrupt0)
    );

    kmeans_flat kmeans_inst1 (
        .ap_clk(ap_clk),
        .ap_rst_n(ap_rst_n),
        .m_axi_mem_AWVALID(axi1_mem_AWVALID),
        .m_axi_mem_AWREADY(axi1_mem_AWREADY),
        .m_axi_mem_AWADDR(axi1_mem_AWADDR),
        .m_axi_mem_AWID(axi1_mem_AWID),
        .m_axi_mem_AWLEN(axi1_mem_AWLEN),
        .m_axi_mem_AWSIZE(axi1_mem_AWSIZE),
        .m_axi_mem_AWBURST(axi1_mem_AWBURST),
        .m_axi_mem_AWLOCK(axi1_mem_AWLOCK),
        .m_axi_mem_AWCACHE(axi1_mem_AWCACHE),
        .m_axi_mem_AWPROT(axi1_mem_AWPROT),
        .m_axi_mem_AWQOS(axi1_mem_AWQOS),
        .m_axi_mem_AWREGION(axi1_mem_AWREGION),
        .m_axi_mem_AWUSER(axi1_mem_AWUSER),
        .m_axi_mem_WVALID(axi1_mem_WVALID),
        .m_axi_mem_WREADY(axi1_mem_WREADY),
        .m_axi_mem_WDATA(axi1_mem_WDATA),
        .m_axi_mem_WSTRB(axi1_mem_WSTRB),
        .m_axi_mem_WLAST(axi1_mem_WLAST),
        .m_axi_mem_WID(axi1_mem_WID),
        .m_axi_mem_WUSER(axi1_mem_WUSER),
        .m_axi_mem_ARVALID(axi1_mem_ARVALID),
        .m_axi_mem_ARREADY(axi1_mem_ARREADY),
        .m_axi_mem_ARADDR(axi1_mem_ARADDR),
        .m_axi_mem_ARID(axi1_mem_ARID),
        .m_axi_mem_ARLEN(axi1_mem_ARLEN),
        .m_axi_mem_ARSIZE(axi1_mem_ARSIZE),
        .m_axi_mem_ARBURST(axi1_mem_ARBURST),
        .m_axi_mem_ARLOCK(axi1_mem_ARLOCK),
        .m_axi_mem_ARCACHE(axi1_mem_ARCACHE),
        .m_axi_mem_ARPROT(axi1_mem_ARPROT),
        .m_axi_mem_ARQOS(axi1_mem_ARQOS),
        .m_axi_mem_ARREGION(axi1_mem_ARREGION),
        .m_axi_mem_ARUSER(axi1_mem_ARUSER),
        .m_axi_mem_RVALID(axi1_mem_RVALID),
        .m_axi_mem_RREADY(axi1_mem_RREADY),
        .m_axi_mem_RDATA(axi1_mem_RDATA),
        .m_axi_mem_RLAST(axi1_mem_RLAST),
        .m_axi_mem_RID(axi1_mem_RID),
        .m_axi_mem_RUSER(axi1_mem_RUSER),
        .m_axi_mem_RRESP(axi1_mem_RRESP),
        .m_axi_mem_BVALID(axi1_mem_BVALID),
        .m_axi_mem_BREADY(axi1_mem_BREADY),
        .m_axi_mem_BRESP(axi1_mem_BRESP),
        .m_axi_mem_BID(axi1_mem_BID),
        .m_axi_mem_BUSER(axi1_mem_BUSER),
        .s_axi_cfg_AWVALID(axi1_cfg_AWVALID),
        .s_axi_cfg_AWREADY(axi1_cfg_AWREADY),
        .s_axi_cfg_AWADDR(axi1_cfg_AWADDR),
        .s_axi_cfg_WVALID(axi1_cfg_WVALID),
        .s_axi_cfg_WREADY(axi1_cfg_WREADY),
        .s_axi_cfg_WDATA(axi1_cfg_WDATA),
        .s_axi_cfg_WSTRB(axi1_cfg_WSTRB),
        .s_axi_cfg_ARVALID(axi1_cfg_ARVALID),
        .s_axi_cfg_ARREADY(axi1_cfg_ARREADY),
        .s_axi_cfg_ARADDR(axi1_cfg_ARADDR),
        .s_axi_cfg_RVALID(axi1_cfg_RVALID),
        .s_axi_cfg_RREADY(axi1_cfg_RREADY),
        .s_axi_cfg_RDATA(axi1_cfg_RDATA),
        .s_axi_cfg_RRESP(axi1_cfg_RRESP),
        .s_axi_cfg_BVALID(axi1_cfg_BVALID),
        .s_axi_cfg_BREADY(axi1_cfg_BREADY),
        .s_axi_cfg_BRESP(axi1_cfg_BRESP),
        .interrupt(interrupt1)
    );

    axi_interconnect_wrap_2x1 #(
        .DATA_WIDTH(64),
        .ADDR_WIDTH(64),
        .STRB_WIDTH(8), // DATA_WIDTH / 8
        .ID_WIDTH(8),
        .AWUSER_ENABLE(1),
        .AWUSER_WIDTH(1),
        .WUSER_ENABLE(1),
        .WUSER_WIDTH(1),
        .BUSER_ENABLE(1),
        .BUSER_WIDTH(1),
        .ARUSER_ENABLE(1),
        .ARUSER_WIDTH(1),
        .RUSER_ENABLE(1),
        .RUSER_WIDTH(1),
        .FORWARD_ID(1),
        .M_REGIONS(1),
        .M00_BASE_ADDR(0),
        .M00_ADDR_WIDTH({1{32'd64}}), // Single region, 24-bit width
        .M00_CONNECT_READ(2'b11),
        .M00_CONNECT_WRITE(2'b11),
        .M00_SECURE(1'b0)
    ) axi_interconnect_inst (
        .clk(ap_clk),
        .rst(~ap_rst_n),

        // Slave 0 Interface
        .s00_axi_awid(axi0_mem_AWID),
        .s00_axi_awaddr(axi0_mem_AWADDR),
        .s00_axi_awlen(axi0_mem_AWLEN),
        .s00_axi_awsize(axi0_mem_AWSIZE),
        .s00_axi_awburst(axi0_mem_AWBURST),
        .s00_axi_awlock(axi0_mem_AWLOCK),
        .s00_axi_awcache(axi0_mem_AWCACHE),
        .s00_axi_awprot(axi0_mem_AWPROT),
        .s00_axi_awqos(axi0_mem_AWQOS),
        .s00_axi_awuser(axi0_mem_AWUSER),
        .s00_axi_awvalid(axi0_mem_AWVALID),
        .s00_axi_awready(axi0_mem_AWREADY),

        .s00_axi_wdata(axi0_mem_WDATA),
        .s00_axi_wstrb(axi0_mem_WSTRB),
        .s00_axi_wlast(axi0_mem_WLAST),
        .s00_axi_wuser(axi0_mem_WUSER),
        .s00_axi_wvalid(axi0_mem_WVALID),
        .s00_axi_wready(axi0_mem_WREADY),

        .s00_axi_bid(axi0_mem_BID),
        .s00_axi_bresp(axi0_mem_BRESP),
        .s00_axi_buser(axi0_mem_BUSER),
        .s00_axi_bvalid(axi0_mem_BVALID),
        .s00_axi_bready(axi0_mem_BREADY),

        .s00_axi_arid(axi0_mem_ARID),
        .s00_axi_araddr(axi0_mem_ARADDR),
        .s00_axi_arlen(axi0_mem_ARLEN),
        .s00_axi_arsize(axi0_mem_ARSIZE),
        .s00_axi_arburst(axi0_mem_ARBURST),
        .s00_axi_arlock(axi0_mem_ARLOCK),
        .s00_axi_arcache(axi0_mem_ARCACHE),
        .s00_axi_arprot(axi0_mem_ARPROT),
        .s00_axi_arqos(axi0_mem_ARQOS),
        .s00_axi_aruser(axi0_mem_ARUSER),
        .s00_axi_arvalid(axi0_mem_ARVALID),
        .s00_axi_arready(axi0_mem_ARREADY),

        .s00_axi_rid(axi0_mem_RID),
        .s00_axi_rdata(axi0_mem_RDATA),
        .s00_axi_rresp(axi0_mem_RRESP),
        .s00_axi_rlast(axi0_mem_RLAST),
        .s00_axi_ruser(axi0_mem_RUSER),
        .s00_axi_rvalid(axi0_mem_RVALID),
        .s00_axi_rready(axi0_mem_RREADY),

        // Slave 1 Interface
        .s01_axi_awid(axi1_mem_AWID),
        .s01_axi_awaddr(axi1_mem_AWADDR),
        .s01_axi_awlen(axi1_mem_AWLEN),
        .s01_axi_awsize(axi1_mem_AWSIZE),
        .s01_axi_awburst(axi1_mem_AWBURST),
        .s01_axi_awlock(axi1_mem_AWLOCK),
        .s01_axi_awcache(axi1_mem_AWCACHE),
        .s01_axi_awprot(axi1_mem_AWPROT),
        .s01_axi_awqos(axi1_mem_AWQOS),
        .s01_axi_awuser(axi1_mem_AWUSER),
        .s01_axi_awvalid(axi1_mem_AWVALID),
        .s01_axi_awready(axi1_mem_AWREADY),

        .s01_axi_wdata(axi1_mem_WDATA),
        .s01_axi_wstrb(axi1_mem_WSTRB),
        .s01_axi_wlast(axi1_mem_WLAST),
        .s01_axi_wuser(axi1_mem_WUSER),
        .s01_axi_wvalid(axi1_mem_WVALID),
        .s01_axi_wready(axi1_mem_WREADY),

        .s01_axi_bid(axi1_mem_BID),
        .s01_axi_bresp(axi1_mem_BRESP),
        .s01_axi_buser(axi1_mem_BUSER),
        .s01_axi_bvalid(axi1_mem_BVALID),
        .s01_axi_bready(axi1_mem_BREADY),

        .s01_axi_arid(axi1_mem_ARID),
        .s01_axi_araddr(axi1_mem_ARADDR),
        .s01_axi_arlen(axi1_mem_ARLEN),
        .s01_axi_arsize(axi1_mem_ARSIZE),
        .s01_axi_arburst(axi1_mem_ARBURST),
        .s01_axi_arlock(axi1_mem_ARLOCK),
        .s01_axi_arcache(axi1_mem_ARCACHE),
        .s01_axi_arprot(axi1_mem_ARPROT),
        .s01_axi_arqos(axi1_mem_ARQOS),
        .s01_axi_aruser(axi1_mem_ARUSER),
        .s01_axi_arvalid(axi1_mem_ARVALID),
        .s01_axi_arready(axi1_mem_ARREADY),

        .s01_axi_rid(axi1_mem_RID),
        .s01_axi_rdata(axi1_mem_RDATA),
        .s01_axi_rresp(axi1_mem_RRESP),
        .s01_axi_rlast(axi1_mem_RLAST),
        .s01_axi_ruser(axi1_mem_RUSER),
        .s01_axi_rvalid(axi1_mem_RVALID),
        .s01_axi_rready(axi1_mem_RREADY),

        // Master 0 Interface
        .m00_axi_awid(m00_axi_awid),
        .m00_axi_awaddr(m00_axi_awaddr),
        .m00_axi_awlen(m00_axi_awlen),
        .m00_axi_awsize(m00_axi_awsize),
        .m00_axi_awburst(m00_axi_awburst),
        .m00_axi_awlock(m00_axi_awlock),
        .m00_axi_awcache(m00_axi_awcache),
        .m00_axi_awprot(m00_axi_awprot),
        .m00_axi_awqos(m00_axi_awqos),
        .m00_axi_awregion(m00_axi_awregion),
        .m00_axi_awuser(m00_axi_awuser),
        .m00_axi_awvalid(m00_axi_awvalid),
        .m00_axi_awready(m00_axi_awready),
        .m00_axi_wdata(m00_axi_wdata),
        .m00_axi_wstrb(m00_axi_wstrb),
        .m00_axi_wlast(m00_axi_wlast),
        .m00_axi_wuser(m00_axi_wuser),
        .m00_axi_wvalid(m00_axi_wvalid),
        .m00_axi_wready(m00_axi_wready),
        .m00_axi_bid(m00_axi_bid),
        .m00_axi_bresp(m00_axi_bresp),
        .m00_axi_buser(m00_axi_buser),
        .m00_axi_bvalid(m00_axi_bvalid),
        .m00_axi_bready(m00_axi_bready),
        .m00_axi_arid(m00_axi_arid),
        .m00_axi_araddr(m00_axi_araddr),
        .m00_axi_arlen(m00_axi_arlen),
        .m00_axi_arsize(m00_axi_arsize),
        .m00_axi_arburst(m00_axi_arburst),
        .m00_axi_arlock(m00_axi_arlock),
        .m00_axi_arcache(m00_axi_arcache),
        .m00_axi_arprot(m00_axi_arprot),
        .m00_axi_arqos(m00_axi_arqos),
        .m00_axi_arregion(m00_axi_arregion),
        .m00_axi_aruser(m00_axi_aruser),
        .m00_axi_arvalid(m00_axi_arvalid),
        .m00_axi_arready(m00_axi_arready),
        .m00_axi_rid(m00_axi_rid),
        .m00_axi_rdata(m00_axi_rdata),
        .m00_axi_rresp(m00_axi_rresp),
        .m00_axi_rlast(m00_axi_rlast),
        .m00_axi_ruser(m00_axi_ruser),
        .m00_axi_rvalid(m00_axi_rvalid),
        .m00_axi_rready(m00_axi_rready)
    );


    axil_interconnect_wrap_1x2 #(
        .DATA_WIDTH(32),
        .ADDR_WIDTH(8),
        .STRB_WIDTH(4), // DATA_WIDTH / 8
        .M_REGIONS(1),
        .M00_BASE_ADDR(8'h00), // Base address for Master 0
        .M00_ADDR_WIDTH({32'd24}), // Address width for Master 0
        .M00_CONNECT_READ(1'b1),  // Enable read connections for Master 0
        .M00_CONNECT_WRITE(1'b1), // Enable write connections for Master 0
        .M00_SECURE(1'b0),        // Security setting for Master 0
        .M01_BASE_ADDR(8'h80),    // Base address for Master 1
        .M01_ADDR_WIDTH({32'd24}), // Address width for Master 1
        .M01_CONNECT_READ(1'b1),  // Enable read connections for Master 1
        .M01_CONNECT_WRITE(1'b1), // Enable write connections for Master 1
        .M01_SECURE(1'b0)         // Security setting for Master 1
    ) axil_interconnect_inst (
        .clk(ap_clk),
        .rst(~ap_rst_n),

        // AXI-Lite Slave Interface
        .s00_axil_awaddr(axi_shared_cfg_AWADDR),
        .s00_axil_awprot(0),
        .s00_axil_awvalid(axi_shared_cfg_AWVALID),
        .s00_axil_awready(axi_shared_cfg_AWREADY),
        .s00_axil_wdata(axi_shared_cfg_WDATA),
        .s00_axil_wstrb(axi_shared_cfg_WSTRB),
        .s00_axil_wvalid(axi_shared_cfg_WVALID),
        .s00_axil_wready(axi_shared_cfg_WREADY),
        .s00_axil_bresp(axi_shared_cfg_BRESP),
        .s00_axil_bvalid(axi_shared_cfg_BVALID),
        .s00_axil_bready(axi_shared_cfg_BREADY),
        .s00_axil_araddr(axi_shared_cfg_ARADDR),
        .s00_axil_arprot(0),
        .s00_axil_arvalid(axi_shared_cfg_ARVALID),
        .s00_axil_arready(axi_shared_cfg_ARREADY),
        .s00_axil_rdata(axi_shared_cfg_RDATA),
        .s00_axil_rresp(axi_shared_cfg_RRESP),
        .s00_axil_rvalid(axi_shared_cfg_RVALID),
        .s00_axil_rready(axi_shared_cfg_RREADY),

        // AXI-Lite Master Interface 0
        .m00_axil_awaddr(axi0_cfg_AWADDR),
        .m00_axil_awprot(),
        .m00_axil_awvalid(axi0_cfg_AWVALID),
        .m00_axil_awready(axi0_cfg_AWREADY),
        .m00_axil_wdata(axi0_cfg_WDATA),
        .m00_axil_wstrb(axi0_cfg_WSTRB),
        .m00_axil_wvalid(axi0_cfg_WVALID),
        .m00_axil_wready(axi0_cfg_WREADY),
        .m00_axil_bresp(axi0_cfg_BRESP),
        .m00_axil_bvalid(axi0_cfg_BVALID),
        .m00_axil_bready(axi0_cfg_BREADY),
        .m00_axil_araddr(axi0_cfg_ARADDR),
        .m00_axil_arprot(),
        .m00_axil_arvalid(axi0_cfg_ARVALID),
        .m00_axil_arready(axi0_cfg_ARREADY),
        .m00_axil_rdata(axi0_cfg_RDATA),
        .m00_axil_rresp(axi0_cfg_RRESP),
        .m00_axil_rvalid(axi0_cfg_RVALID),
        .m00_axil_rready(axi0_cfg_RREADY),

        // AXI-Lite Master Interface 1
        .m01_axil_awaddr(axi1_cfg_AWADDR),
        .m01_axil_awprot(),
        .m01_axil_awvalid(axi1_cfg_AWVALID),
        .m01_axil_awready(axi1_cfg_AWREADY),
        .m01_axil_wdata(axi1_cfg_WDATA),
        .m01_axil_wstrb(axi1_cfg_WSTRB),
        .m01_axil_wvalid(axi1_cfg_WVALID),
        .m01_axil_wready(axi1_cfg_WREADY),
        .m01_axil_bresp(axi1_cfg_BRESP),
        .m01_axil_bvalid(axi1_cfg_BVALID),
        .m01_axil_bready(axi1_cfg_BREADY),
        .m01_axil_araddr(axi1_cfg_ARADDR),
        .m01_axil_arprot(),
        .m01_axil_arvalid(axi1_cfg_ARVALID),
        .m01_axil_arready(axi1_cfg_ARREADY),
        .m01_axil_rdata(axi1_cfg_RDATA),
        .m01_axil_rresp(axi1_cfg_RRESP),
        .m01_axil_rvalid(axi1_cfg_RVALID),
        .m01_axil_rready(axi1_cfg_RREADY)
    );

    axi_axil_adapter #(
        .ADDR_WIDTH(8),
        .AXI_DATA_WIDTH(32),
        .AXI_STRB_WIDTH(4),
        .AXI_ID_WIDTH(8),                 // Slave AXI ID width
        .AXIL_DATA_WIDTH(32),     // Master AXI lite data width
        .AXIL_STRB_WIDTH(4),     // Master AXI lite wstrb width
        .CONVERT_BURST(1),                // Convert full-width burst
        .CONVERT_NARROW_BURST(0)          // Convert narrow burst
    ) axi_axil_adapter_inst (
        .clk(ap_clk),
        .rst(~ap_rst_n),

        // AXI Slave interface
        .s_axi_awid(s_axi_awid),
        .s_axi_awaddr(s_axi_awaddr),
        .s_axi_awlen(s_axi_awlen),
        .s_axi_awsize(s_axi_awsize),
        .s_axi_awburst(s_axi_awburst),
        .s_axi_awlock(s_axi_awlock),
        .s_axi_awcache(s_axi_awcache),
        .s_axi_awprot(s_axi_awprot),
        .s_axi_awvalid(s_axi_awvalid),
        .s_axi_awready(s_axi_awready),
        .s_axi_wdata(s_axi_wdata),
        .s_axi_wstrb(s_axi_wstrb),
        .s_axi_wlast(s_axi_wlast),
        .s_axi_wvalid(s_axi_wvalid),
        .s_axi_wready(s_axi_wready),
        .s_axi_bid(s_axi_bid),
        .s_axi_bresp(s_axi_bresp),
        .s_axi_bvalid(s_axi_bvalid),
        .s_axi_bready(s_axi_bready),
        .s_axi_arid(s_axi_arid),
        .s_axi_araddr(s_axi_araddr),
        .s_axi_arlen(s_axi_arlen),
        .s_axi_arsize(s_axi_arsize),
        .s_axi_arburst(s_axi_arburst),
        .s_axi_arlock(s_axi_arlock),
        .s_axi_arcache(s_axi_arcache),
        .s_axi_arprot(s_axi_arprot),
        .s_axi_arvalid(s_axi_arvalid),
        .s_axi_arready(s_axi_arready),
        .s_axi_rid(s_axi_rid),
        .s_axi_rdata(s_axi_rdata),
        .s_axi_rresp(s_axi_rresp),
        .s_axi_rlast(s_axi_rlast),
        .s_axi_rvalid(s_axi_rvalid),
        .s_axi_rready(s_axi_rready),

        // AXI Lite Master interface
        .m_axil_awaddr(axi_shared_cfg_AWADDR),
        .m_axil_awprot(),
        .m_axil_awvalid(axi_shared_cfg_AWVALID),
        .m_axil_awready(axi_shared_cfg_AWREADY),
        .m_axil_wdata(axi_shared_cfg_WDATA),
        .m_axil_wstrb(axi_shared_cfg_WSTRB),
        .m_axil_wvalid(axi_shared_cfg_WVALID),
        .m_axil_wready(axi_shared_cfg_WREADY),
        .m_axil_bresp(axi_shared_cfg_BRESP),
        .m_axil_bvalid(axi_shared_cfg_BVALID),
        .m_axil_bready(axi_shared_cfg_BREADY),
        .m_axil_araddr(axi_shared_cfg_ARADDR),
        .m_axil_arprot(),
        .m_axil_arvalid(axi_shared_cfg_ARVALID),
        .m_axil_arready(axi_shared_cfg_ARREADY),
        .m_axil_rdata(axi_shared_cfg_RDATA),
        .m_axil_rresp(axi_shared_cfg_RRESP),
        .m_axil_rvalid(axi_shared_cfg_RVALID),
        .m_axil_rready(axi_shared_cfg_RREADY)
    );


endmodule

// Content from axi_interconnect.v
/*

Copyright (c) 2018 Alex Forencich

Permission is hereby granted, free of charge, to any person obtaining a copy
of this software and associated documentation files (the "Software"), to deal
in the Software without restriction, including without limitation the rights
to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
copies of the Software, and to permit persons to whom the Software is
furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in
all copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY
FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
THE SOFTWARE.

*/

// Language: Verilog 2001

/*
 * AXI4 interconnect
 */
module axi_interconnect #
(
    // Number of AXI inputs (slave interfaces)
    parameter S_COUNT = 4,
    // Number of AXI outputs (master interfaces)
    parameter M_COUNT = 4,
    // Width of data bus in bits
    parameter DATA_WIDTH = 32,
    // Width of address bus in bits
    parameter ADDR_WIDTH = 32,
    // Width of wstrb (width of data bus in words)
    parameter STRB_WIDTH = (DATA_WIDTH/8),
    // Width of ID signal
    parameter ID_WIDTH = 8,
    // Propagate awuser signal
    parameter AWUSER_ENABLE = 0,
    // Width of awuser signal
    parameter AWUSER_WIDTH = 1,
    // Propagate wuser signal
    parameter WUSER_ENABLE = 0,
    // Width of wuser signal
    parameter WUSER_WIDTH = 1,
    // Propagate buser signal
    parameter BUSER_ENABLE = 0,
    // Width of buser signal
    parameter BUSER_WIDTH = 1,
    // Propagate aruser signal
    parameter ARUSER_ENABLE = 0,
    // Width of aruser signal
    parameter ARUSER_WIDTH = 1,
    // Propagate ruser signal
    parameter RUSER_ENABLE = 0,
    // Width of ruser signal
    parameter RUSER_WIDTH = 1,
    // Propagate ID field
    parameter FORWARD_ID = 0,
    // Number of regions per master interface
    parameter M_REGIONS = 1,
    // Master interface base addresses
    // M_COUNT concatenated fields of M_REGIONS concatenated fields of ADDR_WIDTH bits
    // set to zero for default addressing based on M_ADDR_WIDTH
    parameter M_BASE_ADDR = 0,
    // Master interface address widths
    // M_COUNT concatenated fields of M_REGIONS concatenated fields of 32 bits
    parameter M_ADDR_WIDTH = {M_COUNT{{M_REGIONS{32'd24}}}},
    // Read connections between interfaces
    // M_COUNT concatenated fields of S_COUNT bits
    parameter M_CONNECT_READ = {M_COUNT{{S_COUNT{1'b1}}}},
    // Write connections between interfaces
    // M_COUNT concatenated fields of S_COUNT bits
    parameter M_CONNECT_WRITE = {M_COUNT{{S_COUNT{1'b1}}}},
    // Secure master (fail operations based on awprot/arprot)
    // M_COUNT bits
    parameter M_SECURE = {M_COUNT{1'b0}}
) (

    input  wire                            clk,
    input  wire                            rst,

    /*
     * AXI slave interfaces
     */
    input  wire [S_COUNT*ID_WIDTH-1:0]     s_axi_awid,
    input  wire [S_COUNT*ADDR_WIDTH-1:0]   s_axi_awaddr,
    input  wire [S_COUNT*8-1:0]            s_axi_awlen,
    input  wire [S_COUNT*3-1:0]            s_axi_awsize,
    input  wire [S_COUNT*2-1:0]            s_axi_awburst,
    input  wire [S_COUNT-1:0]              s_axi_awlock,
    input  wire [S_COUNT*4-1:0]            s_axi_awcache,
    input  wire [S_COUNT*3-1:0]            s_axi_awprot,
    input  wire [S_COUNT*4-1:0]            s_axi_awqos,
    input  wire [S_COUNT*AWUSER_WIDTH-1:0] s_axi_awuser,
    input  wire [S_COUNT-1:0]              s_axi_awvalid,
    output wire [S_COUNT-1:0]              s_axi_awready,
    input  wire [S_COUNT*DATA_WIDTH-1:0]   s_axi_wdata,
    input  wire [S_COUNT*STRB_WIDTH-1:0]   s_axi_wstrb,
    input  wire [S_COUNT-1:0]              s_axi_wlast,
    input  wire [S_COUNT*WUSER_WIDTH-1:0]  s_axi_wuser,
    input  wire [S_COUNT-1:0]              s_axi_wvalid,
    output wire [S_COUNT-1:0]              s_axi_wready,
    output wire [S_COUNT*ID_WIDTH-1:0]     s_axi_bid,
    output wire [S_COUNT*2-1:0]            s_axi_bresp,
    output wire [S_COUNT*BUSER_WIDTH-1:0]  s_axi_buser,
    output wire [S_COUNT-1:0]              s_axi_bvalid,
    input  wire [S_COUNT-1:0]              s_axi_bready,
    input  wire [S_COUNT*ID_WIDTH-1:0]     s_axi_arid,
    input  wire [S_COUNT*ADDR_WIDTH-1:0]   s_axi_araddr,
    input  wire [S_COUNT*8-1:0]            s_axi_arlen,
    input  wire [S_COUNT*3-1:0]            s_axi_arsize,
    input  wire [S_COUNT*2-1:0]            s_axi_arburst,
    input  wire [S_COUNT-1:0]              s_axi_arlock,
    input  wire [S_COUNT*4-1:0]            s_axi_arcache,
    input  wire [S_COUNT*3-1:0]            s_axi_arprot,
    input  wire [S_COUNT*4-1:0]            s_axi_arqos,
    input  wire [S_COUNT*ARUSER_WIDTH-1:0] s_axi_aruser,
    input  wire [S_COUNT-1:0]              s_axi_arvalid,
    output wire [S_COUNT-1:0]              s_axi_arready,
    output wire [S_COUNT*ID_WIDTH-1:0]     s_axi_rid,
    output wire [S_COUNT*DATA_WIDTH-1:0]   s_axi_rdata,
    output wire [S_COUNT*2-1:0]            s_axi_rresp,
    output wire [S_COUNT-1:0]              s_axi_rlast,
    output wire [S_COUNT*RUSER_WIDTH-1:0]  s_axi_ruser,
    output wire [S_COUNT-1:0]              s_axi_rvalid,
    input  wire [S_COUNT-1:0]              s_axi_rready,

    /*
     * AXI master interfaces
     */
    output wire [M_COUNT*ID_WIDTH-1:0]     m_axi_awid,
    output wire [M_COUNT*ADDR_WIDTH-1:0]   m_axi_awaddr,
    output wire [M_COUNT*8-1:0]            m_axi_awlen,
    output wire [M_COUNT*3-1:0]            m_axi_awsize,
    output wire [M_COUNT*2-1:0]            m_axi_awburst,
    output wire [M_COUNT-1:0]              m_axi_awlock,
    output wire [M_COUNT*4-1:0]            m_axi_awcache,
    output wire [M_COUNT*3-1:0]            m_axi_awprot,
    output wire [M_COUNT*4-1:0]            m_axi_awqos,
    output wire [M_COUNT*4-1:0]            m_axi_awregion,
    output wire [M_COUNT*AWUSER_WIDTH-1:0] m_axi_awuser,
    output wire [M_COUNT-1:0]              m_axi_awvalid,
    input  wire [M_COUNT-1:0]              m_axi_awready,
    output wire [M_COUNT*DATA_WIDTH-1:0]   m_axi_wdata,
    output wire [M_COUNT*STRB_WIDTH-1:0]   m_axi_wstrb,
    output wire [M_COUNT-1:0]              m_axi_wlast,
    output wire [M_COUNT*WUSER_WIDTH-1:0]  m_axi_wuser,
    output wire [M_COUNT-1:0]              m_axi_wvalid,
    input  wire [M_COUNT-1:0]              m_axi_wready,
    input  wire [M_COUNT*ID_WIDTH-1:0]     m_axi_bid,
    input  wire [M_COUNT*2-1:0]            m_axi_bresp,
    input  wire [M_COUNT*BUSER_WIDTH-1:0]  m_axi_buser,
    input  wire [M_COUNT-1:0]              m_axi_bvalid,
    output wire [M_COUNT-1:0]              m_axi_bready,
    output wire [M_COUNT*ID_WIDTH-1:0]     m_axi_arid,
    output wire [M_COUNT*ADDR_WIDTH-1:0]   m_axi_araddr,
    output wire [M_COUNT*8-1:0]            m_axi_arlen,
    output wire [M_COUNT*3-1:0]            m_axi_arsize,
    output wire [M_COUNT*2-1:0]            m_axi_arburst,
    output wire [M_COUNT-1:0]              m_axi_arlock,
    output wire [M_COUNT*4-1:0]            m_axi_arcache,
    output wire [M_COUNT*3-1:0]            m_axi_arprot,
    output wire [M_COUNT*4-1:0]            m_axi_arqos,
    output wire [M_COUNT*4-1:0]            m_axi_arregion,
    output wire [M_COUNT*ARUSER_WIDTH-1:0] m_axi_aruser,
    output wire [M_COUNT-1:0]              m_axi_arvalid,
    input  wire [M_COUNT-1:0]              m_axi_arready,
    input  wire [M_COUNT*ID_WIDTH-1:0]     m_axi_rid,
    input  wire [M_COUNT*DATA_WIDTH-1:0]   m_axi_rdata,
    input  wire [M_COUNT*2-1:0]            m_axi_rresp,
    input  wire [M_COUNT-1:0]              m_axi_rlast,
    input  wire [M_COUNT*RUSER_WIDTH-1:0]  m_axi_ruser,
    input  wire [M_COUNT-1:0]              m_axi_rvalid,
    output wire [M_COUNT-1:0]              m_axi_rready
);

parameter CL_S_COUNT = $clog2(S_COUNT);
parameter CL_M_COUNT = $clog2(M_COUNT);

parameter AUSER_WIDTH = AWUSER_WIDTH > ARUSER_WIDTH ? AWUSER_WIDTH : ARUSER_WIDTH;

// default address computation
function [M_COUNT*M_REGIONS*ADDR_WIDTH-1:0] calcBaseAddrs(input [31:0] dummy);
    integer i;
    reg [ADDR_WIDTH-1:0] base;
    reg [ADDR_WIDTH-1:0] width;
    reg [ADDR_WIDTH-1:0] size;
    reg [ADDR_WIDTH-1:0] mask;
    begin
        calcBaseAddrs = {M_COUNT*M_REGIONS*ADDR_WIDTH{1'b0}};
        base = 0;
        for (i = 0; i < M_COUNT*M_REGIONS; i = i + 1) begin
            width = M_ADDR_WIDTH[i*32 +: 32];
            mask = {ADDR_WIDTH{1'b1}} >> (ADDR_WIDTH - width);
            size = mask + 1;
            if (width > 0) begin
                if ((base & mask) != 0) begin
                   base = base + size - (base & mask); // align
                end
                calcBaseAddrs[i * ADDR_WIDTH +: ADDR_WIDTH] = base;
                base = base + size; // increment
            end
        end
    end
endfunction

parameter M_BASE_ADDR_INT = M_BASE_ADDR ? M_BASE_ADDR : calcBaseAddrs(0);

integer i, j;

// check configuration
initial begin
    $display("Addressing configuration for axi_interconnect instance %m");
    for (i = 0; i < M_COUNT*M_REGIONS; i = i + 1) begin
        if (M_ADDR_WIDTH[i*32 +: 32]) begin
            $display("%2d (%2d): %x / %02d -- %x-%x",
                i/M_REGIONS, i%M_REGIONS,
                M_BASE_ADDR_INT[i*ADDR_WIDTH +: ADDR_WIDTH],
                M_ADDR_WIDTH[i*32 +: 32],
                M_BASE_ADDR_INT[i*ADDR_WIDTH +: ADDR_WIDTH] & ({ADDR_WIDTH{1'b1}} << M_ADDR_WIDTH[i*32 +: 32]),
                M_BASE_ADDR_INT[i*ADDR_WIDTH +: ADDR_WIDTH] | ({ADDR_WIDTH{1'b1}} >> (ADDR_WIDTH - M_ADDR_WIDTH[i*32 +: 32]))
            );
        end
    end

    for (i = 0; i < M_COUNT*M_REGIONS; i = i + 1) begin
        if ((M_BASE_ADDR_INT[i*ADDR_WIDTH +: ADDR_WIDTH] & (2**M_ADDR_WIDTH[i*32 +: 32]-1)) != 0) begin
            $display("Region not aligned:");
            $display("%2d (%2d): %x / %2d -- %x-%x",
                i/M_REGIONS, i%M_REGIONS,
                M_BASE_ADDR_INT[i*ADDR_WIDTH +: ADDR_WIDTH],
                M_ADDR_WIDTH[i*32 +: 32],
                M_BASE_ADDR_INT[i*ADDR_WIDTH +: ADDR_WIDTH] & ({ADDR_WIDTH{1'b1}} << M_ADDR_WIDTH[i*32 +: 32]),
                M_BASE_ADDR_INT[i*ADDR_WIDTH +: ADDR_WIDTH] | ({ADDR_WIDTH{1'b1}} >> (ADDR_WIDTH - M_ADDR_WIDTH[i*32 +: 32]))
            );
        end
    end

    for (i = 0; i < M_COUNT*M_REGIONS; i = i + 1) begin
        for (j = i+1; j < M_COUNT*M_REGIONS; j = j + 1) begin
            if (M_ADDR_WIDTH[i*32 +: 32] && M_ADDR_WIDTH[j*32 +: 32]) begin
                if (((M_BASE_ADDR_INT[i*ADDR_WIDTH +: ADDR_WIDTH] & ({ADDR_WIDTH{1'b1}} << M_ADDR_WIDTH[i*32 +: 32])) <= (M_BASE_ADDR_INT[j*ADDR_WIDTH +: ADDR_WIDTH] | ({ADDR_WIDTH{1'b1}} >> (ADDR_WIDTH - M_ADDR_WIDTH[j*32 +: 32]))))
                        && ((M_BASE_ADDR_INT[j*ADDR_WIDTH +: ADDR_WIDTH] & ({ADDR_WIDTH{1'b1}} << M_ADDR_WIDTH[j*32 +: 32])) <= (M_BASE_ADDR_INT[i*ADDR_WIDTH +: ADDR_WIDTH] | ({ADDR_WIDTH{1'b1}} >> (ADDR_WIDTH - M_ADDR_WIDTH[i*32 +: 32]))))) begin
                    $display("Overlapping regions:");
                    $display("%2d (%2d): %x / %2d -- %x-%x",
                        i/M_REGIONS, i%M_REGIONS,
                        M_BASE_ADDR_INT[i*ADDR_WIDTH +: ADDR_WIDTH],
                        M_ADDR_WIDTH[i*32 +: 32],
                        M_BASE_ADDR_INT[i*ADDR_WIDTH +: ADDR_WIDTH] & ({ADDR_WIDTH{1'b1}} << M_ADDR_WIDTH[i*32 +: 32]),
                        M_BASE_ADDR_INT[i*ADDR_WIDTH +: ADDR_WIDTH] | ({ADDR_WIDTH{1'b1}} >> (ADDR_WIDTH - M_ADDR_WIDTH[i*32 +: 32]))
                    );
                    $display("%2d (%2d): %x / %2d -- %x-%x",
                        j/M_REGIONS, j%M_REGIONS,
                        M_BASE_ADDR_INT[j*ADDR_WIDTH +: ADDR_WIDTH],
                        M_ADDR_WIDTH[j*32 +: 32],
                        M_BASE_ADDR_INT[j*ADDR_WIDTH +: ADDR_WIDTH] & ({ADDR_WIDTH{1'b1}} << M_ADDR_WIDTH[j*32 +: 32]),
                        M_BASE_ADDR_INT[j*ADDR_WIDTH +: ADDR_WIDTH] | ({ADDR_WIDTH{1'b1}} >> (ADDR_WIDTH - M_ADDR_WIDTH[j*32 +: 32]))
                    );
                end
            end
        end
    end
end

localparam [2:0]
    STATE_IDLE = 3'd0,
    STATE_DECODE = 3'd1,
    STATE_WRITE = 3'd2,
    STATE_WRITE_RESP = 3'd3,
    STATE_WRITE_DROP = 3'd4,
    STATE_READ = 3'd5,
    STATE_READ_DROP = 3'd6,
    STATE_WAIT_IDLE = 3'd7;

reg [2:0] state_reg = STATE_IDLE, state_next;

reg match;

reg [CL_M_COUNT-1:0] m_select_reg = 2'd0, m_select_next;
reg [ID_WIDTH-1:0] axi_id_reg = {ID_WIDTH{1'b0}}, axi_id_next;
reg [ADDR_WIDTH-1:0] axi_addr_reg = {ADDR_WIDTH{1'b0}}, axi_addr_next;
reg axi_addr_valid_reg = 1'b0, axi_addr_valid_next;
reg [7:0] axi_len_reg = 8'd0, axi_len_next;
reg [2:0] axi_size_reg = 3'd0, axi_size_next;
reg [1:0] axi_burst_reg = 2'd0, axi_burst_next;
reg axi_lock_reg = 1'b0, axi_lock_next;
reg [3:0] axi_cache_reg = 4'd0, axi_cache_next;
reg [2:0] axi_prot_reg = 3'b000, axi_prot_next;
reg [3:0] axi_qos_reg = 4'd0, axi_qos_next;
reg [3:0] axi_region_reg = 4'd0, axi_region_next;
reg [AUSER_WIDTH-1:0] axi_auser_reg = {AUSER_WIDTH{1'b0}}, axi_auser_next;
reg [1:0] axi_bresp_reg = 2'b00, axi_bresp_next;
reg [BUSER_WIDTH-1:0] axi_buser_reg = {BUSER_WIDTH{1'b0}}, axi_buser_next;

reg [S_COUNT-1:0] s_axi_awready_reg = 0, s_axi_awready_next;
reg [S_COUNT-1:0] s_axi_wready_reg = 0, s_axi_wready_next;
reg [S_COUNT-1:0] s_axi_bvalid_reg = 0, s_axi_bvalid_next;
reg [S_COUNT-1:0] s_axi_arready_reg = 0, s_axi_arready_next;

reg [M_COUNT-1:0] m_axi_awvalid_reg = 0, m_axi_awvalid_next;
reg [M_COUNT-1:0] m_axi_bready_reg = 0, m_axi_bready_next;
reg [M_COUNT-1:0] m_axi_arvalid_reg = 0, m_axi_arvalid_next;
reg [M_COUNT-1:0] m_axi_rready_reg = 0, m_axi_rready_next;

// internal datapath
reg  [ID_WIDTH-1:0]    s_axi_rid_int;
reg  [DATA_WIDTH-1:0]  s_axi_rdata_int;
reg  [1:0]             s_axi_rresp_int;
reg                    s_axi_rlast_int;
reg  [RUSER_WIDTH-1:0] s_axi_ruser_int;
reg                    s_axi_rvalid_int;
reg                    s_axi_rready_int_reg = 1'b0;
wire                   s_axi_rready_int_early;

reg  [DATA_WIDTH-1:0]  m_axi_wdata_int;
reg  [STRB_WIDTH-1:0]  m_axi_wstrb_int;
reg                    m_axi_wlast_int;
reg  [WUSER_WIDTH-1:0] m_axi_wuser_int;
reg                    m_axi_wvalid_int;
reg                    m_axi_wready_int_reg = 1'b0;
wire                   m_axi_wready_int_early;

assign s_axi_awready = s_axi_awready_reg;
assign s_axi_wready = s_axi_wready_reg;
assign s_axi_bid = {S_COUNT{axi_id_reg}};
assign s_axi_bresp = {S_COUNT{axi_bresp_reg}};
assign s_axi_buser = {S_COUNT{BUSER_ENABLE ? axi_buser_reg : {BUSER_WIDTH{1'b0}}}};
assign s_axi_bvalid = s_axi_bvalid_reg;
assign s_axi_arready = s_axi_arready_reg;

assign m_axi_awid = {M_COUNT{FORWARD_ID ? axi_id_reg : {ID_WIDTH{1'b0}}}};
assign m_axi_awaddr = {M_COUNT{axi_addr_reg}};
assign m_axi_awlen = {M_COUNT{axi_len_reg}};
assign m_axi_awsize = {M_COUNT{axi_size_reg}};
assign m_axi_awburst = {M_COUNT{axi_burst_reg}};
assign m_axi_awlock = {M_COUNT{axi_lock_reg}};
assign m_axi_awcache = {M_COUNT{axi_cache_reg}};
assign m_axi_awprot = {M_COUNT{axi_prot_reg}};
assign m_axi_awqos = {M_COUNT{axi_qos_reg}};
assign m_axi_awregion = {M_COUNT{axi_region_reg}};
assign m_axi_awuser = {M_COUNT{AWUSER_ENABLE ? axi_auser_reg[AWUSER_WIDTH-1:0] : {AWUSER_WIDTH{1'b0}}}};
assign m_axi_awvalid = m_axi_awvalid_reg;
assign m_axi_bready = m_axi_bready_reg;
assign m_axi_arid = {M_COUNT{FORWARD_ID ? axi_id_reg : {ID_WIDTH{1'b0}}}};
assign m_axi_araddr = {M_COUNT{axi_addr_reg}};
assign m_axi_arlen = {M_COUNT{axi_len_reg}};
assign m_axi_arsize = {M_COUNT{axi_size_reg}};
assign m_axi_arburst = {M_COUNT{axi_burst_reg}};
assign m_axi_arlock = {M_COUNT{axi_lock_reg}};
assign m_axi_arcache = {M_COUNT{axi_cache_reg}};
assign m_axi_arprot = {M_COUNT{axi_prot_reg}};
assign m_axi_arqos = {M_COUNT{axi_qos_reg}};
assign m_axi_arregion = {M_COUNT{axi_region_reg}};
assign m_axi_aruser = {M_COUNT{ARUSER_ENABLE ? axi_auser_reg[ARUSER_WIDTH-1:0] : {ARUSER_WIDTH{1'b0}}}};
assign m_axi_arvalid = m_axi_arvalid_reg;
assign m_axi_rready = m_axi_rready_reg;

// slave side mux
wire [(CL_S_COUNT > 0 ? CL_S_COUNT-1 : 0):0] s_select;

wire [ID_WIDTH-1:0]     current_s_axi_awid      = s_axi_awid[s_select*ID_WIDTH +: ID_WIDTH];
wire [ADDR_WIDTH-1:0]   current_s_axi_awaddr    = s_axi_awaddr[s_select*ADDR_WIDTH +: ADDR_WIDTH];
wire [7:0]              current_s_axi_awlen     = s_axi_awlen[s_select*8 +: 8];
wire [2:0]              current_s_axi_awsize    = s_axi_awsize[s_select*3 +: 3];
wire [1:0]              current_s_axi_awburst   = s_axi_awburst[s_select*2 +: 2];
wire                    current_s_axi_awlock    = s_axi_awlock[s_select];
wire [3:0]              current_s_axi_awcache   = s_axi_awcache[s_select*4 +: 4];
wire [2:0]              current_s_axi_awprot    = s_axi_awprot[s_select*3 +: 3];
wire [3:0]              current_s_axi_awqos     = s_axi_awqos[s_select*4 +: 4];
wire [AWUSER_WIDTH-1:0] current_s_axi_awuser    = s_axi_awuser[s_select*AWUSER_WIDTH +: AWUSER_WIDTH];
wire                    current_s_axi_awvalid   = s_axi_awvalid[s_select];
wire                    current_s_axi_awready   = s_axi_awready[s_select];
wire [DATA_WIDTH-1:0]   current_s_axi_wdata     = s_axi_wdata[s_select*DATA_WIDTH +: DATA_WIDTH];
wire [STRB_WIDTH-1:0]   current_s_axi_wstrb     = s_axi_wstrb[s_select*STRB_WIDTH +: STRB_WIDTH];
wire                    current_s_axi_wlast     = s_axi_wlast[s_select];
wire [WUSER_WIDTH-1:0]  current_s_axi_wuser     = s_axi_wuser[s_select*WUSER_WIDTH +: WUSER_WIDTH];
wire                    current_s_axi_wvalid    = s_axi_wvalid[s_select];
wire                    current_s_axi_wready    = s_axi_wready[s_select];
wire [ID_WIDTH-1:0]     current_s_axi_bid       = s_axi_bid[s_select*ID_WIDTH +: ID_WIDTH];
wire [1:0]              current_s_axi_bresp     = s_axi_bresp[s_select*2 +: 2];
wire [BUSER_WIDTH-1:0]  current_s_axi_buser     = s_axi_buser[s_select*BUSER_WIDTH +: BUSER_WIDTH];
wire                    current_s_axi_bvalid    = s_axi_bvalid[s_select];
wire                    current_s_axi_bready    = s_axi_bready[s_select];
wire [ID_WIDTH-1:0]     current_s_axi_arid      = s_axi_arid[s_select*ID_WIDTH +: ID_WIDTH];
wire [ADDR_WIDTH-1:0]   current_s_axi_araddr    = s_axi_araddr[s_select*ADDR_WIDTH +: ADDR_WIDTH];
wire [7:0]              current_s_axi_arlen     = s_axi_arlen[s_select*8 +: 8];
wire [2:0]              current_s_axi_arsize    = s_axi_arsize[s_select*3 +: 3];
wire [1:0]              current_s_axi_arburst   = s_axi_arburst[s_select*2 +: 2];
wire                    current_s_axi_arlock    = s_axi_arlock[s_select];
wire [3:0]              current_s_axi_arcache   = s_axi_arcache[s_select*4 +: 4];
wire [2:0]              current_s_axi_arprot    = s_axi_arprot[s_select*3 +: 3];
wire [3:0]              current_s_axi_arqos     = s_axi_arqos[s_select*4 +: 4];
wire [ARUSER_WIDTH-1:0] current_s_axi_aruser    = s_axi_aruser[s_select*ARUSER_WIDTH +: ARUSER_WIDTH];
wire                    current_s_axi_arvalid   = s_axi_arvalid[s_select];
wire                    current_s_axi_arready   = s_axi_arready[s_select];
wire [ID_WIDTH-1:0]     current_s_axi_rid       = s_axi_rid[s_select*ID_WIDTH +: ID_WIDTH];
wire [DATA_WIDTH-1:0]   current_s_axi_rdata     = s_axi_rdata[s_select*DATA_WIDTH +: DATA_WIDTH];
wire [1:0]              current_s_axi_rresp     = s_axi_rresp[s_select*2 +: 2];
wire                    current_s_axi_rlast     = s_axi_rlast[s_select];
wire [RUSER_WIDTH-1:0]  current_s_axi_ruser     = s_axi_ruser[s_select*RUSER_WIDTH +: RUSER_WIDTH];
wire                    current_s_axi_rvalid    = s_axi_rvalid[s_select];
wire                    current_s_axi_rready    = s_axi_rready[s_select];

// master side mux
wire [ID_WIDTH-1:0]     current_m_axi_awid      = m_axi_awid[m_select_reg*ID_WIDTH +: ID_WIDTH];
wire [ADDR_WIDTH-1:0]   current_m_axi_awaddr    = m_axi_awaddr[m_select_reg*ADDR_WIDTH +: ADDR_WIDTH];
wire [7:0]              current_m_axi_awlen     = m_axi_awlen[m_select_reg*8 +: 8];
wire [2:0]              current_m_axi_awsize    = m_axi_awsize[m_select_reg*3 +: 3];
wire [1:0]              current_m_axi_awburst   = m_axi_awburst[m_select_reg*2 +: 2];
wire                    current_m_axi_awlock    = m_axi_awlock[m_select_reg];
wire [3:0]              current_m_axi_awcache   = m_axi_awcache[m_select_reg*4 +: 4];
wire [2:0]              current_m_axi_awprot    = m_axi_awprot[m_select_reg*3 +: 3];
wire [3:0]              current_m_axi_awqos     = m_axi_awqos[m_select_reg*4 +: 4];
wire [3:0]              current_m_axi_awregion  = m_axi_awregion[m_select_reg*4 +: 4];
wire [AWUSER_WIDTH-1:0] current_m_axi_awuser    = m_axi_awuser[m_select_reg*AWUSER_WIDTH +: AWUSER_WIDTH];
wire                    current_m_axi_awvalid   = m_axi_awvalid[m_select_reg];
wire                    current_m_axi_awready   = m_axi_awready[m_select_reg];
wire [DATA_WIDTH-1:0]   current_m_axi_wdata     = m_axi_wdata[m_select_reg*DATA_WIDTH +: DATA_WIDTH];
wire [STRB_WIDTH-1:0]   current_m_axi_wstrb     = m_axi_wstrb[m_select_reg*STRB_WIDTH +: STRB_WIDTH];
wire                    current_m_axi_wlast     = m_axi_wlast[m_select_reg];
wire [WUSER_WIDTH-1:0]  current_m_axi_wuser     = m_axi_wuser[m_select_reg*WUSER_WIDTH +: WUSER_WIDTH];
wire                    current_m_axi_wvalid    = m_axi_wvalid[m_select_reg];
wire                    current_m_axi_wready    = m_axi_wready[m_select_reg];
wire [ID_WIDTH-1:0]     current_m_axi_bid       = m_axi_bid[m_select_reg*ID_WIDTH +: ID_WIDTH];
wire [1:0]              current_m_axi_bresp     = m_axi_bresp[m_select_reg*2 +: 2];
wire [BUSER_WIDTH-1:0]  current_m_axi_buser     = m_axi_buser[m_select_reg*BUSER_WIDTH +: BUSER_WIDTH];
wire                    current_m_axi_bvalid    = m_axi_bvalid[m_select_reg];
wire                    current_m_axi_bready    = m_axi_bready[m_select_reg];
wire [ID_WIDTH-1:0]     current_m_axi_arid      = m_axi_arid[m_select_reg*ID_WIDTH +: ID_WIDTH];
wire [ADDR_WIDTH-1:0]   current_m_axi_araddr    = m_axi_araddr[m_select_reg*ADDR_WIDTH +: ADDR_WIDTH];
wire [7:0]              current_m_axi_arlen     = m_axi_arlen[m_select_reg*8 +: 8];
wire [2:0]              current_m_axi_arsize    = m_axi_arsize[m_select_reg*3 +: 3];
wire [1:0]              current_m_axi_arburst   = m_axi_arburst[m_select_reg*2 +: 2];
wire                    current_m_axi_arlock    = m_axi_arlock[m_select_reg];
wire [3:0]              current_m_axi_arcache   = m_axi_arcache[m_select_reg*4 +: 4];
wire [2:0]              current_m_axi_arprot    = m_axi_arprot[m_select_reg*3 +: 3];
wire [3:0]              current_m_axi_arqos     = m_axi_arqos[m_select_reg*4 +: 4];
wire [3:0]              current_m_axi_arregion  = m_axi_arregion[m_select_reg*4 +: 4];
wire [ARUSER_WIDTH-1:0] current_m_axi_aruser    = m_axi_aruser[m_select_reg*ARUSER_WIDTH +: ARUSER_WIDTH];
wire                    current_m_axi_arvalid   = m_axi_arvalid[m_select_reg];
wire                    current_m_axi_arready   = m_axi_arready[m_select_reg];
wire [ID_WIDTH-1:0]     current_m_axi_rid       = m_axi_rid[m_select_reg*ID_WIDTH +: ID_WIDTH];
wire [DATA_WIDTH-1:0]   current_m_axi_rdata     = m_axi_rdata[m_select_reg*DATA_WIDTH +: DATA_WIDTH];
wire [1:0]              current_m_axi_rresp     = m_axi_rresp[m_select_reg*2 +: 2];
wire                    current_m_axi_rlast     = m_axi_rlast[m_select_reg];
wire [RUSER_WIDTH-1:0]  current_m_axi_ruser     = m_axi_ruser[m_select_reg*RUSER_WIDTH +: RUSER_WIDTH];
wire                    current_m_axi_rvalid    = m_axi_rvalid[m_select_reg];
wire                    current_m_axi_rready    = m_axi_rready[m_select_reg];

// arbiter instance
wire [S_COUNT*2-1:0] request;
wire [S_COUNT*2-1:0] acknowledge;
wire [S_COUNT*2-1:0] grant;
wire grant_valid;
wire [CL_S_COUNT:0] grant_encoded;

wire read = grant_encoded[0];
assign s_select = grant_encoded >> 1;

arbiter #(
    .PORTS(S_COUNT*2),
    .ARB_TYPE_ROUND_ROBIN(1),
    .ARB_BLOCK(1),
    .ARB_BLOCK_ACK(1),
    .ARB_LSB_HIGH_PRIORITY(1)
)
arb_inst (
    .clk(clk),
    .rst(rst),
    .request(request),
    .acknowledge(acknowledge),
    .grant(grant),
    .grant_valid(grant_valid),
    .grant_encoded(grant_encoded)
);

genvar n;

// request generation
generate
for (n = 0; n < S_COUNT; n = n + 1) begin
    assign request[2*n]   = s_axi_awvalid[n];
    assign request[2*n+1] = s_axi_arvalid[n];
end
endgenerate

// acknowledge generation
generate
for (n = 0; n < S_COUNT; n = n + 1) begin
    assign acknowledge[2*n]   = grant[2*n]   && s_axi_bvalid[n] && s_axi_bready[n];
    assign acknowledge[2*n+1] = grant[2*n+1] && s_axi_rvalid[n] && s_axi_rready[n] && s_axi_rlast[n];
end
endgenerate

always @* begin
    state_next = STATE_IDLE;

    match = 1'b0;

    m_select_next = m_select_reg;
    axi_id_next = axi_id_reg;
    axi_addr_next = axi_addr_reg;
    axi_addr_valid_next = axi_addr_valid_reg;
    axi_len_next = axi_len_reg;
    axi_size_next = axi_size_reg;
    axi_burst_next = axi_burst_reg;
    axi_lock_next = axi_lock_reg;
    axi_cache_next = axi_cache_reg;
    axi_prot_next = axi_prot_reg;
    axi_qos_next = axi_qos_reg;
    axi_region_next = axi_region_reg;
    axi_auser_next = axi_auser_reg;
    axi_bresp_next = axi_bresp_reg;
    axi_buser_next = axi_buser_reg;

    s_axi_awready_next = 0;
    s_axi_wready_next = 0;
    s_axi_bvalid_next = s_axi_bvalid_reg & ~s_axi_bready;
    s_axi_arready_next = 0;

    m_axi_awvalid_next = m_axi_awvalid_reg & ~m_axi_awready;
    m_axi_bready_next = 0;
    m_axi_arvalid_next = m_axi_arvalid_reg & ~m_axi_arready;
    m_axi_rready_next = 0;

    s_axi_rid_int = axi_id_reg;
    s_axi_rdata_int = current_m_axi_rdata;
    s_axi_rresp_int = current_m_axi_rresp;
    s_axi_rlast_int = current_m_axi_rlast;
    s_axi_ruser_int = current_m_axi_ruser;
    s_axi_rvalid_int = 1'b0;

    m_axi_wdata_int = current_s_axi_wdata;
    m_axi_wstrb_int = current_s_axi_wstrb;
    m_axi_wlast_int = current_s_axi_wlast;
    m_axi_wuser_int = current_s_axi_wuser;
    m_axi_wvalid_int = 1'b0;

    case (state_reg)
        STATE_IDLE: begin
            // idle state; wait for arbitration

            if (grant_valid) begin

                axi_addr_valid_next = 1'b1;

                if (read) begin
                    // reading
                    axi_addr_next = current_s_axi_araddr;
                    axi_prot_next = current_s_axi_arprot;
                    axi_id_next = current_s_axi_arid;
                    axi_addr_next = current_s_axi_araddr;
                    axi_len_next = current_s_axi_arlen;
                    axi_size_next = current_s_axi_arsize;
                    axi_burst_next = current_s_axi_arburst;
                    axi_lock_next = current_s_axi_arlock;
                    axi_cache_next = current_s_axi_arcache;
                    axi_prot_next = current_s_axi_arprot;
                    axi_qos_next = current_s_axi_arqos;
                    axi_auser_next = current_s_axi_aruser;
                    s_axi_arready_next[s_select] = 1'b1;
                end else  begin
                    // writing
                    axi_addr_next = current_s_axi_awaddr;
                    axi_prot_next = current_s_axi_awprot;
                    axi_id_next = current_s_axi_awid;
                    axi_addr_next = current_s_axi_awaddr;
                    axi_len_next = current_s_axi_awlen;
                    axi_size_next = current_s_axi_awsize;
                    axi_burst_next = current_s_axi_awburst;
                    axi_lock_next = current_s_axi_awlock;
                    axi_cache_next = current_s_axi_awcache;
                    axi_prot_next = current_s_axi_awprot;
                    axi_qos_next = current_s_axi_awqos;
                    axi_auser_next = current_s_axi_awuser;
                    s_axi_awready_next[s_select] = 1'b1;
                end

                state_next = STATE_DECODE;
            end else begin
                state_next = STATE_IDLE;
            end
        end
        STATE_DECODE: begin
            // decode state; determine master interface

            match = 1'b0;
            for (i = 0; i < M_COUNT; i = i + 1) begin
                for (j = 0; j < M_REGIONS; j = j + 1) begin
                    if (M_ADDR_WIDTH[(i*M_REGIONS+j)*32 +: 32] && (!M_SECURE[i] || !axi_prot_reg[1]) && ((read ? M_CONNECT_READ : M_CONNECT_WRITE) & (1 << (s_select+i*S_COUNT))) && (axi_addr_reg >> M_ADDR_WIDTH[(i*M_REGIONS+j)*32 +: 32]) == (M_BASE_ADDR_INT[(i*M_REGIONS+j)*ADDR_WIDTH +: ADDR_WIDTH] >> M_ADDR_WIDTH[(i*M_REGIONS+j)*32 +: 32])) begin
                        m_select_next = i;
                        axi_region_next = j;
                        match = 1'b1;
                    end
                end
            end

            if (match) begin
                if (read) begin
                    // reading
                    m_axi_rready_next[m_select_reg] = s_axi_rready_int_early;
                    state_next = STATE_READ;
                end else begin
                    // writing
                    s_axi_wready_next[s_select] = m_axi_wready_int_early;
                    state_next = STATE_WRITE;
                end
            end else begin
                // no match; return decode error
                if (read) begin
                    // reading
                    state_next = STATE_READ_DROP;
                end else begin
                    // writing
                    axi_bresp_next = 2'b11;
                    s_axi_wready_next[s_select] = 1'b1;
                    state_next = STATE_WRITE_DROP;
                end
            end
        end
        STATE_WRITE: begin
            // write state; store and forward write data
            s_axi_wready_next[s_select] = m_axi_wready_int_early;

            if (axi_addr_valid_reg) begin
                m_axi_awvalid_next[m_select_reg] = 1'b1;
            end
            axi_addr_valid_next = 1'b0;

            if (current_s_axi_wready && current_s_axi_wvalid) begin
                m_axi_wdata_int = current_s_axi_wdata;
                m_axi_wstrb_int = current_s_axi_wstrb;
                m_axi_wlast_int = current_s_axi_wlast;
                m_axi_wuser_int = current_s_axi_wuser;
                m_axi_wvalid_int = 1'b1;

                if (current_s_axi_wlast) begin
                    s_axi_wready_next[s_select] = 1'b0;
                    m_axi_bready_next[m_select_reg] = 1'b1;
                    state_next = STATE_WRITE_RESP;
                end else begin
                    state_next = STATE_WRITE;
                end
            end else begin
                state_next = STATE_WRITE;
            end
        end
        STATE_WRITE_RESP: begin
            // write response state; store and forward write response
            m_axi_bready_next[m_select_reg] = 1'b1;

            if (current_m_axi_bready && current_m_axi_bvalid) begin
                m_axi_bready_next[m_select_reg] = 1'b0;
                axi_bresp_next = current_m_axi_bresp;
                s_axi_bvalid_next[s_select] = 1'b1;
                state_next = STATE_WAIT_IDLE;
            end else begin
                state_next = STATE_WRITE_RESP;
            end
        end
        STATE_WRITE_DROP: begin
            // write drop state; drop write data
            s_axi_wready_next[s_select] = 1'b1;

            axi_addr_valid_next = 1'b0;

            if (current_s_axi_wready && current_s_axi_wvalid && current_s_axi_wlast) begin
                s_axi_wready_next[s_select] = 1'b0;
                s_axi_bvalid_next[s_select] = 1'b1;
                state_next = STATE_WAIT_IDLE;
            end else begin
                state_next = STATE_WRITE_DROP;
            end
        end
        STATE_READ: begin
            // read state; store and forward read response
            m_axi_rready_next[m_select_reg] = s_axi_rready_int_early;

            if (axi_addr_valid_reg) begin
                m_axi_arvalid_next[m_select_reg] = 1'b1;
            end
            axi_addr_valid_next = 1'b0;

            if (current_m_axi_rready && current_m_axi_rvalid) begin
                s_axi_rid_int = axi_id_reg;
                s_axi_rdata_int = current_m_axi_rdata;
                s_axi_rresp_int = current_m_axi_rresp;
                s_axi_rlast_int = current_m_axi_rlast;
                s_axi_ruser_int = current_m_axi_ruser;
                s_axi_rvalid_int = 1'b1;

                if (current_m_axi_rlast) begin
                    m_axi_rready_next[m_select_reg] = 1'b0;
                    state_next = STATE_WAIT_IDLE;
                end else begin
                    state_next = STATE_READ;
                end
            end else begin
                state_next = STATE_READ;
            end
        end
        STATE_READ_DROP: begin
            // read drop state; generate decode error read response

            s_axi_rid_int = axi_id_reg;
            s_axi_rdata_int = {DATA_WIDTH{1'b0}};
            s_axi_rresp_int = 2'b11;
            s_axi_rlast_int = axi_len_reg == 0;
            s_axi_ruser_int = {RUSER_WIDTH{1'b0}};
            s_axi_rvalid_int = 1'b1;

            if (s_axi_rready_int_reg) begin
                axi_len_next = axi_len_reg - 1;
                if (axi_len_reg == 0) begin
                    state_next = STATE_WAIT_IDLE;
                end else begin
                    state_next = STATE_READ_DROP;
                end
            end else begin
                state_next = STATE_READ_DROP;
            end
        end
        STATE_WAIT_IDLE: begin
            // wait for idle state; wait untl grant valid is deasserted

            if (!grant_valid || acknowledge) begin
                state_next = STATE_IDLE;
            end else begin
                state_next = STATE_WAIT_IDLE;
            end
        end
    endcase
end

always @(posedge clk) begin
    if (rst) begin
        state_reg <= STATE_IDLE;

        s_axi_awready_reg <= 0;
        s_axi_wready_reg <= 0;
        s_axi_bvalid_reg <= 0;
        s_axi_arready_reg <= 0;

        m_axi_awvalid_reg <= 0;
        m_axi_bready_reg <= 0;
        m_axi_arvalid_reg <= 0;
        m_axi_rready_reg <= 0;
    end else begin
        state_reg <= state_next;

        s_axi_awready_reg <= s_axi_awready_next;
        s_axi_wready_reg <= s_axi_wready_next;
        s_axi_bvalid_reg <= s_axi_bvalid_next;
        s_axi_arready_reg <= s_axi_arready_next;

        m_axi_awvalid_reg <= m_axi_awvalid_next;
        m_axi_bready_reg <= m_axi_bready_next;
        m_axi_arvalid_reg <= m_axi_arvalid_next;
        m_axi_rready_reg <= m_axi_rready_next;
    end

    m_select_reg <= m_select_next;
    axi_id_reg <= axi_id_next;
    axi_addr_reg <= axi_addr_next;
    axi_addr_valid_reg <= axi_addr_valid_next;
    axi_len_reg <= axi_len_next;
    axi_size_reg <= axi_size_next;
    axi_burst_reg <= axi_burst_next;
    axi_lock_reg <= axi_lock_next;
    axi_cache_reg <= axi_cache_next;
    axi_prot_reg <= axi_prot_next;
    axi_qos_reg <= axi_qos_next;
    axi_region_reg <= axi_region_next;
    axi_auser_reg <= axi_auser_next;
    axi_bresp_reg <= axi_bresp_next;
    axi_buser_reg <= axi_buser_next;
end

// output datapath logic (R channel)
reg [ID_WIDTH-1:0]    s_axi_rid_reg    = {ID_WIDTH{1'b0}};
reg [DATA_WIDTH-1:0]  s_axi_rdata_reg  = {DATA_WIDTH{1'b0}};
reg [1:0]             s_axi_rresp_reg  = 2'd0;
reg                   s_axi_rlast_reg  = 1'b0;
reg [RUSER_WIDTH-1:0] s_axi_ruser_reg  = 1'b0;
reg [S_COUNT-1:0]     s_axi_rvalid_reg = 1'b0, s_axi_rvalid_next;

reg [ID_WIDTH-1:0]    temp_s_axi_rid_reg    = {ID_WIDTH{1'b0}};
reg [DATA_WIDTH-1:0]  temp_s_axi_rdata_reg  = {DATA_WIDTH{1'b0}};
reg [1:0]             temp_s_axi_rresp_reg  = 2'd0;
reg                   temp_s_axi_rlast_reg  = 1'b0;
reg [RUSER_WIDTH-1:0] temp_s_axi_ruser_reg  = 1'b0;
reg                   temp_s_axi_rvalid_reg = 1'b0, temp_s_axi_rvalid_next;

// datapath control
reg store_axi_r_int_to_output;
reg store_axi_r_int_to_temp;
reg store_axi_r_temp_to_output;

assign s_axi_rid = {S_COUNT{s_axi_rid_reg}};
assign s_axi_rdata = {S_COUNT{s_axi_rdata_reg}};
assign s_axi_rresp = {S_COUNT{s_axi_rresp_reg}};
assign s_axi_rlast = {S_COUNT{s_axi_rlast_reg}};
assign s_axi_ruser = {S_COUNT{RUSER_ENABLE ? s_axi_ruser_reg : {RUSER_WIDTH{1'b0}}}};
assign s_axi_rvalid = s_axi_rvalid_reg;

// enable ready input next cycle if output is ready or the temp reg will not be filled on the next cycle (output reg empty or no input)
assign s_axi_rready_int_early = current_s_axi_rready | (~temp_s_axi_rvalid_reg & (~current_s_axi_rvalid | ~s_axi_rvalid_int));

always @* begin
    // transfer sink ready state to source
    s_axi_rvalid_next = s_axi_rvalid_reg;
    temp_s_axi_rvalid_next = temp_s_axi_rvalid_reg;

    store_axi_r_int_to_output = 1'b0;
    store_axi_r_int_to_temp = 1'b0;
    store_axi_r_temp_to_output = 1'b0;

    if (s_axi_rready_int_reg) begin
        // input is ready
        if (current_s_axi_rready | ~current_s_axi_rvalid) begin
            // output is ready or currently not valid, transfer data to output
            s_axi_rvalid_next[s_select] = s_axi_rvalid_int;
            store_axi_r_int_to_output = 1'b1;
        end else begin
            // output is not ready, store input in temp
            temp_s_axi_rvalid_next = s_axi_rvalid_int;
            store_axi_r_int_to_temp = 1'b1;
        end
    end else if (current_s_axi_rready) begin
        // input is not ready, but output is ready
        s_axi_rvalid_next[s_select] = temp_s_axi_rvalid_reg;
        temp_s_axi_rvalid_next = 1'b0;
        store_axi_r_temp_to_output = 1'b1;
    end
end

always @(posedge clk) begin
    if (rst) begin
        s_axi_rvalid_reg <= 1'b0;
        s_axi_rready_int_reg <= 1'b0;
        temp_s_axi_rvalid_reg <= 1'b0;
    end else begin
        s_axi_rvalid_reg <= s_axi_rvalid_next;
        s_axi_rready_int_reg <= s_axi_rready_int_early;
        temp_s_axi_rvalid_reg <= temp_s_axi_rvalid_next;
    end

    // datapath
    if (store_axi_r_int_to_output) begin
        s_axi_rid_reg <= s_axi_rid_int;
        s_axi_rdata_reg <= s_axi_rdata_int;
        s_axi_rresp_reg <= s_axi_rresp_int;
        s_axi_rlast_reg <= s_axi_rlast_int;
        s_axi_ruser_reg <= s_axi_ruser_int;
    end else if (store_axi_r_temp_to_output) begin
        s_axi_rid_reg <= temp_s_axi_rid_reg;
        s_axi_rdata_reg <= temp_s_axi_rdata_reg;
        s_axi_rresp_reg <= temp_s_axi_rresp_reg;
        s_axi_rlast_reg <= temp_s_axi_rlast_reg;
        s_axi_ruser_reg <= temp_s_axi_ruser_reg;
    end

    if (store_axi_r_int_to_temp) begin
        temp_s_axi_rid_reg <= s_axi_rid_int;
        temp_s_axi_rdata_reg <= s_axi_rdata_int;
        temp_s_axi_rresp_reg <= s_axi_rresp_int;
        temp_s_axi_rlast_reg <= s_axi_rlast_int;
        temp_s_axi_ruser_reg <= s_axi_ruser_int;
    end
end

// output datapath logic (W channel)
reg [DATA_WIDTH-1:0]  m_axi_wdata_reg  = {DATA_WIDTH{1'b0}};
reg [STRB_WIDTH-1:0]  m_axi_wstrb_reg  = {STRB_WIDTH{1'b0}};
reg                   m_axi_wlast_reg  = 1'b0;
reg [WUSER_WIDTH-1:0] m_axi_wuser_reg  = 1'b0;
reg [M_COUNT-1:0]     m_axi_wvalid_reg = 1'b0, m_axi_wvalid_next;

reg [DATA_WIDTH-1:0]  temp_m_axi_wdata_reg  = {DATA_WIDTH{1'b0}};
reg [STRB_WIDTH-1:0]  temp_m_axi_wstrb_reg  = {STRB_WIDTH{1'b0}};
reg                   temp_m_axi_wlast_reg  = 1'b0;
reg [WUSER_WIDTH-1:0] temp_m_axi_wuser_reg  = 1'b0;
reg                   temp_m_axi_wvalid_reg = 1'b0, temp_m_axi_wvalid_next;

// datapath control
reg store_axi_w_int_to_output;
reg store_axi_w_int_to_temp;
reg store_axi_w_temp_to_output;

assign m_axi_wdata = {M_COUNT{m_axi_wdata_reg}};
assign m_axi_wstrb = {M_COUNT{m_axi_wstrb_reg}};
assign m_axi_wlast = {M_COUNT{m_axi_wlast_reg}};
assign m_axi_wuser = {M_COUNT{WUSER_ENABLE ? m_axi_wuser_reg : {WUSER_WIDTH{1'b0}}}};
assign m_axi_wvalid = m_axi_wvalid_reg;

// enable ready input next cycle if output is ready or the temp reg will not be filled on the next cycle (output reg empty or no input)
assign m_axi_wready_int_early = current_m_axi_wready | (~temp_m_axi_wvalid_reg & (~current_m_axi_wvalid | ~m_axi_wvalid_int));

always @* begin
    // transfer sink ready state to source
    m_axi_wvalid_next = m_axi_wvalid_reg;
    temp_m_axi_wvalid_next = temp_m_axi_wvalid_reg;

    store_axi_w_int_to_output = 1'b0;
    store_axi_w_int_to_temp = 1'b0;
    store_axi_w_temp_to_output = 1'b0;

    if (m_axi_wready_int_reg) begin
        // input is ready
        if (current_m_axi_wready | ~current_m_axi_wvalid) begin
            // output is ready or currently not valid, transfer data to output
            m_axi_wvalid_next[m_select_reg] = m_axi_wvalid_int;
            store_axi_w_int_to_output = 1'b1;
        end else begin
            // output is not ready, store input in temp
            temp_m_axi_wvalid_next = m_axi_wvalid_int;
            store_axi_w_int_to_temp = 1'b1;
        end
    end else if (current_m_axi_wready) begin
        // input is not ready, but output is ready
        m_axi_wvalid_next[m_select_reg] = temp_m_axi_wvalid_reg;
        temp_m_axi_wvalid_next = 1'b0;
        store_axi_w_temp_to_output = 1'b1;
    end
end

always @(posedge clk) begin
    if (rst) begin
        m_axi_wvalid_reg <= 1'b0;
        m_axi_wready_int_reg <= 1'b0;
        temp_m_axi_wvalid_reg <= 1'b0;
    end else begin
        m_axi_wvalid_reg <= m_axi_wvalid_next;
        m_axi_wready_int_reg <= m_axi_wready_int_early;
        temp_m_axi_wvalid_reg <= temp_m_axi_wvalid_next;
    end

    // datapath
    if (store_axi_w_int_to_output) begin
        m_axi_wdata_reg <= m_axi_wdata_int;
        m_axi_wstrb_reg <= m_axi_wstrb_int;
        m_axi_wlast_reg <= m_axi_wlast_int;
        m_axi_wuser_reg <= m_axi_wuser_int;
    end else if (store_axi_w_temp_to_output) begin
        m_axi_wdata_reg <= temp_m_axi_wdata_reg;
        m_axi_wstrb_reg <= temp_m_axi_wstrb_reg;
        m_axi_wlast_reg <= temp_m_axi_wlast_reg;
        m_axi_wuser_reg <= temp_m_axi_wuser_reg;
    end

    if (store_axi_w_int_to_temp) begin
        temp_m_axi_wdata_reg <= m_axi_wdata_int;
        temp_m_axi_wstrb_reg <= m_axi_wstrb_int;
        temp_m_axi_wlast_reg <= m_axi_wlast_int;
        temp_m_axi_wuser_reg <= m_axi_wuser_int;
    end
end

endmodule

`resetall


// Content from axi_axil_adapter_wr.v
/*

Copyright (c) 2019 Alex Forencich

Permission is hereby granted, free of charge, to any person obtaining a copy
of this software and associated documentation files (the "Software"), to deal
in the Software without restriction, including without limitation the rights
to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
copies of the Software, and to permit persons to whom the Software is
furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in
all copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY
FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
THE SOFTWARE.

*/

// Language: Verilog 2001
/*
 * AXI4 to AXI4-Lite adapter (write)
 */
module axi_axil_adapter_wr #
(
    // Width of address bus in bits
    parameter ADDR_WIDTH = 32,
    // Width of input (slave) AXI interface data bus in bits
    parameter AXI_DATA_WIDTH = 32,
    // Width of input (slave) AXI interface wstrb (width of data bus in words)
    parameter AXI_STRB_WIDTH = (AXI_DATA_WIDTH/8),
    // Width of AXI ID signal
    parameter AXI_ID_WIDTH = 8,
    // Width of output (master) AXI lite interface data bus in bits
    parameter AXIL_DATA_WIDTH = 32,
    // Width of output (master) AXI lite interface wstrb (width of data bus in words)
    parameter AXIL_STRB_WIDTH = (AXIL_DATA_WIDTH/8),
    // When adapting to a wider bus, re-pack full-width burst instead of passing through narrow burst if possible
    parameter CONVERT_BURST = 1,
    // When adapting to a wider bus, re-pack all bursts instead of passing through narrow burst if possible
    parameter CONVERT_NARROW_BURST = 0
)
(
    input  wire                        clk,
    input  wire                        rst,

    /*
     * AXI slave interface
     */
    input  wire [AXI_ID_WIDTH-1:0]     s_axi_awid,
    input  wire [ADDR_WIDTH-1:0]       s_axi_awaddr,
    input  wire [7:0]                  s_axi_awlen,
    input  wire [2:0]                  s_axi_awsize,
    input  wire [1:0]                  s_axi_awburst,
    input  wire                        s_axi_awlock,
    input  wire [3:0]                  s_axi_awcache,
    input  wire [2:0]                  s_axi_awprot,
    input  wire                        s_axi_awvalid,
    output wire                        s_axi_awready,
    input  wire [AXI_DATA_WIDTH-1:0]   s_axi_wdata,
    input  wire [AXI_STRB_WIDTH-1:0]   s_axi_wstrb,
    input  wire                        s_axi_wlast,
    input  wire                        s_axi_wvalid,
    output wire                        s_axi_wready,
    output wire [AXI_ID_WIDTH-1:0]     s_axi_bid,
    output wire [1:0]                  s_axi_bresp,
    output wire                        s_axi_bvalid,
    input  wire                        s_axi_bready,

    /*
     * AXI lite master interface
     */
    output wire [ADDR_WIDTH-1:0]       m_axil_awaddr,
    output wire [2:0]                  m_axil_awprot,
    output wire                        m_axil_awvalid,
    input  wire                        m_axil_awready,
    output wire [AXIL_DATA_WIDTH-1:0]  m_axil_wdata,
    output wire [AXIL_STRB_WIDTH-1:0]  m_axil_wstrb,
    output wire                        m_axil_wvalid,
    input  wire                        m_axil_wready,
    input  wire [1:0]                  m_axil_bresp,
    input  wire                        m_axil_bvalid,
    output wire                        m_axil_bready
);

parameter AXI_ADDR_BIT_OFFSET = $clog2(AXI_STRB_WIDTH);
parameter AXIL_ADDR_BIT_OFFSET = $clog2(AXIL_STRB_WIDTH);
parameter AXI_WORD_WIDTH = AXI_STRB_WIDTH;
parameter AXIL_WORD_WIDTH = AXIL_STRB_WIDTH;
parameter AXI_WORD_SIZE = AXI_DATA_WIDTH/AXI_WORD_WIDTH;
parameter AXIL_WORD_SIZE = AXIL_DATA_WIDTH/AXIL_WORD_WIDTH;
parameter AXI_BURST_SIZE = $clog2(AXI_STRB_WIDTH);
parameter AXIL_BURST_SIZE = $clog2(AXIL_STRB_WIDTH);

// output bus is wider
parameter EXPAND = AXIL_STRB_WIDTH > AXI_STRB_WIDTH;
parameter DATA_WIDTH = EXPAND ? AXIL_DATA_WIDTH : AXI_DATA_WIDTH;
parameter STRB_WIDTH = EXPAND ? AXIL_STRB_WIDTH : AXI_STRB_WIDTH;
// required number of segments in wider bus
parameter SEGMENT_COUNT = EXPAND ? (AXIL_STRB_WIDTH / AXI_STRB_WIDTH) : (AXI_STRB_WIDTH / AXIL_STRB_WIDTH);
// data width and keep width per segment
parameter SEGMENT_DATA_WIDTH = DATA_WIDTH / SEGMENT_COUNT;
parameter SEGMENT_STRB_WIDTH = STRB_WIDTH / SEGMENT_COUNT;

localparam [1:0]
    STATE_IDLE = 2'd0,
    STATE_DATA = 2'd1,
    STATE_DATA_2 = 2'd2,
    STATE_RESP = 2'd3;

reg [1:0] state_reg = STATE_IDLE, state_next;

reg [AXI_ID_WIDTH-1:0] id_reg = {AXI_ID_WIDTH{1'b0}}, id_next;
reg [ADDR_WIDTH-1:0] addr_reg = {ADDR_WIDTH{1'b0}}, addr_next;
reg [DATA_WIDTH-1:0] data_reg = {DATA_WIDTH{1'b0}}, data_next;
reg [STRB_WIDTH-1:0] strb_reg = {STRB_WIDTH{1'b0}}, strb_next;
reg [7:0] burst_reg = 8'd0, burst_next;
reg [2:0] burst_size_reg = 3'd0, burst_size_next;
reg [2:0] master_burst_size_reg = 3'd0, master_burst_size_next;
reg burst_active_reg = 1'b0, burst_active_next;
reg convert_burst_reg = 1'b0, convert_burst_next;
reg first_transfer_reg = 1'b0, first_transfer_next;
reg last_segment_reg = 1'b0, last_segment_next;

reg s_axi_awready_reg = 1'b0, s_axi_awready_next;
reg s_axi_wready_reg = 1'b0, s_axi_wready_next;
reg [AXI_ID_WIDTH-1:0] s_axi_bid_reg = {AXI_ID_WIDTH{1'b0}}, s_axi_bid_next;
reg [1:0] s_axi_bresp_reg = 2'd0, s_axi_bresp_next;
reg s_axi_bvalid_reg = 1'b0, s_axi_bvalid_next;

reg [ADDR_WIDTH-1:0] m_axil_awaddr_reg = {ADDR_WIDTH{1'b0}}, m_axil_awaddr_next;
reg [2:0] m_axil_awprot_reg = 3'd0, m_axil_awprot_next;
reg m_axil_awvalid_reg = 1'b0, m_axil_awvalid_next;
reg [AXIL_DATA_WIDTH-1:0] m_axil_wdata_reg = {AXIL_DATA_WIDTH{1'b0}}, m_axil_wdata_next;
reg [AXIL_STRB_WIDTH-1:0] m_axil_wstrb_reg = {AXIL_STRB_WIDTH{1'b0}}, m_axil_wstrb_next;
reg m_axil_wvalid_reg = 1'b0, m_axil_wvalid_next;
reg m_axil_bready_reg = 1'b0, m_axil_bready_next;

assign s_axi_awready = s_axi_awready_reg;
assign s_axi_wready = s_axi_wready_reg;
assign s_axi_bid = s_axi_bid_reg;
assign s_axi_bresp = s_axi_bresp_reg;
assign s_axi_bvalid = s_axi_bvalid_reg;

assign m_axil_awaddr = m_axil_awaddr_reg;
//assign m_axil_awlen = m_axil_awlen_reg;
//assign m_axil_awsize = m_axil_awsize_reg;
//assign m_axil_awburst = m_axil_awburst_reg;
assign m_axil_awprot = m_axil_awprot_reg;
assign m_axil_awvalid = m_axil_awvalid_reg;
assign m_axil_wdata = m_axil_wdata_reg;
assign m_axil_wstrb = m_axil_wstrb_reg;
assign m_axil_wvalid = m_axil_wvalid_reg;
assign m_axil_bready = m_axil_bready_reg;

integer i;

always @* begin
    state_next = STATE_IDLE;

    id_next = id_reg;
    addr_next = addr_reg;
    data_next = data_reg;
    strb_next = strb_reg;
    burst_next = burst_reg;
    burst_size_next = burst_size_reg;
    master_burst_size_next = master_burst_size_reg;
    burst_active_next = burst_active_reg;
    convert_burst_next = convert_burst_reg;
    first_transfer_next = first_transfer_reg;
    last_segment_next = last_segment_reg;

    s_axi_awready_next = 1'b0;
    s_axi_wready_next = 1'b0;
    s_axi_bid_next = s_axi_bid_reg;
    s_axi_bresp_next = s_axi_bresp_reg;
    s_axi_bvalid_next = s_axi_bvalid_reg && !s_axi_bready;
    m_axil_awaddr_next = m_axil_awaddr_reg;
    m_axil_awprot_next = m_axil_awprot_reg;
    m_axil_awvalid_next = m_axil_awvalid_reg && !m_axil_awready;
    m_axil_wdata_next = m_axil_wdata_reg;
    m_axil_wstrb_next = m_axil_wstrb_reg;
    m_axil_wvalid_next = m_axil_wvalid_reg && !m_axil_wready;
    m_axil_bready_next = 1'b0;

    if (SEGMENT_COUNT == 1) begin
        // master output is same width; direct transfer with no splitting/merging
        case (state_reg)
            STATE_IDLE: begin
                // idle state; wait for new burst
                s_axi_awready_next = !m_axil_awvalid;
                first_transfer_next = 1'b1;

                if (s_axi_awready && s_axi_awvalid) begin
                    s_axi_awready_next = 1'b0;
                    id_next = s_axi_awid;
                    m_axil_awaddr_next = s_axi_awaddr;
                    addr_next = s_axi_awaddr;
                    burst_next = s_axi_awlen;
                    burst_size_next = s_axi_awsize;
                    burst_active_next = 1'b1;
                    m_axil_awprot_next = s_axi_awprot;
                    m_axil_awvalid_next = 1'b1;
                    s_axi_wready_next = !m_axil_wvalid;
                    state_next = STATE_DATA;
                end else begin
                    state_next = STATE_IDLE;
                end
            end
            STATE_DATA: begin
                // data state; transfer write data
                s_axi_wready_next = !m_axil_wvalid;

                if (s_axi_wready && s_axi_wvalid) begin
                    m_axil_wdata_next = s_axi_wdata;
                    m_axil_wstrb_next = s_axi_wstrb;
                    m_axil_wvalid_next = 1'b1;
                    burst_next = burst_reg - 1;
                    burst_active_next = burst_reg != 0;
                    addr_next = addr_reg + (1 << burst_size_reg);
                    s_axi_wready_next = 1'b0;
                    m_axil_bready_next = !s_axi_bvalid && !m_axil_awvalid;
                    state_next = STATE_RESP;
                end else begin
                    state_next = STATE_DATA;
                end
            end
            STATE_RESP: begin
                // resp state; transfer write response
                m_axil_bready_next = !s_axi_bvalid && !m_axil_awvalid;

                if (m_axil_bready && m_axil_bvalid) begin
                    m_axil_bready_next = 1'b0;
                    s_axi_bid_next = id_reg;
                    first_transfer_next = 1'b0;
                    if (first_transfer_reg || m_axil_bresp != 0) begin
                        s_axi_bresp_next = m_axil_bresp;
                    end
                    if (burst_active_reg) begin
                        // burst on slave interface still active; start new AXI lite write
                        m_axil_awaddr_next = addr_reg;
                        m_axil_awvalid_next = 1'b1;
                        s_axi_wready_next = !m_axil_wvalid;
                        state_next = STATE_DATA;
                    end else begin
                        // burst on slave interface finished; return to idle
                        s_axi_bvalid_next = 1'b1;
                        s_axi_awready_next = !m_axil_awvalid;
                        state_next = STATE_IDLE;
                    end
                end else begin
                    state_next = STATE_RESP;
                end
            end
        endcase
    end else if (EXPAND) begin
        // master output is wider; merge writes
        case (state_reg)
            STATE_IDLE: begin
                // idle state; wait for new burst
                s_axi_awready_next = !m_axil_awvalid;

                first_transfer_next = 1'b1;

                data_next = {DATA_WIDTH{1'b0}};
                strb_next = {STRB_WIDTH{1'b0}};

                if (s_axi_awready && s_axi_awvalid) begin
                    s_axi_awready_next = 1'b0;
                    id_next = s_axi_awid;
                    m_axil_awaddr_next = s_axi_awaddr;
                    addr_next = s_axi_awaddr;
                    burst_next = s_axi_awlen;
                    burst_size_next = s_axi_awsize;
                    if (CONVERT_BURST && s_axi_awcache[1] && (CONVERT_NARROW_BURST || s_axi_awsize == AXI_BURST_SIZE)) begin
                        // merge writes
                        // require CONVERT_BURST and awcache[1] set
                        convert_burst_next = 1'b1;
                        master_burst_size_next = AXIL_BURST_SIZE;
                        state_next = STATE_DATA_2;
                    end else begin
                        // output narrow burst
                        convert_burst_next = 1'b0;
                        master_burst_size_next = s_axi_awsize;
                        state_next = STATE_DATA;
                    end
                    m_axil_awprot_next = s_axi_awprot;
                    m_axil_awvalid_next = 1'b1;
                    s_axi_wready_next = !m_axil_wvalid;
                end else begin
                    state_next = STATE_IDLE;
                end
            end
            STATE_DATA: begin
                // data state; transfer write data
                s_axi_wready_next = !m_axil_wvalid || m_axil_wready;

                if (s_axi_wready && s_axi_wvalid) begin
                    m_axil_wdata_next = {(AXIL_WORD_WIDTH/AXI_WORD_WIDTH){s_axi_wdata}};
                    m_axil_wstrb_next = s_axi_wstrb << (addr_reg[AXIL_ADDR_BIT_OFFSET-1:AXI_ADDR_BIT_OFFSET] * AXI_STRB_WIDTH);
                    m_axil_wvalid_next = 1'b1;
                    burst_next = burst_reg - 1;
                    burst_active_next = burst_reg != 0;
                    addr_next = addr_reg + (1 << burst_size_reg);
                    s_axi_wready_next = 1'b0;
                    m_axil_bready_next = !s_axi_bvalid && !m_axil_awvalid;
                    state_next = STATE_RESP;
                end else begin
                    state_next = STATE_DATA;
                end
            end
            STATE_DATA_2: begin
                s_axi_wready_next = !m_axil_wvalid;

                if (s_axi_wready && s_axi_wvalid) begin
                    if (CONVERT_NARROW_BURST) begin
                        for (i = 0; i < AXI_WORD_WIDTH; i = i + 1) begin
                            if (s_axi_wstrb[i]) begin
                                data_next[addr_reg[AXIL_ADDR_BIT_OFFSET-1:AXI_ADDR_BIT_OFFSET]*SEGMENT_DATA_WIDTH+i*AXIL_WORD_SIZE +: AXIL_WORD_SIZE] = s_axi_wdata[i*AXIL_WORD_SIZE +: AXIL_WORD_SIZE];
                                strb_next[addr_reg[AXIL_ADDR_BIT_OFFSET-1:AXI_ADDR_BIT_OFFSET]*SEGMENT_STRB_WIDTH+i] = 1'b1;
                            end
                        end
                    end else begin
                        data_next[addr_reg[AXIL_ADDR_BIT_OFFSET-1:AXI_ADDR_BIT_OFFSET]*SEGMENT_DATA_WIDTH +: SEGMENT_DATA_WIDTH] = s_axi_wdata;
                        strb_next[addr_reg[AXIL_ADDR_BIT_OFFSET-1:AXI_ADDR_BIT_OFFSET]*SEGMENT_STRB_WIDTH +: SEGMENT_STRB_WIDTH] = s_axi_wstrb;
                    end
                    m_axil_wdata_next = data_next;
                    m_axil_wstrb_next = strb_next;
                    burst_next = burst_reg - 1;
                    burst_active_next = burst_reg != 0;
                    addr_next = addr_reg + (1 << burst_size_reg);
                    if (burst_reg == 0 || addr_next[master_burst_size_reg] != addr_reg[master_burst_size_reg]) begin
                        data_next = {DATA_WIDTH{1'b0}};
                        strb_next = {STRB_WIDTH{1'b0}};
                        m_axil_wvalid_next = 1'b1;
                        s_axi_wready_next = 1'b0;
                        m_axil_bready_next = !s_axi_bvalid && !m_axil_awvalid;
                        state_next = STATE_RESP;
                    end else begin
                        state_next = STATE_DATA_2;
                    end
                end else begin
                    state_next = STATE_DATA_2;
                end
            end
            STATE_RESP: begin
                // resp state; transfer write response
                m_axil_bready_next = !s_axi_bvalid && !m_axil_awvalid;

                if (m_axil_bready && m_axil_bvalid) begin
                    m_axil_bready_next = 1'b0;
                    s_axi_bid_next = id_reg;
                    first_transfer_next = 1'b0;
                    if (first_transfer_reg || m_axil_bresp != 0) begin
                        s_axi_bresp_next = m_axil_bresp;
                    end
                    if (burst_active_reg) begin
                        // burst on slave interface still active; start new AXI lite write
                        m_axil_awaddr_next = addr_reg;
                        m_axil_awvalid_next = 1'b1;
                        s_axi_wready_next = !m_axil_wvalid || m_axil_wready;
                        if (convert_burst_reg) begin
                            state_next = STATE_DATA_2;
                        end else begin
                            state_next = STATE_DATA;
                        end
                    end else begin
                        // burst on slave interface finished; return to idle
                        s_axi_bvalid_next = 1'b1;
                        s_axi_awready_next = !m_axil_awvalid;
                        state_next = STATE_IDLE;
                    end
                end else begin
                    state_next = STATE_RESP;
                end
            end
        endcase
    end else begin
        // master output is narrower; split writes, and possibly split burst
        case (state_reg)
            STATE_IDLE: begin
                // idle state; wait for new burst
                s_axi_awready_next = !m_axil_awvalid;

                first_transfer_next = 1'b1;

                if (s_axi_awready && s_axi_awvalid) begin
                    s_axi_awready_next = 1'b0;
                    id_next = s_axi_awid;
                    m_axil_awaddr_next = s_axi_awaddr;
                    addr_next = s_axi_awaddr;
                    burst_next = s_axi_awlen;
                    burst_size_next = s_axi_awsize;
                    burst_active_next = 1'b1;
                    if (s_axi_awsize > AXIL_BURST_SIZE) begin
                        // need to adjust burst size
                        master_burst_size_next = AXIL_BURST_SIZE;
                    end else begin
                        // pass through narrow (enough) burst
                        master_burst_size_next = s_axi_awsize;
                    end
                    m_axil_awprot_next = s_axi_awprot;
                    m_axil_awvalid_next = 1'b1;
                    s_axi_wready_next = !m_axil_wvalid;
                    state_next = STATE_DATA;
                end else begin
                    state_next = STATE_IDLE;
                end
            end
            STATE_DATA: begin
                s_axi_wready_next = !m_axil_wvalid;

                if (s_axi_wready && s_axi_wvalid) begin
                    data_next = s_axi_wdata;
                    strb_next = s_axi_wstrb;
                    m_axil_wdata_next = s_axi_wdata >> (addr_reg[AXI_ADDR_BIT_OFFSET-1:AXIL_ADDR_BIT_OFFSET] * AXIL_DATA_WIDTH);
                    m_axil_wstrb_next = s_axi_wstrb >> (addr_reg[AXI_ADDR_BIT_OFFSET-1:AXIL_ADDR_BIT_OFFSET] * AXIL_STRB_WIDTH);
                    m_axil_wvalid_next = 1'b1;
                    burst_next = burst_reg - 1;
                    burst_active_next = burst_reg != 0;
                    addr_next = (addr_reg + (1 << master_burst_size_reg)) & ({ADDR_WIDTH{1'b1}} << master_burst_size_reg);
                    last_segment_next = addr_next[burst_size_reg] != addr_reg[burst_size_reg];
                    s_axi_wready_next = 1'b0;
                    m_axil_bready_next = !s_axi_bvalid && !m_axil_awvalid;
                    state_next = STATE_RESP;
                end else begin
                    state_next = STATE_DATA;
                end
            end
            STATE_DATA_2: begin
                s_axi_wready_next = 1'b0;

                if (!m_axil_wvalid || m_axil_wready) begin
                    m_axil_wdata_next = data_reg >> (addr_reg[AXI_ADDR_BIT_OFFSET-1:AXIL_ADDR_BIT_OFFSET] * AXIL_DATA_WIDTH);
                    m_axil_wstrb_next = strb_reg >> (addr_reg[AXI_ADDR_BIT_OFFSET-1:AXIL_ADDR_BIT_OFFSET] * AXIL_STRB_WIDTH);
                    m_axil_wvalid_next = 1'b1;
                    addr_next = (addr_reg + (1 << master_burst_size_reg)) & ({ADDR_WIDTH{1'b1}} << master_burst_size_reg);
                    last_segment_next = addr_next[burst_size_reg] != addr_reg[burst_size_reg];
                    s_axi_wready_next = 1'b0;
                    m_axil_bready_next = !s_axi_bvalid && !m_axil_awvalid;
                    state_next = STATE_RESP;
                end else begin
                    state_next = STATE_DATA_2;
                end
            end
            STATE_RESP: begin
                // resp state; transfer write response
                m_axil_bready_next = !s_axi_bvalid && !m_axil_awvalid;

                if (m_axil_bready && m_axil_bvalid) begin
                    first_transfer_next = 1'b0;
                    m_axil_awaddr_next = addr_reg;
                    m_axil_bready_next = 1'b0;
                    s_axi_bid_next = id_reg;
                    if (first_transfer_reg || m_axil_bresp != 0) begin
                        s_axi_bresp_next = m_axil_bresp;
                    end
                    if (burst_active_reg || !last_segment_reg) begin
                        // burst on slave interface still active; start new burst
                        m_axil_awvalid_next = 1'b1;
                        if (last_segment_reg) begin
                            s_axi_wready_next = !m_axil_wvalid;
                            state_next = STATE_DATA;
                        end else begin
                            s_axi_wready_next = 1'b0;
                            state_next = STATE_DATA_2;
                        end
                    end else begin
                        // burst on slave interface finished; return to idle
                        s_axi_bvalid_next = 1'b1;
                        s_axi_awready_next = !m_axil_awvalid;
                        state_next = STATE_IDLE;
                    end
                end else begin
                    state_next = STATE_RESP;
                end
            end
        endcase
    end
end

always @(posedge clk) begin
    state_reg <= state_next;

    id_reg <= id_next;
    addr_reg <= addr_next;
    data_reg <= data_next;
    strb_reg <= strb_next;
    burst_reg <= burst_next;
    burst_size_reg <= burst_size_next;
    master_burst_size_reg <= master_burst_size_next;
    burst_active_reg <= burst_active_next;
    convert_burst_reg <= convert_burst_next;
    first_transfer_reg <= first_transfer_next;
    last_segment_reg <= last_segment_next;

    s_axi_awready_reg <= s_axi_awready_next;
    s_axi_wready_reg <= s_axi_wready_next;
    s_axi_bid_reg <= s_axi_bid_next;
    s_axi_bresp_reg <= s_axi_bresp_next;
    s_axi_bvalid_reg <= s_axi_bvalid_next;

    m_axil_awaddr_reg <= m_axil_awaddr_next;
    m_axil_awprot_reg <= m_axil_awprot_next;
    m_axil_awvalid_reg <= m_axil_awvalid_next;
    m_axil_wdata_reg <= m_axil_wdata_next;
    m_axil_wstrb_reg <= m_axil_wstrb_next;
    m_axil_wvalid_reg <= m_axil_wvalid_next;
    m_axil_bready_reg <= m_axil_bready_next;

    if (rst) begin
        state_reg <= STATE_IDLE;

        s_axi_awready_reg <= 1'b0;
        s_axi_wready_reg <= 1'b0;
        s_axi_bvalid_reg <= 1'b0;

        m_axil_awvalid_reg <= 1'b0;
        m_axil_wvalid_reg <= 1'b0;
        m_axil_bready_reg <= 1'b0;
    end
end

endmodule

`resetall


// Content from priority_encoder.v
/*

Copyright (c) 2014-2021 Alex Forencich

Permission is hereby granted, free of charge, to any person obtaining a copy
of this software and associated documentation files (the "Software"), to deal
in the Software without restriction, including without limitation the rights
to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
copies of the Software, and to permit persons to whom the Software is
furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in
all copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY
FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
THE SOFTWARE.

*/

// Language: Verilog 2001

`resetall
`timescale 1ns / 1ps
`default_nettype none

/*
 * Priority encoder module
 */
module priority_encoder #
(
    parameter WIDTH = 4,
    // LSB priority selection
    parameter LSB_HIGH_PRIORITY = 0
)
(
    input  wire [WIDTH-1:0]         input_unencoded,
    output wire                     output_valid,
    output wire [$clog2(WIDTH)-1:0] output_encoded,
    output wire [WIDTH-1:0]         output_unencoded
);

parameter LEVELS = WIDTH > 2 ? $clog2(WIDTH) : 1;
parameter W = 2**LEVELS;

// pad input to even power of two
wire [W-1:0] input_padded = {{W-WIDTH{1'b0}}, input_unencoded};

wire [W/2-1:0] stage_valid[LEVELS-1:0];
wire [W/2-1:0] stage_enc[LEVELS-1:0];

generate
    genvar l, n;

    // process input bits; generate valid bit and encoded bit for each pair
    for (n = 0; n < W/2; n = n + 1) begin : loop_in
        assign stage_valid[0][n] = |input_padded[n*2+1:n*2];
        if (LSB_HIGH_PRIORITY) begin
            // bit 0 is highest priority
            assign stage_enc[0][n] = !input_padded[n*2+0];
        end else begin
            // bit 0 is lowest priority
            assign stage_enc[0][n] = input_padded[n*2+1];
        end
    end

    // compress down to single valid bit and encoded bus
    for (l = 1; l < LEVELS; l = l + 1) begin : loop_levels
        for (n = 0; n < W/(2*2**l); n = n + 1) begin : loop_compress
            assign stage_valid[l][n] = |stage_valid[l-1][n*2+1:n*2];
            if (LSB_HIGH_PRIORITY) begin
                // bit 0 is highest priority
                assign stage_enc[l][(n+1)*(l+1)-1:n*(l+1)] = stage_valid[l-1][n*2+0] ? {1'b0, stage_enc[l-1][(n*2+1)*l-1:(n*2+0)*l]} : {1'b1, stage_enc[l-1][(n*2+2)*l-1:(n*2+1)*l]};
            end else begin
                // bit 0 is lowest priority
                assign stage_enc[l][(n+1)*(l+1)-1:n*(l+1)] = stage_valid[l-1][n*2+1] ? {1'b1, stage_enc[l-1][(n*2+2)*l-1:(n*2+1)*l]} : {1'b0, stage_enc[l-1][(n*2+1)*l-1:(n*2+0)*l]};
            end
        end
    end
endgenerate

assign output_valid = stage_valid[LEVELS-1];
assign output_encoded = stage_enc[LEVELS-1];
assign output_unencoded = 1 << output_encoded;

endmodule

`resetall


// Content from axil_interconnect_wrap_1x2.v
/*

Copyright (c) 2020 Alex Forencich

Permission is hereby granted, free of charge, to any person obtaining a copy
of this software and associated documentation files (the "Software"), to deal
in the Software without restriction, including without limitation the rights
to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
copies of the Software, and to permit persons to whom the Software is
furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in
all copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY
FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
THE SOFTWARE.

*/

// Language: Verilog 2001

/*
 * AXI4 lite 1x2 interconnect (wrapper)
 */
module axil_interconnect_wrap_1x2 #
(
    parameter DATA_WIDTH = 32,
    parameter ADDR_WIDTH = 16,
    parameter STRB_WIDTH = (DATA_WIDTH/8),
    parameter M_REGIONS = 1,
    parameter M00_BASE_ADDR = 0,
    parameter M00_ADDR_WIDTH = {M_REGIONS{32'd24}},
    parameter M00_CONNECT_READ = 1'b1,
    parameter M00_CONNECT_WRITE = 1'b1,
    parameter M00_SECURE = 1'b0,
    parameter M01_BASE_ADDR = 0,
    parameter M01_ADDR_WIDTH = {M_REGIONS{32'd24}},
    parameter M01_CONNECT_READ = 1'b1,
    parameter M01_CONNECT_WRITE = 1'b1,
    parameter M01_SECURE = 1'b0
)
(
    input  wire                     clk,
    input  wire                     rst,

    /*
     * AXI lite slave interfaces
     */
    input  wire [ADDR_WIDTH-1:0]    s00_axil_awaddr,
    input  wire [2:0]               s00_axil_awprot,
    input  wire                     s00_axil_awvalid,
    output wire                     s00_axil_awready,
    input  wire [DATA_WIDTH-1:0]    s00_axil_wdata,
    input  wire [STRB_WIDTH-1:0]    s00_axil_wstrb,
    input  wire                     s00_axil_wvalid,
    output wire                     s00_axil_wready,
    output wire [1:0]               s00_axil_bresp,
    output wire                     s00_axil_bvalid,
    input  wire                     s00_axil_bready,
    input  wire [ADDR_WIDTH-1:0]    s00_axil_araddr,
    input  wire [2:0]               s00_axil_arprot,
    input  wire                     s00_axil_arvalid,
    output wire                     s00_axil_arready,
    output wire [DATA_WIDTH-1:0]    s00_axil_rdata,
    output wire [1:0]               s00_axil_rresp,
    output wire                     s00_axil_rvalid,
    input  wire                     s00_axil_rready,

    /*
     * AXI lite master interfaces
     */
    output wire [ADDR_WIDTH-1:0]    m00_axil_awaddr,
    output wire [2:0]               m00_axil_awprot,
    output wire                     m00_axil_awvalid,
    input  wire                     m00_axil_awready,
    output wire [DATA_WIDTH-1:0]    m00_axil_wdata,
    output wire [STRB_WIDTH-1:0]    m00_axil_wstrb,
    output wire                     m00_axil_wvalid,
    input  wire                     m00_axil_wready,
    input  wire [1:0]               m00_axil_bresp,
    input  wire                     m00_axil_bvalid,
    output wire                     m00_axil_bready,
    output wire [ADDR_WIDTH-1:0]    m00_axil_araddr,
    output wire [2:0]               m00_axil_arprot,
    output wire                     m00_axil_arvalid,
    input  wire                     m00_axil_arready,
    input  wire [DATA_WIDTH-1:0]    m00_axil_rdata,
    input  wire [1:0]               m00_axil_rresp,
    input  wire                     m00_axil_rvalid,
    output wire                     m00_axil_rready,

    output wire [ADDR_WIDTH-1:0]    m01_axil_awaddr,
    output wire [2:0]               m01_axil_awprot,
    output wire                     m01_axil_awvalid,
    input  wire                     m01_axil_awready,
    output wire [DATA_WIDTH-1:0]    m01_axil_wdata,
    output wire [STRB_WIDTH-1:0]    m01_axil_wstrb,
    output wire                     m01_axil_wvalid,
    input  wire                     m01_axil_wready,
    input  wire [1:0]               m01_axil_bresp,
    input  wire                     m01_axil_bvalid,
    output wire                     m01_axil_bready,
    output wire [ADDR_WIDTH-1:0]    m01_axil_araddr,
    output wire [2:0]               m01_axil_arprot,
    output wire                     m01_axil_arvalid,
    input  wire                     m01_axil_arready,
    input  wire [DATA_WIDTH-1:0]    m01_axil_rdata,
    input  wire [1:0]               m01_axil_rresp,
    input  wire                     m01_axil_rvalid,
    output wire                     m01_axil_rready
);

localparam S_COUNT = 1;
localparam M_COUNT = 2;

// parameter sizing helpers
function [ADDR_WIDTH*M_REGIONS-1:0] w_a_r(input [ADDR_WIDTH*M_REGIONS-1:0] val);
    w_a_r = val;
endfunction

function [32*M_REGIONS-1:0] w_32_r(input [32*M_REGIONS-1:0] val);
    w_32_r = val;
endfunction

function [S_COUNT-1:0] w_s(input [S_COUNT-1:0] val);
    w_s = val;
endfunction

function w_1(input val);
    w_1 = val;
endfunction

axil_interconnect #(
    .S_COUNT(S_COUNT),
    .M_COUNT(M_COUNT),
    .DATA_WIDTH(DATA_WIDTH),
    .ADDR_WIDTH(ADDR_WIDTH),
    .STRB_WIDTH(STRB_WIDTH),
    .M_REGIONS(M_REGIONS),
    .M_BASE_ADDR({ w_a_r(M01_BASE_ADDR), w_a_r(M00_BASE_ADDR) }),
    .M_ADDR_WIDTH({ w_32_r(M01_ADDR_WIDTH), w_32_r(M00_ADDR_WIDTH) }),
    .M_CONNECT_READ({ w_s(M01_CONNECT_READ), w_s(M00_CONNECT_READ) }),
    .M_CONNECT_WRITE({ w_s(M01_CONNECT_WRITE), w_s(M00_CONNECT_WRITE) }),
    .M_SECURE({ w_1(M01_SECURE), w_1(M00_SECURE) })
)
axil_interconnect_inst (
    .clk(clk),
    .rst(rst),
    .s_axil_awaddr({ s00_axil_awaddr }),
    .s_axil_awprot({ s00_axil_awprot }),
    .s_axil_awvalid({ s00_axil_awvalid }),
    .s_axil_awready({ s00_axil_awready }),
    .s_axil_wdata({ s00_axil_wdata }),
    .s_axil_wstrb({ s00_axil_wstrb }),
    .s_axil_wvalid({ s00_axil_wvalid }),
    .s_axil_wready({ s00_axil_wready }),
    .s_axil_bresp({ s00_axil_bresp }),
    .s_axil_bvalid({ s00_axil_bvalid }),
    .s_axil_bready({ s00_axil_bready }),
    .s_axil_araddr({ s00_axil_araddr }),
    .s_axil_arprot({ s00_axil_arprot }),
    .s_axil_arvalid({ s00_axil_arvalid }),
    .s_axil_arready({ s00_axil_arready }),
    .s_axil_rdata({ s00_axil_rdata }),
    .s_axil_rresp({ s00_axil_rresp }),
    .s_axil_rvalid({ s00_axil_rvalid }),
    .s_axil_rready({ s00_axil_rready }),
    .m_axil_awaddr({ m01_axil_awaddr, m00_axil_awaddr }),
    .m_axil_awprot({ m01_axil_awprot, m00_axil_awprot }),
    .m_axil_awvalid({ m01_axil_awvalid, m00_axil_awvalid }),
    .m_axil_awready({ m01_axil_awready, m00_axil_awready }),
    .m_axil_wdata({ m01_axil_wdata, m00_axil_wdata }),
    .m_axil_wstrb({ m01_axil_wstrb, m00_axil_wstrb }),
    .m_axil_wvalid({ m01_axil_wvalid, m00_axil_wvalid }),
    .m_axil_wready({ m01_axil_wready, m00_axil_wready }),
    .m_axil_bresp({ m01_axil_bresp, m00_axil_bresp }),
    .m_axil_bvalid({ m01_axil_bvalid, m00_axil_bvalid }),
    .m_axil_bready({ m01_axil_bready, m00_axil_bready }),
    .m_axil_araddr({ m01_axil_araddr, m00_axil_araddr }),
    .m_axil_arprot({ m01_axil_arprot, m00_axil_arprot }),
    .m_axil_arvalid({ m01_axil_arvalid, m00_axil_arvalid }),
    .m_axil_arready({ m01_axil_arready, m00_axil_arready }),
    .m_axil_rdata({ m01_axil_rdata, m00_axil_rdata }),
    .m_axil_rresp({ m01_axil_rresp, m00_axil_rresp }),
    .m_axil_rvalid({ m01_axil_rvalid, m00_axil_rvalid }),
    .m_axil_rready({ m01_axil_rready, m00_axil_rready })
);

endmodule

`resetall


// Content from axi_axil_adapter_rd.v
/*

Copyright (c) 2019 Alex Forencich

Permission is hereby granted, free of charge, to any person obtaining a copy
of this software and associated documentation files (the "Software"), to deal
in the Software without restriction, including without limitation the rights
to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
copies of the Software, and to permit persons to whom the Software is
furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in
all copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY
FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
THE SOFTWARE.

*/

// Language: Verilog 2001

/*
 * AXI4 to AXI4-Lite adapter (read)
 */
module axi_axil_adapter_rd #
(
    // Width of address bus in bits
    parameter ADDR_WIDTH = 32,
    // Width of input (slave) AXI interface data bus in bits
    parameter AXI_DATA_WIDTH = 32,
    // Width of input (slave) AXI interface wstrb (width of data bus in words)
    parameter AXI_STRB_WIDTH = (AXI_DATA_WIDTH/8),
    // Width of AXI ID signal
    parameter AXI_ID_WIDTH = 8,
    // Width of output (master) AXI lite interface data bus in bits
    parameter AXIL_DATA_WIDTH = 32,
    // Width of output (master) AXI lite interface wstrb (width of data bus in words)
    parameter AXIL_STRB_WIDTH = (AXIL_DATA_WIDTH/8),
    // When adapting to a wider bus, re-pack full-width burst instead of passing through narrow burst if possible
    parameter CONVERT_BURST = 1,
    // When adapting to a wider bus, re-pack all bursts instead of passing through narrow burst if possible
    parameter CONVERT_NARROW_BURST = 0
)
(
    input  wire                        clk,
    input  wire                        rst,

    /*
     * AXI slave interface
     */
    input  wire [AXI_ID_WIDTH-1:0]     s_axi_arid,
    input  wire [ADDR_WIDTH-1:0]       s_axi_araddr,
    input  wire [7:0]                  s_axi_arlen,
    input  wire [2:0]                  s_axi_arsize,
    input  wire [1:0]                  s_axi_arburst,
    input  wire                        s_axi_arlock,
    input  wire [3:0]                  s_axi_arcache,
    input  wire [2:0]                  s_axi_arprot,
    input  wire                        s_axi_arvalid,
    output wire                        s_axi_arready,
    output wire [AXI_ID_WIDTH-1:0]     s_axi_rid,
    output wire [AXI_DATA_WIDTH-1:0]   s_axi_rdata,
    output wire [1:0]                  s_axi_rresp,
    output wire                        s_axi_rlast,
    output wire                        s_axi_rvalid,
    input  wire                        s_axi_rready,

    /*
     * AXI lite master interface
     */
    output wire [ADDR_WIDTH-1:0]       m_axil_araddr,
    output wire [2:0]                  m_axil_arprot,
    output wire                        m_axil_arvalid,
    input  wire                        m_axil_arready,
    input  wire [AXIL_DATA_WIDTH-1:0]  m_axil_rdata,
    input  wire [1:0]                  m_axil_rresp,
    input  wire                        m_axil_rvalid,
    output wire                        m_axil_rready
);

parameter AXI_ADDR_BIT_OFFSET = $clog2(AXI_STRB_WIDTH);
parameter AXIL_ADDR_BIT_OFFSET = $clog2(AXIL_STRB_WIDTH);
parameter AXI_WORD_WIDTH = AXI_STRB_WIDTH;
parameter AXIL_WORD_WIDTH = AXIL_STRB_WIDTH;
parameter AXI_WORD_SIZE = AXI_DATA_WIDTH/AXI_WORD_WIDTH;
parameter AXIL_WORD_SIZE = AXIL_DATA_WIDTH/AXIL_WORD_WIDTH;
parameter AXI_BURST_SIZE = $clog2(AXI_STRB_WIDTH);
parameter AXIL_BURST_SIZE = $clog2(AXIL_STRB_WIDTH);

// output bus is wider
parameter EXPAND = AXIL_STRB_WIDTH > AXI_STRB_WIDTH;
parameter DATA_WIDTH = EXPAND ? AXIL_DATA_WIDTH : AXI_DATA_WIDTH;
parameter STRB_WIDTH = EXPAND ? AXIL_STRB_WIDTH : AXI_STRB_WIDTH;
// required number of segments in wider bus
parameter SEGMENT_COUNT = EXPAND ? (AXIL_STRB_WIDTH / AXI_STRB_WIDTH) : (AXI_STRB_WIDTH / AXIL_STRB_WIDTH);
// data width and keep width per segment
parameter SEGMENT_DATA_WIDTH = DATA_WIDTH / SEGMENT_COUNT;
parameter SEGMENT_STRB_WIDTH = STRB_WIDTH / SEGMENT_COUNT;



localparam [1:0]
    STATE_IDLE = 2'd0,
    STATE_DATA = 2'd1,
    STATE_DATA_READ = 2'd2,
    STATE_DATA_SPLIT = 2'd3;

reg [1:0] state_reg = STATE_IDLE, state_next;

reg [AXI_ID_WIDTH-1:0] id_reg = {AXI_ID_WIDTH{1'b0}}, id_next;
reg [ADDR_WIDTH-1:0] addr_reg = {ADDR_WIDTH{1'b0}}, addr_next;
reg [DATA_WIDTH-1:0] data_reg = {DATA_WIDTH{1'b0}}, data_next;
reg [1:0] resp_reg = 2'd0, resp_next;
reg [7:0] burst_reg = 8'd0, burst_next;
reg [2:0] burst_size_reg = 3'd0, burst_size_next;
reg [7:0] master_burst_reg = 8'd0, master_burst_next;
reg [2:0] master_burst_size_reg = 3'd0, master_burst_size_next;

reg s_axi_arready_reg = 1'b0, s_axi_arready_next;
reg [AXI_ID_WIDTH-1:0] s_axi_rid_reg = {AXI_ID_WIDTH{1'b0}}, s_axi_rid_next;
reg [AXI_DATA_WIDTH-1:0] s_axi_rdata_reg = {AXI_DATA_WIDTH{1'b0}}, s_axi_rdata_next;
reg [1:0] s_axi_rresp_reg = 2'd0, s_axi_rresp_next;
reg s_axi_rlast_reg = 1'b0, s_axi_rlast_next;
reg s_axi_rvalid_reg = 1'b0, s_axi_rvalid_next;

reg [ADDR_WIDTH-1:0] m_axil_araddr_reg = {ADDR_WIDTH{1'b0}}, m_axil_araddr_next;
reg [2:0] m_axil_arprot_reg = 3'd0, m_axil_arprot_next;
reg m_axil_arvalid_reg = 1'b0, m_axil_arvalid_next;
reg m_axil_rready_reg = 1'b0, m_axil_rready_next;

assign s_axi_arready = s_axi_arready_reg;
assign s_axi_rid = s_axi_rid_reg;
assign s_axi_rdata = s_axi_rdata_reg;
assign s_axi_rresp = s_axi_rresp_reg;
assign s_axi_rlast = s_axi_rlast_reg;
assign s_axi_rvalid = s_axi_rvalid_reg;

assign m_axil_araddr = m_axil_araddr_reg;
assign m_axil_arprot = m_axil_arprot_reg;
assign m_axil_arvalid = m_axil_arvalid_reg;
assign m_axil_rready = m_axil_rready_reg;

always @* begin
    state_next = STATE_IDLE;

    id_next = id_reg;
    addr_next = addr_reg;
    data_next = data_reg;
    resp_next = resp_reg;
    burst_next = burst_reg;
    burst_size_next = burst_size_reg;
    master_burst_next = master_burst_reg;
    master_burst_size_next = master_burst_size_reg;

    s_axi_arready_next = 1'b0;
    s_axi_rid_next = s_axi_rid_reg;
    s_axi_rdata_next = s_axi_rdata_reg;
    s_axi_rresp_next = s_axi_rresp_reg;
    s_axi_rlast_next = s_axi_rlast_reg;
    s_axi_rvalid_next = s_axi_rvalid_reg && !s_axi_rready;
    m_axil_araddr_next = m_axil_araddr_reg;
    m_axil_arprot_next = m_axil_arprot_reg;
    m_axil_arvalid_next = m_axil_arvalid_reg && !m_axil_arready;
    m_axil_rready_next = 1'b0;

    if (SEGMENT_COUNT == 1) begin
        // master output is same width; direct transfer with no splitting/merging
        case (state_reg)
            STATE_IDLE: begin
                // idle state; wait for new burst
                s_axi_arready_next = !m_axil_arvalid;

                if (s_axi_arready && s_axi_arvalid) begin
                    s_axi_arready_next = 1'b0;
                    id_next = s_axi_arid;
                    m_axil_araddr_next = s_axi_araddr;
                    addr_next = s_axi_araddr;
                    burst_next = s_axi_arlen;
                    burst_size_next = s_axi_arsize;
                    m_axil_arprot_next = s_axi_arprot;
                    m_axil_arvalid_next = 1'b1;
                    m_axil_rready_next = 1'b0;
                    state_next = STATE_DATA;
                end else begin
                    state_next = STATE_IDLE;
                end
            end
            STATE_DATA: begin
                // data state; transfer read data
                m_axil_rready_next = !s_axi_rvalid && !m_axil_arvalid;

                if (m_axil_rready && m_axil_rvalid) begin
                    s_axi_rid_next = id_reg;
                    s_axi_rdata_next = m_axil_rdata;
                    s_axi_rresp_next = m_axil_rresp;
                    s_axi_rlast_next = 1'b0;
                    s_axi_rvalid_next = 1'b1;
                    burst_next = burst_reg - 1;
                    addr_next = addr_reg + (1 << burst_size_reg);
                    if (burst_reg == 0) begin
                        // last data word, return to idle
                        m_axil_rready_next = 1'b0;
                        s_axi_rlast_next = 1'b1;
                        s_axi_arready_next = !m_axil_arvalid;
                        state_next = STATE_IDLE;
                    end else begin
                        // start new AXI lite read
                        m_axil_araddr_next = addr_next;
                        m_axil_arvalid_next = 1'b1;
                        m_axil_rready_next = 1'b0;
                        state_next = STATE_DATA;
                    end
                end else begin
                    state_next = STATE_DATA;
                end
            end
        endcase
    end else if (EXPAND) begin
        // master output is wider; split reads
        case (state_reg)
            STATE_IDLE: begin
                // idle state; wait for new burst
                s_axi_arready_next = !m_axil_arvalid;

                if (s_axi_arready && s_axi_arvalid) begin
                    s_axi_arready_next = 1'b0;
                    id_next = s_axi_arid;
                    m_axil_araddr_next = s_axi_araddr;
                    addr_next = s_axi_araddr;
                    burst_next = s_axi_arlen;
                    burst_size_next = s_axi_arsize;
                    if (CONVERT_BURST && s_axi_arcache[1] && (CONVERT_NARROW_BURST || s_axi_arsize == AXI_BURST_SIZE)) begin
                        // split reads
                        // require CONVERT_BURST and arcache[1] set
                        master_burst_size_next = AXIL_BURST_SIZE;
                        state_next = STATE_DATA_READ;
                    end else begin
                        // output narrow burst
                        master_burst_size_next = s_axi_arsize;
                        state_next = STATE_DATA;
                    end
                    m_axil_arprot_next = s_axi_arprot;
                    m_axil_arvalid_next = 1'b1;
                    m_axil_rready_next = 1'b0;
                end else begin
                    state_next = STATE_IDLE;
                end
            end
            STATE_DATA: begin
                m_axil_rready_next = !s_axi_rvalid && !m_axil_arvalid;

                if (m_axil_rready && m_axil_rvalid) begin
                    s_axi_rid_next = id_reg;
                    s_axi_rdata_next = m_axil_rdata >> (addr_reg[AXIL_ADDR_BIT_OFFSET-1:AXI_ADDR_BIT_OFFSET] * AXI_DATA_WIDTH);
                    s_axi_rresp_next = m_axil_rresp;
                    s_axi_rlast_next = 1'b0;
                    s_axi_rvalid_next = 1'b1;
                    burst_next = burst_reg - 1;
                    addr_next = addr_reg + (1 << burst_size_reg);
                    if (burst_reg == 0) begin
                        // last data word, return to idle
                        m_axil_rready_next = 1'b0;
                        s_axi_rlast_next = 1'b1;
                        s_axi_arready_next = !m_axil_arvalid;
                        state_next = STATE_IDLE;
                    end else begin
                        // start new AXI lite read
                        m_axil_araddr_next = addr_next;
                        m_axil_arvalid_next = 1'b1;
                        m_axil_rready_next = 1'b0;
                        state_next = STATE_DATA;
                    end
                end else begin
                    state_next = STATE_DATA;
                end
            end
            STATE_DATA_READ: begin
                m_axil_rready_next = !s_axi_rvalid && !m_axil_arvalid;

                if (m_axil_rready && m_axil_rvalid) begin
                    s_axi_rid_next = id_reg;
                    data_next = m_axil_rdata;
                    resp_next = m_axil_rresp;
                    s_axi_rdata_next = m_axil_rdata >> (addr_reg[AXIL_ADDR_BIT_OFFSET-1:AXI_ADDR_BIT_OFFSET] * AXI_DATA_WIDTH);
                    s_axi_rresp_next = m_axil_rresp;
                    s_axi_rlast_next = 1'b0;
                    s_axi_rvalid_next = 1'b1;
                    burst_next = burst_reg - 1;
                    addr_next = addr_reg + (1 << burst_size_reg);
                    if (burst_reg == 0) begin
                        m_axil_rready_next = 1'b0;
                        s_axi_arready_next = !m_axil_arvalid;
                        s_axi_rlast_next = 1'b1;
                        state_next = STATE_IDLE;
                    end else if (addr_next[master_burst_size_reg] != addr_reg[master_burst_size_reg]) begin
                        // start new AXI lite read
                        m_axil_araddr_next = addr_next;
                        m_axil_arvalid_next = 1'b1;
                        m_axil_rready_next = 1'b0;
                        state_next = STATE_DATA_READ;
                    end else begin
                        m_axil_rready_next = 1'b0;
                        state_next = STATE_DATA_SPLIT;
                    end
                end else begin
                    state_next = STATE_DATA_READ;
                end
            end
            STATE_DATA_SPLIT: begin
                m_axil_rready_next = 1'b0;

                if (s_axi_rready || !s_axi_rvalid) begin
                    s_axi_rid_next = id_reg;
                    s_axi_rdata_next = data_reg >> (addr_reg[AXIL_ADDR_BIT_OFFSET-1:AXI_ADDR_BIT_OFFSET] * AXI_DATA_WIDTH);
                    s_axi_rresp_next = resp_reg;
                    s_axi_rlast_next = 1'b0;
                    s_axi_rvalid_next = 1'b1;
                    burst_next = burst_reg - 1;
                    addr_next = addr_reg + (1 << burst_size_reg);
                    if (burst_reg == 0) begin
                        s_axi_arready_next = !m_axil_arvalid;
                        s_axi_rlast_next = 1'b1;
                        state_next = STATE_IDLE;
                    end else if (addr_next[master_burst_size_reg] != addr_reg[master_burst_size_reg]) begin
                        // start new AXI lite read
                        m_axil_araddr_next = addr_next;
                        m_axil_arvalid_next = 1'b1;
                        m_axil_rready_next = 1'b0;
                        state_next = STATE_DATA_READ;
                    end else begin
                        state_next = STATE_DATA_SPLIT;
                    end
                end else begin
                    state_next = STATE_DATA_SPLIT;
                end
            end
        endcase
    end else begin
        // master output is narrower; merge reads and possibly split burst
        case (state_reg)
            STATE_IDLE: begin
                // idle state; wait for new burst
                s_axi_arready_next = !m_axil_arvalid;

                resp_next = 2'd0;

                if (s_axi_arready && s_axi_arvalid) begin
                    s_axi_arready_next = 1'b0;
                    id_next = s_axi_arid;
                    m_axil_araddr_next = s_axi_araddr;
                    addr_next = s_axi_araddr;
                    burst_next = s_axi_arlen;
                    burst_size_next = s_axi_arsize;
                    if (s_axi_arsize > AXIL_BURST_SIZE) begin
                        // need to adjust burst size
                        if (s_axi_arlen >> (8+AXIL_BURST_SIZE-s_axi_arsize) != 0) begin
                            // limit burst length to max
                            master_burst_next = (8'd255 << (s_axi_arsize-AXIL_BURST_SIZE)) | ((~s_axi_araddr & (8'hff >> (8-s_axi_arsize))) >> AXIL_BURST_SIZE);
                        end else begin
                            master_burst_next = (s_axi_arlen << (s_axi_arsize-AXIL_BURST_SIZE)) | ((~s_axi_araddr & (8'hff >> (8-s_axi_arsize))) >> AXIL_BURST_SIZE);
                        end
                        master_burst_size_next = AXIL_BURST_SIZE;
                    end else begin
                        // pass through narrow (enough) burst
                        master_burst_next = s_axi_arlen;
                        master_burst_size_next = s_axi_arsize;
                    end
                    m_axil_arprot_next = s_axi_arprot;
                    m_axil_arvalid_next = 1'b1;
                    m_axil_rready_next = 1'b0;
                    state_next = STATE_DATA;
                end else begin
                    state_next = STATE_IDLE;
                end
            end
            STATE_DATA: begin
                m_axil_rready_next = !s_axi_rvalid && !m_axil_arvalid;

                if (m_axil_rready && m_axil_rvalid) begin
                    data_next[addr_reg[AXI_ADDR_BIT_OFFSET-1:AXIL_ADDR_BIT_OFFSET]*SEGMENT_DATA_WIDTH +: SEGMENT_DATA_WIDTH] = m_axil_rdata;
                    if (m_axil_rresp) begin
                        resp_next = m_axil_rresp;
                    end
                    s_axi_rid_next = id_reg;
                    s_axi_rdata_next = data_next;
                    s_axi_rresp_next = resp_next;
                    s_axi_rlast_next = 1'b0;
                    s_axi_rvalid_next = 1'b0;
                    master_burst_next = master_burst_reg - 1;
                    addr_next = (addr_reg + (1 << master_burst_size_reg)) & ({ADDR_WIDTH{1'b1}} << master_burst_size_reg);
                    m_axil_araddr_next = addr_next;
                    if (addr_next[burst_size_reg] != addr_reg[burst_size_reg]) begin
                        data_next = {DATA_WIDTH{1'b0}};
                        burst_next = burst_reg - 1;
                        s_axi_rvalid_next = 1'b1;
                    end
                    if (master_burst_reg == 0) begin
                        if (burst_next >> (8+AXIL_BURST_SIZE-burst_size_reg) != 0) begin
                            // limit burst length to max
                            master_burst_next = 8'd255;
                        end else begin
                            master_burst_next = (burst_next << (burst_size_reg-AXIL_BURST_SIZE)) | (8'hff >> (8-burst_size_reg) >> AXIL_BURST_SIZE);
                        end

                        if (burst_reg == 0) begin
                            m_axil_rready_next = 1'b0;
                            s_axi_rlast_next = 1'b1;
                            s_axi_rvalid_next = 1'b1;
                            s_axi_arready_next = !m_axil_arvalid;
                            state_next = STATE_IDLE;
                        end else begin
                            m_axil_arvalid_next = 1'b1;
                            m_axil_rready_next = 1'b0;
                            state_next = STATE_DATA;
                        end
                    end else begin
                        m_axil_arvalid_next = 1'b1;
                        m_axil_rready_next = 1'b0;
                        state_next = STATE_DATA;
                    end
                end else begin
                    state_next = STATE_DATA;
                end
            end
        endcase
    end
end

always @(posedge clk) begin
    state_reg <= state_next;

    id_reg <= id_next;
    addr_reg <= addr_next;
    data_reg <= data_next;
    resp_reg <= resp_next;
    burst_reg <= burst_next;
    burst_size_reg <= burst_size_next;
    master_burst_reg <= master_burst_next;
    master_burst_size_reg <= master_burst_size_next;

    s_axi_arready_reg <= s_axi_arready_next;
    s_axi_rid_reg <= s_axi_rid_next;
    s_axi_rdata_reg <= s_axi_rdata_next;
    s_axi_rresp_reg <= s_axi_rresp_next;
    s_axi_rlast_reg <= s_axi_rlast_next;
    s_axi_rvalid_reg <= s_axi_rvalid_next;

    m_axil_araddr_reg <= m_axil_araddr_next;
    m_axil_arprot_reg <= m_axil_arprot_next;
    m_axil_arvalid_reg <= m_axil_arvalid_next;
    m_axil_rready_reg <= m_axil_rready_next;

    if (rst) begin
        state_reg <= STATE_IDLE;

        s_axi_arready_reg <= 1'b0;
        s_axi_rvalid_reg <= 1'b0;

        m_axil_arvalid_reg <= 1'b0;
        m_axil_rready_reg <= 1'b0;
    end
end

endmodule

`resetall


// Content from axi_axil_adapter.v
/*

Copyright (c) 2019 Alex Forencich

Permission is hereby granted, free of charge, to any person obtaining a copy
of this software and associated documentation files (the "Software"), to deal
in the Software without restriction, including without limitation the rights
to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
copies of the Software, and to permit persons to whom the Software is
furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in
all copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY
FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
THE SOFTWARE.

*/

// Language: Verilog 2001

/*
 * AXI4 to AXI4-Lite adapter
 */
module axi_axil_adapter #
(
    // Width of address bus in bits
    parameter ADDR_WIDTH = 32,
    // Width of input (slave) AXI interface data bus in bits
    parameter AXI_DATA_WIDTH = 32,
    // Width of input (slave) AXI interface wstrb (width of data bus in words)
    parameter AXI_STRB_WIDTH = (AXI_DATA_WIDTH/8),
    // Width of AXI ID signal
    parameter AXI_ID_WIDTH = 8,
    // Width of output (master) AXI lite interface data bus in bits
    parameter AXIL_DATA_WIDTH = 32,
    // Width of output (master) AXI lite interface wstrb (width of data bus in words)
    parameter AXIL_STRB_WIDTH = (AXIL_DATA_WIDTH/8),
    // When adapting to a wider bus, re-pack full-width burst instead of passing through narrow burst if possible
    parameter CONVERT_BURST = 1,
    // When adapting to a wider bus, re-pack all bursts instead of passing through narrow burst if possible
    parameter CONVERT_NARROW_BURST = 0
)
(
    input  wire                        clk,
    input  wire                        rst,

    /*
     * AXI slave interface
     */
    input  wire [AXI_ID_WIDTH-1:0]     s_axi_awid,
    input  wire [ADDR_WIDTH-1:0]       s_axi_awaddr,
    input  wire [7:0]                  s_axi_awlen,
    input  wire [2:0]                  s_axi_awsize,
    input  wire [1:0]                  s_axi_awburst,
    input  wire                        s_axi_awlock,
    input  wire [3:0]                  s_axi_awcache,
    input  wire [2:0]                  s_axi_awprot,
    input  wire                        s_axi_awvalid,
    output wire                        s_axi_awready,
    input  wire [AXI_DATA_WIDTH-1:0]   s_axi_wdata,
    input  wire [AXI_STRB_WIDTH-1:0]   s_axi_wstrb,
    input  wire                        s_axi_wlast,
    input  wire                        s_axi_wvalid,
    output wire                        s_axi_wready,
    output wire [AXI_ID_WIDTH-1:0]     s_axi_bid,
    output wire [1:0]                  s_axi_bresp,
    output wire                        s_axi_bvalid,
    input  wire                        s_axi_bready,
    input  wire [AXI_ID_WIDTH-1:0]     s_axi_arid,
    input  wire [ADDR_WIDTH-1:0]       s_axi_araddr,
    input  wire [7:0]                  s_axi_arlen,
    input  wire [2:0]                  s_axi_arsize,
    input  wire [1:0]                  s_axi_arburst,
    input  wire                        s_axi_arlock,
    input  wire [3:0]                  s_axi_arcache,
    input  wire [2:0]                  s_axi_arprot,
    input  wire                        s_axi_arvalid,
    output wire                        s_axi_arready,
    output wire [AXI_ID_WIDTH-1:0]     s_axi_rid,
    output wire [AXI_DATA_WIDTH-1:0]   s_axi_rdata,
    output wire [1:0]                  s_axi_rresp,
    output wire                        s_axi_rlast,
    output wire                        s_axi_rvalid,
    input  wire                        s_axi_rready,

    /*
     * AXI lite master interface
     */
    output wire [ADDR_WIDTH-1:0]       m_axil_awaddr,
    output wire [2:0]                  m_axil_awprot,
    output wire                        m_axil_awvalid,
    input  wire                        m_axil_awready,
    output wire [AXIL_DATA_WIDTH-1:0]  m_axil_wdata,
    output wire [AXIL_STRB_WIDTH-1:0]  m_axil_wstrb,
    output wire                        m_axil_wvalid,
    input  wire                        m_axil_wready,
    input  wire [1:0]                  m_axil_bresp,
    input  wire                        m_axil_bvalid,
    output wire                        m_axil_bready,
    output wire [ADDR_WIDTH-1:0]       m_axil_araddr,
    output wire [2:0]                  m_axil_arprot,
    output wire                        m_axil_arvalid,
    input  wire                        m_axil_arready,
    input  wire [AXIL_DATA_WIDTH-1:0]  m_axil_rdata,
    input  wire [1:0]                  m_axil_rresp,
    input  wire                        m_axil_rvalid,
    output wire                        m_axil_rready
);


axi_axil_adapter_wr #(
    .ADDR_WIDTH(ADDR_WIDTH),
    .AXI_DATA_WIDTH(AXI_DATA_WIDTH),
    .AXI_STRB_WIDTH(AXI_STRB_WIDTH),
    .AXI_ID_WIDTH(AXI_ID_WIDTH),
    .AXIL_DATA_WIDTH(AXIL_DATA_WIDTH),
    .AXIL_STRB_WIDTH(AXIL_STRB_WIDTH),
    .CONVERT_BURST(CONVERT_BURST),
    .CONVERT_NARROW_BURST(CONVERT_NARROW_BURST)
)
axi_axil_adapter_wr_inst (
    .clk(clk),
    .rst(rst),

    /*
     * AXI slave interface
     */
    .s_axi_awid(s_axi_awid),
    .s_axi_awaddr(s_axi_awaddr),
    .s_axi_awlen(s_axi_awlen),
    .s_axi_awsize(s_axi_awsize),
    .s_axi_awburst(s_axi_awburst),
    .s_axi_awlock(s_axi_awlock),
    .s_axi_awcache(s_axi_awcache),
    .s_axi_awprot(s_axi_awprot),
    .s_axi_awvalid(s_axi_awvalid),
    .s_axi_awready(s_axi_awready),
    .s_axi_wdata(s_axi_wdata),
    .s_axi_wstrb(s_axi_wstrb),
    .s_axi_wlast(s_axi_wlast),
    .s_axi_wvalid(s_axi_wvalid),
    .s_axi_wready(s_axi_wready),
    .s_axi_bid(s_axi_bid),
    .s_axi_bresp(s_axi_bresp),
    .s_axi_bvalid(s_axi_bvalid),
    .s_axi_bready(s_axi_bready),

    /*
     * AXI lite master interface
     */
    .m_axil_awaddr(m_axil_awaddr),
    .m_axil_awprot(m_axil_awprot),
    .m_axil_awvalid(m_axil_awvalid),
    .m_axil_awready(m_axil_awready),
    .m_axil_wdata(m_axil_wdata),
    .m_axil_wstrb(m_axil_wstrb),
    .m_axil_wvalid(m_axil_wvalid),
    .m_axil_wready(m_axil_wready),
    .m_axil_bresp(m_axil_bresp),
    .m_axil_bvalid(m_axil_bvalid),
    .m_axil_bready(m_axil_bready)
);

axi_axil_adapter_rd #(
    .ADDR_WIDTH(ADDR_WIDTH),
    .AXI_DATA_WIDTH(AXI_DATA_WIDTH),
    .AXI_STRB_WIDTH(AXI_STRB_WIDTH),
    .AXI_ID_WIDTH(AXI_ID_WIDTH),
    .AXIL_DATA_WIDTH(AXIL_DATA_WIDTH),
    .AXIL_STRB_WIDTH(AXIL_STRB_WIDTH),
    .CONVERT_BURST(CONVERT_BURST),
    .CONVERT_NARROW_BURST(CONVERT_NARROW_BURST)
)
axi_axil_adapter_rd_inst (
    .clk(clk),
    .rst(rst),

    /*
     * AXI slave interface
     */
    .s_axi_arid(s_axi_arid),
    .s_axi_araddr(s_axi_araddr),
    .s_axi_arlen(s_axi_arlen),
    .s_axi_arsize(s_axi_arsize),
    .s_axi_arburst(s_axi_arburst),
    .s_axi_arlock(s_axi_arlock),
    .s_axi_arcache(s_axi_arcache),
    .s_axi_arprot(s_axi_arprot),
    .s_axi_arvalid(s_axi_arvalid),
    .s_axi_arready(s_axi_arready),
    .s_axi_rid(s_axi_rid),
    .s_axi_rdata(s_axi_rdata),
    .s_axi_rresp(s_axi_rresp),
    .s_axi_rlast(s_axi_rlast),
    .s_axi_rvalid(s_axi_rvalid),
    .s_axi_rready(s_axi_rready),

    /*
     * AXI lite master interface
     */
    .m_axil_araddr(m_axil_araddr),
    .m_axil_arprot(m_axil_arprot),
    .m_axil_arvalid(m_axil_arvalid),
    .m_axil_arready(m_axil_arready),
    .m_axil_rdata(m_axil_rdata),
    .m_axil_rresp(m_axil_rresp),
    .m_axil_rvalid(m_axil_rvalid),
    .m_axil_rready(m_axil_rready)
);

endmodule

`resetall


// Content from axil_interconnect.v
/*

Copyright (c) 2018 Alex Forencich

Permission is hereby granted, free of charge, to any person obtaining a copy
of this software and associated documentation files (the "Software"), to deal
in the Software without restriction, including without limitation the rights
to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
copies of the Software, and to permit persons to whom the Software is
furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in
all copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY
FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
THE SOFTWARE.

*/

// Language: Verilog 2001

/*
 * AXI4 lite interconnect
 */
module axil_interconnect #
(
    // Number of AXI inputs (slave interfaces)
    parameter S_COUNT = 4,
    // Number of AXI outputs (master interfaces)
    parameter M_COUNT = 4,
    // Width of data bus in bits
    parameter DATA_WIDTH = 32,
    // Width of address bus in bits
    parameter ADDR_WIDTH = 32,
    // Width of wstrb (width of data bus in words)
    parameter STRB_WIDTH = (DATA_WIDTH/8),
    // Number of regions per master interface
    parameter M_REGIONS = 1,
    // Master interface base addresses
    // M_COUNT concatenated fields of M_REGIONS concatenated fields of ADDR_WIDTH bits
    // set to zero for default addressing based on M_ADDR_WIDTH
    parameter M_BASE_ADDR = 0,
    // Master interface address widths
    // M_COUNT concatenated fields of M_REGIONS concatenated fields of 32 bits
    parameter M_ADDR_WIDTH = {M_COUNT{{M_REGIONS{32'd24}}}},
    // Read connections between interfaces
    // M_COUNT concatenated fields of S_COUNT bits
    parameter M_CONNECT_READ = {M_COUNT{{S_COUNT{1'b1}}}},
    // Write connections between interfaces
    // M_COUNT concatenated fields of S_COUNT bits
    parameter M_CONNECT_WRITE = {M_COUNT{{S_COUNT{1'b1}}}},
    // Secure master (fail operations based on awprot/arprot)
    // M_COUNT bits
    parameter M_SECURE = {M_COUNT{1'b0}}
)
(
    input  wire                           clk,
    input  wire                           rst,

    /*
     * AXI lite slave interfaces
     */
    input  wire [S_COUNT*ADDR_WIDTH-1:0]  s_axil_awaddr,
    input  wire [S_COUNT*3-1:0]           s_axil_awprot,
    input  wire [S_COUNT-1:0]             s_axil_awvalid,
    output wire [S_COUNT-1:0]             s_axil_awready,
    input  wire [S_COUNT*DATA_WIDTH-1:0]  s_axil_wdata,
    input  wire [S_COUNT*STRB_WIDTH-1:0]  s_axil_wstrb,
    input  wire [S_COUNT-1:0]             s_axil_wvalid,
    output wire [S_COUNT-1:0]             s_axil_wready,
    output wire [S_COUNT*2-1:0]           s_axil_bresp,
    output wire [S_COUNT-1:0]             s_axil_bvalid,
    input  wire [S_COUNT-1:0]             s_axil_bready,
    input  wire [S_COUNT*ADDR_WIDTH-1:0]  s_axil_araddr,
    input  wire [S_COUNT*3-1:0]           s_axil_arprot,
    input  wire [S_COUNT-1:0]             s_axil_arvalid,
    output wire [S_COUNT-1:0]             s_axil_arready,
    output wire [S_COUNT*DATA_WIDTH-1:0]  s_axil_rdata,
    output wire [S_COUNT*2-1:0]           s_axil_rresp,
    output wire [S_COUNT-1:0]             s_axil_rvalid,
    input  wire [S_COUNT-1:0]             s_axil_rready,

    /*
     * AXI lite master interfaces
     */
    output wire [M_COUNT*ADDR_WIDTH-1:0]  m_axil_awaddr,
    output wire [M_COUNT*3-1:0]           m_axil_awprot,
    output wire [M_COUNT-1:0]             m_axil_awvalid,
    input  wire [M_COUNT-1:0]             m_axil_awready,
    output wire [M_COUNT*DATA_WIDTH-1:0]  m_axil_wdata,
    output wire [M_COUNT*STRB_WIDTH-1:0]  m_axil_wstrb,
    output wire [M_COUNT-1:0]             m_axil_wvalid,
    input  wire [M_COUNT-1:0]             m_axil_wready,
    input  wire [M_COUNT*2-1:0]           m_axil_bresp,
    input  wire [M_COUNT-1:0]             m_axil_bvalid,
    output wire [M_COUNT-1:0]             m_axil_bready,
    output wire [M_COUNT*ADDR_WIDTH-1:0]  m_axil_araddr,
    output wire [M_COUNT*3-1:0]           m_axil_arprot,
    output wire [M_COUNT-1:0]             m_axil_arvalid,
    input  wire [M_COUNT-1:0]             m_axil_arready,
    input  wire [M_COUNT*DATA_WIDTH-1:0]  m_axil_rdata,
    input  wire [M_COUNT*2-1:0]           m_axil_rresp,
    input  wire [M_COUNT-1:0]             m_axil_rvalid,
    output wire [M_COUNT-1:0]             m_axil_rready
);

parameter CL_S_COUNT = $clog2(S_COUNT);
parameter CL_M_COUNT = $clog2(M_COUNT);

// default address computation
function [M_COUNT*M_REGIONS*ADDR_WIDTH-1:0] calcBaseAddrs(input [31:0] dummy);
    integer i;
    reg [ADDR_WIDTH-1:0] base;
    reg [ADDR_WIDTH-1:0] width;
    reg [ADDR_WIDTH-1:0] size;
    reg [ADDR_WIDTH-1:0] mask;
    begin
        calcBaseAddrs = {M_COUNT*M_REGIONS*ADDR_WIDTH{1'b0}};
        base = 0;
        for (i = 0; i < M_COUNT*M_REGIONS; i = i + 1) begin
            width = M_ADDR_WIDTH[i*32 +: 32];
            mask = {ADDR_WIDTH{1'b1}} >> (ADDR_WIDTH - width);
            size = mask + 1;
            if (width > 0) begin
                if ((base & mask) != 0) begin
                   base = base + size - (base & mask); // align
                end
                calcBaseAddrs[i * ADDR_WIDTH +: ADDR_WIDTH] = base;
                base = base + size; // increment
            end
        end
    end
endfunction

parameter M_BASE_ADDR_INT = M_BASE_ADDR ? M_BASE_ADDR : calcBaseAddrs(0);

integer i, j;

// check configuration
initial begin
    $display("Addressing configuration for axil_interconnect instance %m");
    for (i = 0; i < M_COUNT*M_REGIONS; i = i + 1) begin
        if (M_ADDR_WIDTH[i*32 +: 32]) begin
            $display("%2d (%2d): %x / %02d -- %x-%x",
                i/M_REGIONS, i%M_REGIONS,
                M_BASE_ADDR_INT[i*ADDR_WIDTH +: ADDR_WIDTH],
                M_ADDR_WIDTH[i*32 +: 32],
                M_BASE_ADDR_INT[i*ADDR_WIDTH +: ADDR_WIDTH] & ({ADDR_WIDTH{1'b1}} << M_ADDR_WIDTH[i*32 +: 32]),
                M_BASE_ADDR_INT[i*ADDR_WIDTH +: ADDR_WIDTH] | ({ADDR_WIDTH{1'b1}} >> (ADDR_WIDTH - M_ADDR_WIDTH[i*32 +: 32]))
            );
        end
    end

    for (i = 0; i < M_COUNT*M_REGIONS; i = i + 1) begin
        if ((M_BASE_ADDR_INT[i*ADDR_WIDTH +: ADDR_WIDTH] & (2**M_ADDR_WIDTH[i*32 +: 32]-1)) != 0) begin
            $display("Region not aligned:");
            $display("%2d (%2d): %x / %2d -- %x-%x",
                i/M_REGIONS, i%M_REGIONS,
                M_BASE_ADDR_INT[i*ADDR_WIDTH +: ADDR_WIDTH],
                M_ADDR_WIDTH[i*32 +: 32],
                M_BASE_ADDR_INT[i*ADDR_WIDTH +: ADDR_WIDTH] & ({ADDR_WIDTH{1'b1}} << M_ADDR_WIDTH[i*32 +: 32]),
                M_BASE_ADDR_INT[i*ADDR_WIDTH +: ADDR_WIDTH] | ({ADDR_WIDTH{1'b1}} >> (ADDR_WIDTH - M_ADDR_WIDTH[i*32 +: 32]))
            );
        end
    end

    for (i = 0; i < M_COUNT*M_REGIONS; i = i + 1) begin
        for (j = i+1; j < M_COUNT*M_REGIONS; j = j + 1) begin
            if (M_ADDR_WIDTH[i*32 +: 32] && M_ADDR_WIDTH[j*32 +: 32]) begin
                if (((M_BASE_ADDR_INT[i*ADDR_WIDTH +: ADDR_WIDTH] & ({ADDR_WIDTH{1'b1}} << M_ADDR_WIDTH[i*32 +: 32])) <= (M_BASE_ADDR_INT[j*ADDR_WIDTH +: ADDR_WIDTH] | ({ADDR_WIDTH{1'b1}} >> (ADDR_WIDTH - M_ADDR_WIDTH[j*32 +: 32]))))
                        && ((M_BASE_ADDR_INT[j*ADDR_WIDTH +: ADDR_WIDTH] & ({ADDR_WIDTH{1'b1}} << M_ADDR_WIDTH[j*32 +: 32])) <= (M_BASE_ADDR_INT[i*ADDR_WIDTH +: ADDR_WIDTH] | ({ADDR_WIDTH{1'b1}} >> (ADDR_WIDTH - M_ADDR_WIDTH[i*32 +: 32]))))) begin
                    $display("Overlapping regions:");
                    $display("%2d (%2d): %x / %2d -- %x-%x",
                        i/M_REGIONS, i%M_REGIONS,
                        M_BASE_ADDR_INT[i*ADDR_WIDTH +: ADDR_WIDTH],
                        M_ADDR_WIDTH[i*32 +: 32],
                        M_BASE_ADDR_INT[i*ADDR_WIDTH +: ADDR_WIDTH] & ({ADDR_WIDTH{1'b1}} << M_ADDR_WIDTH[i*32 +: 32]),
                        M_BASE_ADDR_INT[i*ADDR_WIDTH +: ADDR_WIDTH] | ({ADDR_WIDTH{1'b1}} >> (ADDR_WIDTH - M_ADDR_WIDTH[i*32 +: 32]))
                    );
                    $display("%2d (%2d): %x / %2d -- %x-%x",
                        j/M_REGIONS, j%M_REGIONS,
                        M_BASE_ADDR_INT[j*ADDR_WIDTH +: ADDR_WIDTH],
                        M_ADDR_WIDTH[j*32 +: 32],
                        M_BASE_ADDR_INT[j*ADDR_WIDTH +: ADDR_WIDTH] & ({ADDR_WIDTH{1'b1}} << M_ADDR_WIDTH[j*32 +: 32]),
                        M_BASE_ADDR_INT[j*ADDR_WIDTH +: ADDR_WIDTH] | ({ADDR_WIDTH{1'b1}} >> (ADDR_WIDTH - M_ADDR_WIDTH[j*32 +: 32]))
                    );
                end
            end
        end
    end
end

localparam [2:0]
    STATE_IDLE = 3'd0,
    STATE_DECODE = 3'd1,
    STATE_WRITE = 3'd2,
    STATE_WRITE_RESP = 3'd3,
    STATE_WRITE_DROP = 3'd4,
    STATE_READ = 3'd5,
    STATE_WAIT_IDLE = 3'd6;

reg [2:0] state_reg = STATE_IDLE, state_next;

reg match;

reg [CL_M_COUNT-1:0] m_select_reg = 2'd0, m_select_next;
reg [ADDR_WIDTH-1:0] axil_addr_reg = {ADDR_WIDTH{1'b0}}, axil_addr_next;
reg axil_addr_valid_reg = 1'b0, axil_addr_valid_next;
reg [2:0] axil_prot_reg = 3'b000, axil_prot_next;
reg [DATA_WIDTH-1:0] axil_data_reg = {DATA_WIDTH{1'b0}}, axil_data_next;
reg [STRB_WIDTH-1:0] axil_wstrb_reg = {STRB_WIDTH{1'b0}}, axil_wstrb_next;
reg [1:0] axil_resp_reg = 2'b00, axil_resp_next;

reg [S_COUNT-1:0] s_axil_awready_reg = 0, s_axil_awready_next;
reg [S_COUNT-1:0] s_axil_wready_reg = 0, s_axil_wready_next;
reg [S_COUNT-1:0] s_axil_bvalid_reg = 0, s_axil_bvalid_next;
reg [S_COUNT-1:0] s_axil_arready_reg = 0, s_axil_arready_next;
reg [S_COUNT-1:0] s_axil_rvalid_reg = 0, s_axil_rvalid_next;

reg [M_COUNT-1:0] m_axil_awvalid_reg = 0, m_axil_awvalid_next;
reg [M_COUNT-1:0] m_axil_wvalid_reg = 0, m_axil_wvalid_next;
reg [M_COUNT-1:0] m_axil_bready_reg = 0, m_axil_bready_next;
reg [M_COUNT-1:0] m_axil_arvalid_reg = 0, m_axil_arvalid_next;
reg [M_COUNT-1:0] m_axil_rready_reg = 0, m_axil_rready_next;

assign s_axil_awready = s_axil_awready_reg;
assign s_axil_wready = s_axil_wready_reg;
assign s_axil_bresp = {S_COUNT{axil_resp_reg}};
assign s_axil_bvalid = s_axil_bvalid_reg;
assign s_axil_arready = s_axil_arready_reg;
assign s_axil_rdata = {S_COUNT{axil_data_reg}};
assign s_axil_rresp = {S_COUNT{axil_resp_reg}};
assign s_axil_rvalid = s_axil_rvalid_reg;

assign m_axil_awaddr = {M_COUNT{axil_addr_reg}};
assign m_axil_awprot = {M_COUNT{axil_prot_reg}};
assign m_axil_awvalid = m_axil_awvalid_reg;
assign m_axil_wdata = {M_COUNT{axil_data_reg}};
assign m_axil_wstrb = {M_COUNT{axil_wstrb_reg}};
assign m_axil_wvalid = m_axil_wvalid_reg;
assign m_axil_bready = m_axil_bready_reg;
assign m_axil_araddr = {M_COUNT{axil_addr_reg}};
assign m_axil_arprot = {M_COUNT{axil_prot_reg}};
assign m_axil_arvalid = m_axil_arvalid_reg;
assign m_axil_rready = m_axil_rready_reg;

// slave side mux
wire [(CL_S_COUNT > 0 ? CL_S_COUNT-1 : 0):0] s_select;

wire [ADDR_WIDTH-1:0] current_s_axil_awaddr  = s_axil_awaddr[s_select*ADDR_WIDTH +: ADDR_WIDTH];
wire [2:0]            current_s_axil_awprot  = s_axil_awprot[s_select*3 +: 3];
wire                  current_s_axil_awvalid = s_axil_awvalid[s_select];
wire                  current_s_axil_awready = s_axil_awready[s_select];
wire [DATA_WIDTH-1:0] current_s_axil_wdata   = s_axil_wdata[s_select*DATA_WIDTH +: DATA_WIDTH];
wire [STRB_WIDTH-1:0] current_s_axil_wstrb   = s_axil_wstrb[s_select*STRB_WIDTH +: STRB_WIDTH];
wire                  current_s_axil_wvalid  = s_axil_wvalid[s_select];
wire                  current_s_axil_wready  = s_axil_wready[s_select];
wire [1:0]            current_s_axil_bresp   = s_axil_bresp[s_select*2 +: 2];
wire                  current_s_axil_bvalid  = s_axil_bvalid[s_select];
wire                  current_s_axil_bready  = s_axil_bready[s_select];
wire [ADDR_WIDTH-1:0] current_s_axil_araddr  = s_axil_araddr[s_select*ADDR_WIDTH +: ADDR_WIDTH];
wire [2:0]            current_s_axil_arprot  = s_axil_arprot[s_select*3 +: 3];
wire                  current_s_axil_arvalid = s_axil_arvalid[s_select];
wire                  current_s_axil_arready = s_axil_arready[s_select];
wire [DATA_WIDTH-1:0] current_s_axil_rdata   = s_axil_rdata[s_select*DATA_WIDTH +: DATA_WIDTH];
wire [1:0]            current_s_axil_rresp   = s_axil_rresp[s_select*2 +: 2];
wire                  current_s_axil_rvalid  = s_axil_rvalid[s_select];
wire                  current_s_axil_rready  = s_axil_rready[s_select];

// master side mux
wire [ADDR_WIDTH-1:0] current_m_axil_awaddr  = m_axil_awaddr[m_select_reg*ADDR_WIDTH +: ADDR_WIDTH];
wire [2:0]            current_m_axil_awprot  = m_axil_awprot[m_select_reg*3 +: 3];
wire                  current_m_axil_awvalid = m_axil_awvalid[m_select_reg];
wire                  current_m_axil_awready = m_axil_awready[m_select_reg];
wire [DATA_WIDTH-1:0] current_m_axil_wdata   = m_axil_wdata[m_select_reg*DATA_WIDTH +: DATA_WIDTH];
wire [STRB_WIDTH-1:0] current_m_axil_wstrb   = m_axil_wstrb[m_select_reg*STRB_WIDTH +: STRB_WIDTH];
wire                  current_m_axil_wvalid  = m_axil_wvalid[m_select_reg];
wire                  current_m_axil_wready  = m_axil_wready[m_select_reg];
wire [1:0]            current_m_axil_bresp   = m_axil_bresp[m_select_reg*2 +: 2];
wire                  current_m_axil_bvalid  = m_axil_bvalid[m_select_reg];
wire                  current_m_axil_bready  = m_axil_bready[m_select_reg];
wire [ADDR_WIDTH-1:0] current_m_axil_araddr  = m_axil_araddr[m_select_reg*ADDR_WIDTH +: ADDR_WIDTH];
wire [2:0]            current_m_axil_arprot  = m_axil_arprot[m_select_reg*3 +: 3];
wire                  current_m_axil_arvalid = m_axil_arvalid[m_select_reg];
wire                  current_m_axil_arready = m_axil_arready[m_select_reg];
wire [DATA_WIDTH-1:0] current_m_axil_rdata   = m_axil_rdata[m_select_reg*DATA_WIDTH +: DATA_WIDTH];
wire [1:0]            current_m_axil_rresp   = m_axil_rresp[m_select_reg*2 +: 2];
wire                  current_m_axil_rvalid  = m_axil_rvalid[m_select_reg];
wire                  current_m_axil_rready  = m_axil_rready[m_select_reg];

// arbiter instance
wire [S_COUNT*2-1:0] request;
wire [S_COUNT*2-1:0] acknowledge;
wire [S_COUNT*2-1:0] grant;
wire grant_valid;
wire [CL_S_COUNT:0] grant_encoded;

wire read = grant_encoded[0];
assign s_select = grant_encoded >> 1;

arbiter #(
    .PORTS(S_COUNT*2),
    .ARB_TYPE_ROUND_ROBIN(1),
    .ARB_BLOCK(1),
    .ARB_BLOCK_ACK(1),
    .ARB_LSB_HIGH_PRIORITY(1)
)
arb_inst (
    .clk(clk),
    .rst(rst),
    .request(request),
    .acknowledge(acknowledge),
    .grant(grant),
    .grant_valid(grant_valid),
    .grant_encoded(grant_encoded)
);

genvar n;

// request generation
generate
for (n = 0; n < S_COUNT; n = n + 1) begin
    assign request[2*n]   = s_axil_awvalid[n];
    assign request[2*n+1] = s_axil_arvalid[n];
end
endgenerate

// acknowledge generation
generate
for (n = 0; n < S_COUNT; n = n + 1) begin
    assign acknowledge[2*n]   = grant[2*n]   && s_axil_bvalid[n] && s_axil_bready[n];
    assign acknowledge[2*n+1] = grant[2*n+1] && s_axil_rvalid[n] && s_axil_rready[n];
end
endgenerate

always @* begin
    state_next = STATE_IDLE;

    match = 1'b0;

    m_select_next = m_select_reg;
    axil_addr_next = axil_addr_reg;
    axil_addr_valid_next = axil_addr_valid_reg;
    axil_prot_next = axil_prot_reg;
    axil_data_next = axil_data_reg;
    axil_wstrb_next = axil_wstrb_reg;
    axil_resp_next = axil_resp_reg;

    s_axil_awready_next = 0;
    s_axil_wready_next = 0;
    s_axil_bvalid_next = s_axil_bvalid_reg & ~s_axil_bready;
    s_axil_arready_next = 0;
    s_axil_rvalid_next = s_axil_rvalid_reg & ~s_axil_rready;

    m_axil_awvalid_next = m_axil_awvalid_reg & ~m_axil_awready;
    m_axil_wvalid_next = m_axil_wvalid_reg & ~m_axil_wready;
    m_axil_bready_next = 0;
    m_axil_arvalid_next = m_axil_arvalid_reg & ~m_axil_arready;
    m_axil_rready_next = 0;

    case (state_reg)
        STATE_IDLE: begin
            // idle state; wait for arbitration

            if (grant_valid) begin

                axil_addr_valid_next = 1'b1;

                if (read) begin
                    // reading
                    axil_addr_next = current_s_axil_araddr;
                    axil_prot_next = current_s_axil_arprot;
                    s_axil_arready_next[s_select] = 1'b1;
                end else  begin
                    // writing
                    axil_addr_next = current_s_axil_awaddr;
                    axil_prot_next = current_s_axil_awprot;
                    s_axil_awready_next[s_select] = 1'b1;
                end

                state_next = STATE_DECODE;
            end else begin
                state_next = STATE_IDLE;
            end
        end
        STATE_DECODE: begin
            // decode state; determine master interface

            match = 1'b0;
            for (i = 0; i < M_COUNT; i = i + 1) begin
                for (j = 0; j < M_REGIONS; j = j + 1) begin
                    if (M_ADDR_WIDTH[(i*M_REGIONS+j)*32 +: 32] && (!M_SECURE[i] || !axil_prot_reg[1]) && ((read ? M_CONNECT_READ : M_CONNECT_WRITE) & (1 << (s_select+i*S_COUNT))) && (axil_addr_reg >> M_ADDR_WIDTH[(i*M_REGIONS+j)*32 +: 32]) == (M_BASE_ADDR_INT[(i*M_REGIONS+j)*ADDR_WIDTH +: ADDR_WIDTH] >> M_ADDR_WIDTH[(i*M_REGIONS+j)*32 +: 32])) begin
                        m_select_next = i;
                        match = 1'b1;
                    end
                end
            end

            if (match) begin
                if (read) begin
                    // reading
                    m_axil_rready_next[m_select_next] = 1'b1;
                    state_next = STATE_READ;
                end else begin
                    // writing
                    s_axil_wready_next[s_select] = 1'b1;
                    state_next = STATE_WRITE;
                end
            end else begin
                // no match; return decode error
                axil_data_next = {DATA_WIDTH{1'b0}};
                axil_resp_next = 2'b11;
                if (read) begin
                    // reading
                    s_axil_rvalid_next[s_select] = 1'b1;
                    state_next = STATE_WAIT_IDLE;
                end else begin
                    // writing
                    s_axil_wready_next[s_select] = 1'b1;
                    state_next = STATE_WRITE_DROP;
                end
            end
        end
        STATE_WRITE: begin
            // write state; store and forward write data
            s_axil_wready_next[s_select] = 1'b1;

            if (axil_addr_valid_reg) begin
                m_axil_awvalid_next[m_select_reg] = 1'b1;
            end
            axil_addr_valid_next = 1'b0;

            if (current_s_axil_wready && current_s_axil_wvalid) begin
                s_axil_wready_next[s_select] = 1'b0;
                axil_data_next = current_s_axil_wdata;
                axil_wstrb_next = current_s_axil_wstrb;
                m_axil_wvalid_next[m_select_reg] = 1'b1;
                m_axil_bready_next[m_select_reg] = 1'b1;
                state_next = STATE_WRITE_RESP;
            end else begin
                state_next = STATE_WRITE;
            end
        end
        STATE_WRITE_RESP: begin
            // write response state; store and forward write response
            m_axil_bready_next[m_select_reg] = 1'b1;

            if (current_m_axil_bready && current_m_axil_bvalid) begin
                m_axil_bready_next[m_select_reg] = 1'b0;
                axil_resp_next = current_m_axil_bresp;
                s_axil_bvalid_next[s_select] = 1'b1;
                state_next = STATE_WAIT_IDLE;
            end else begin
                state_next = STATE_WRITE_RESP;
            end
        end
        STATE_WRITE_DROP: begin
            // write drop state; drop write data
            s_axil_wready_next[s_select] = 1'b1;

            axil_addr_valid_next = 1'b0;

            if (current_s_axil_wready && current_s_axil_wvalid) begin
                s_axil_wready_next[s_select] = 1'b0;
                s_axil_bvalid_next[s_select] = 1'b1;
                state_next = STATE_WAIT_IDLE;
            end else begin
                state_next = STATE_WRITE_DROP;
            end
        end
        STATE_READ: begin
            // read state; store and forward read response
            m_axil_rready_next[m_select_reg] = 1'b1;

            if (axil_addr_valid_reg) begin
                m_axil_arvalid_next[m_select_reg] = 1'b1;
            end
            axil_addr_valid_next = 1'b0;

            if (current_m_axil_rready && current_m_axil_rvalid) begin
                m_axil_rready_next[m_select_reg] = 1'b0;
                axil_data_next = current_m_axil_rdata;
                axil_resp_next = current_m_axil_rresp;
                s_axil_rvalid_next[s_select] = 1'b1;
                state_next = STATE_WAIT_IDLE;
            end else begin
                state_next = STATE_READ;
            end
        end
        STATE_WAIT_IDLE: begin
            // wait for idle state; wait untl grant valid is deasserted

            if (!grant_valid || acknowledge) begin
                state_next = STATE_IDLE;
            end else begin
                state_next = STATE_WAIT_IDLE;
            end
        end
    endcase
end

always @(posedge clk) begin
    if (rst) begin
        state_reg <= STATE_IDLE;

        s_axil_awready_reg <= 0;
        s_axil_wready_reg <= 0;
        s_axil_bvalid_reg <= 0;
        s_axil_arready_reg <= 0;
        s_axil_rvalid_reg <= 0;

        m_axil_awvalid_reg <= 0;
        m_axil_wvalid_reg <= 0;
        m_axil_bready_reg <= 0;
        m_axil_arvalid_reg <= 0;
        m_axil_rready_reg <= 0;
    end else begin
        state_reg <= state_next;

        s_axil_awready_reg <= s_axil_awready_next;
        s_axil_wready_reg <= s_axil_wready_next;
        s_axil_bvalid_reg <= s_axil_bvalid_next;
        s_axil_arready_reg <= s_axil_arready_next;
        s_axil_rvalid_reg <= s_axil_rvalid_next;

        m_axil_awvalid_reg <= m_axil_awvalid_next;
        m_axil_wvalid_reg <= m_axil_wvalid_next;
        m_axil_bready_reg <= m_axil_bready_next;
        m_axil_arvalid_reg <= m_axil_arvalid_next;
        m_axil_rready_reg <= m_axil_rready_next;
    end

    m_select_reg <= m_select_next;
    axil_addr_reg <= axil_addr_next;
    axil_addr_valid_reg <= axil_addr_valid_next;
    axil_prot_reg <= axil_prot_next;
    axil_data_reg <= axil_data_next;
    axil_wstrb_reg <= axil_wstrb_next;
    axil_resp_reg <= axil_resp_next;
end

endmodule

`resetall


// Content from kmeans.v
// Content from kmeans_top.v
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2022.2 (64-bit)
// Version: 2022.2
// Copyright (C) Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

(* CORE_GENERATION_INFO="kmeans_top_kmeans_top,hls_ip_2022_2,{HLS_INPUT_TYPE=cxx,HLS_INPUT_FLOAT=0,HLS_INPUT_FIXED=0,HLS_INPUT_PART=xcvc1902-vsva2197-2MP-e-S,HLS_INPUT_CLOCK=5.000000,HLS_INPUT_ARCH=others,HLS_SYN_CLOCK=4.950000,HLS_SYN_LAT=-1,HLS_SYN_TPT=none,HLS_SYN_MEM=11,HLS_SYN_DSP=0,HLS_SYN_FF=9239,HLS_SYN_LUT=12196,HLS_VERSION=2022_2}" *)

module kmeans_flat (
        ap_clk,
        ap_rst_n,
        m_axi_mem_AWVALID,
        m_axi_mem_AWREADY,
        m_axi_mem_AWADDR,
        m_axi_mem_AWID,
        m_axi_mem_AWLEN,
        m_axi_mem_AWSIZE,
        m_axi_mem_AWBURST,
        m_axi_mem_AWLOCK,
        m_axi_mem_AWCACHE,
        m_axi_mem_AWPROT,
        m_axi_mem_AWQOS,
        m_axi_mem_AWREGION,
        m_axi_mem_AWUSER,
        m_axi_mem_WVALID,
        m_axi_mem_WREADY,
        m_axi_mem_WDATA,
        m_axi_mem_WSTRB,
        m_axi_mem_WLAST,
        m_axi_mem_WID,
        m_axi_mem_WUSER,
        m_axi_mem_ARVALID,
        m_axi_mem_ARREADY,
        m_axi_mem_ARADDR,
        m_axi_mem_ARID,
        m_axi_mem_ARLEN,
        m_axi_mem_ARSIZE,
        m_axi_mem_ARBURST,
        m_axi_mem_ARLOCK,
        m_axi_mem_ARCACHE,
        m_axi_mem_ARPROT,
        m_axi_mem_ARQOS,
        m_axi_mem_ARREGION,
        m_axi_mem_ARUSER,
        m_axi_mem_RVALID,
        m_axi_mem_RREADY,
        m_axi_mem_RDATA,
        m_axi_mem_RLAST,
        m_axi_mem_RID,
        m_axi_mem_RUSER,
        m_axi_mem_RRESP,
        m_axi_mem_BVALID,
        m_axi_mem_BREADY,
        m_axi_mem_BRESP,
        m_axi_mem_BID,
        m_axi_mem_BUSER,
        s_axi_cfg_AWVALID,
        s_axi_cfg_AWREADY,
        s_axi_cfg_AWADDR,
        s_axi_cfg_WVALID,
        s_axi_cfg_WREADY,
        s_axi_cfg_WDATA,
        s_axi_cfg_WSTRB,
        s_axi_cfg_ARVALID,
        s_axi_cfg_ARREADY,
        s_axi_cfg_ARADDR,
        s_axi_cfg_RVALID,
        s_axi_cfg_RREADY,
        s_axi_cfg_RDATA,
        s_axi_cfg_RRESP,
        s_axi_cfg_BVALID,
        s_axi_cfg_BREADY,
        s_axi_cfg_BRESP,
        interrupt
);

parameter    ap_ST_fsm_state1 = 107'd1;
parameter    ap_ST_fsm_state2 = 107'd2;
parameter    ap_ST_fsm_state3 = 107'd4;
parameter    ap_ST_fsm_state4 = 107'd8;
parameter    ap_ST_fsm_state5 = 107'd16;
parameter    ap_ST_fsm_state6 = 107'd32;
parameter    ap_ST_fsm_state7 = 107'd64;
parameter    ap_ST_fsm_state8 = 107'd128;
parameter    ap_ST_fsm_state9 = 107'd256;
parameter    ap_ST_fsm_state10 = 107'd512;
parameter    ap_ST_fsm_state11 = 107'd1024;
parameter    ap_ST_fsm_state12 = 107'd2048;
parameter    ap_ST_fsm_state13 = 107'd4096;
parameter    ap_ST_fsm_state14 = 107'd8192;
parameter    ap_ST_fsm_state15 = 107'd16384;
parameter    ap_ST_fsm_state16 = 107'd32768;
parameter    ap_ST_fsm_state17 = 107'd65536;
parameter    ap_ST_fsm_state18 = 107'd131072;
parameter    ap_ST_fsm_state19 = 107'd262144;
parameter    ap_ST_fsm_state20 = 107'd524288;
parameter    ap_ST_fsm_state21 = 107'd1048576;
parameter    ap_ST_fsm_state22 = 107'd2097152;
parameter    ap_ST_fsm_state23 = 107'd4194304;
parameter    ap_ST_fsm_state24 = 107'd8388608;
parameter    ap_ST_fsm_state25 = 107'd16777216;
parameter    ap_ST_fsm_state26 = 107'd33554432;
parameter    ap_ST_fsm_state27 = 107'd67108864;
parameter    ap_ST_fsm_state28 = 107'd134217728;
parameter    ap_ST_fsm_state29 = 107'd268435456;
parameter    ap_ST_fsm_state30 = 107'd536870912;
parameter    ap_ST_fsm_state31 = 107'd1073741824;
parameter    ap_ST_fsm_state32 = 107'd2147483648;
parameter    ap_ST_fsm_state33 = 107'd4294967296;
parameter    ap_ST_fsm_state34 = 107'd8589934592;
parameter    ap_ST_fsm_state35 = 107'd17179869184;
parameter    ap_ST_fsm_state36 = 107'd34359738368;
parameter    ap_ST_fsm_state37 = 107'd68719476736;
parameter    ap_ST_fsm_state38 = 107'd137438953472;
parameter    ap_ST_fsm_state39 = 107'd274877906944;
parameter    ap_ST_fsm_state40 = 107'd549755813888;
parameter    ap_ST_fsm_state41 = 107'd1099511627776;
parameter    ap_ST_fsm_state42 = 107'd2199023255552;
parameter    ap_ST_fsm_state43 = 107'd4398046511104;
parameter    ap_ST_fsm_state44 = 107'd8796093022208;
parameter    ap_ST_fsm_state45 = 107'd17592186044416;
parameter    ap_ST_fsm_state46 = 107'd35184372088832;
parameter    ap_ST_fsm_state47 = 107'd70368744177664;
parameter    ap_ST_fsm_state48 = 107'd140737488355328;
parameter    ap_ST_fsm_state49 = 107'd281474976710656;
parameter    ap_ST_fsm_state50 = 107'd562949953421312;
parameter    ap_ST_fsm_state51 = 107'd1125899906842624;
parameter    ap_ST_fsm_state52 = 107'd2251799813685248;
parameter    ap_ST_fsm_state53 = 107'd4503599627370496;
parameter    ap_ST_fsm_state54 = 107'd9007199254740992;
parameter    ap_ST_fsm_state55 = 107'd18014398509481984;
parameter    ap_ST_fsm_state56 = 107'd36028797018963968;
parameter    ap_ST_fsm_state57 = 107'd72057594037927936;
parameter    ap_ST_fsm_state58 = 107'd144115188075855872;
parameter    ap_ST_fsm_state59 = 107'd288230376151711744;
parameter    ap_ST_fsm_state60 = 107'd576460752303423488;
parameter    ap_ST_fsm_state61 = 107'd1152921504606846976;
parameter    ap_ST_fsm_state62 = 107'd2305843009213693952;
parameter    ap_ST_fsm_state63 = 107'd4611686018427387904;
parameter    ap_ST_fsm_state64 = 107'd9223372036854775808;
parameter    ap_ST_fsm_state65 = 107'd18446744073709551616;
parameter    ap_ST_fsm_state66 = 107'd36893488147419103232;
parameter    ap_ST_fsm_state67 = 107'd73786976294838206464;
parameter    ap_ST_fsm_state68 = 107'd147573952589676412928;
parameter    ap_ST_fsm_state69 = 107'd295147905179352825856;
parameter    ap_ST_fsm_state70 = 107'd590295810358705651712;
parameter    ap_ST_fsm_state71 = 107'd1180591620717411303424;
parameter    ap_ST_fsm_state72 = 107'd2361183241434822606848;
parameter    ap_ST_fsm_state73 = 107'd4722366482869645213696;
parameter    ap_ST_fsm_state74 = 107'd9444732965739290427392;
parameter    ap_ST_fsm_state75 = 107'd18889465931478580854784;
parameter    ap_ST_fsm_state76 = 107'd37778931862957161709568;
parameter    ap_ST_fsm_state77 = 107'd75557863725914323419136;
parameter    ap_ST_fsm_state78 = 107'd151115727451828646838272;
parameter    ap_ST_fsm_state79 = 107'd302231454903657293676544;
parameter    ap_ST_fsm_state80 = 107'd604462909807314587353088;
parameter    ap_ST_fsm_state81 = 107'd1208925819614629174706176;
parameter    ap_ST_fsm_state82 = 107'd2417851639229258349412352;
parameter    ap_ST_fsm_state83 = 107'd4835703278458516698824704;
parameter    ap_ST_fsm_state84 = 107'd9671406556917033397649408;
parameter    ap_ST_fsm_state85 = 107'd19342813113834066795298816;
parameter    ap_ST_fsm_state86 = 107'd38685626227668133590597632;
parameter    ap_ST_fsm_state87 = 107'd77371252455336267181195264;
parameter    ap_ST_fsm_state88 = 107'd154742504910672534362390528;
parameter    ap_ST_fsm_state89 = 107'd309485009821345068724781056;
parameter    ap_ST_fsm_state90 = 107'd618970019642690137449562112;
parameter    ap_ST_fsm_state91 = 107'd1237940039285380274899124224;
parameter    ap_ST_fsm_state92 = 107'd2475880078570760549798248448;
parameter    ap_ST_fsm_state93 = 107'd4951760157141521099596496896;
parameter    ap_ST_fsm_state94 = 107'd9903520314283042199192993792;
parameter    ap_ST_fsm_state95 = 107'd19807040628566084398385987584;
parameter    ap_ST_fsm_state96 = 107'd39614081257132168796771975168;
parameter    ap_ST_fsm_state97 = 107'd79228162514264337593543950336;
parameter    ap_ST_fsm_state98 = 107'd158456325028528675187087900672;
parameter    ap_ST_fsm_state99 = 107'd316912650057057350374175801344;
parameter    ap_ST_fsm_state100 = 107'd633825300114114700748351602688;
parameter    ap_ST_fsm_state101 = 107'd1267650600228229401496703205376;
parameter    ap_ST_fsm_state102 = 107'd2535301200456458802993406410752;
parameter    ap_ST_fsm_state103 = 107'd5070602400912917605986812821504;
parameter    ap_ST_fsm_state104 = 107'd10141204801825835211973625643008;
parameter    ap_ST_fsm_state105 = 107'd20282409603651670423947251286016;
parameter    ap_ST_fsm_state106 = 107'd40564819207303340847894502572032;
parameter    ap_ST_fsm_state107 = 107'd81129638414606681695789005144064;
parameter    C_S_AXI_CFG_DATA_WIDTH = 32;
parameter    C_S_AXI_CFG_ADDR_WIDTH = 8;
parameter    C_S_AXI_DATA_WIDTH = 32;
parameter    C_M_AXI_MEM_ID_WIDTH = 1;
parameter    C_M_AXI_MEM_ADDR_WIDTH = 64;
parameter    C_M_AXI_MEM_DATA_WIDTH = 64;
parameter    C_M_AXI_MEM_AWUSER_WIDTH = 1;
parameter    C_M_AXI_MEM_ARUSER_WIDTH = 1;
parameter    C_M_AXI_MEM_WUSER_WIDTH = 1;
parameter    C_M_AXI_MEM_RUSER_WIDTH = 1;
parameter    C_M_AXI_MEM_BUSER_WIDTH = 1;
parameter    C_M_AXI_MEM_USER_VALUE = 0;
parameter    C_M_AXI_MEM_PROT_VALUE = 0;
parameter    C_M_AXI_MEM_CACHE_VALUE = 3;
parameter    C_M_AXI_DATA_WIDTH = 32;

parameter C_S_AXI_CFG_WSTRB_WIDTH = (32 / 8);
parameter C_S_AXI_WSTRB_WIDTH = (32 / 8);
parameter C_M_AXI_MEM_WSTRB_WIDTH = (64 / 8);
parameter C_M_AXI_WSTRB_WIDTH = (32 / 8);

input   ap_clk;
input   ap_rst_n;
output   m_axi_mem_AWVALID;
input   m_axi_mem_AWREADY;
output  [C_M_AXI_MEM_ADDR_WIDTH - 1:0] m_axi_mem_AWADDR;
output  [C_M_AXI_MEM_ID_WIDTH - 1:0] m_axi_mem_AWID;
output  [7:0] m_axi_mem_AWLEN;
output  [2:0] m_axi_mem_AWSIZE;
output  [1:0] m_axi_mem_AWBURST;
output  [1:0] m_axi_mem_AWLOCK;
output  [3:0] m_axi_mem_AWCACHE;
output  [2:0] m_axi_mem_AWPROT;
output  [3:0] m_axi_mem_AWQOS;
output  [3:0] m_axi_mem_AWREGION;
output  [C_M_AXI_MEM_AWUSER_WIDTH - 1:0] m_axi_mem_AWUSER;
output   m_axi_mem_WVALID;
input   m_axi_mem_WREADY;
output  [C_M_AXI_MEM_DATA_WIDTH - 1:0] m_axi_mem_WDATA;
output  [C_M_AXI_MEM_WSTRB_WIDTH - 1:0] m_axi_mem_WSTRB;
output   m_axi_mem_WLAST;
output  [C_M_AXI_MEM_ID_WIDTH - 1:0] m_axi_mem_WID;
output  [C_M_AXI_MEM_WUSER_WIDTH - 1:0] m_axi_mem_WUSER;
output   m_axi_mem_ARVALID;
input   m_axi_mem_ARREADY;
output  [C_M_AXI_MEM_ADDR_WIDTH - 1:0] m_axi_mem_ARADDR;
output  [C_M_AXI_MEM_ID_WIDTH - 1:0] m_axi_mem_ARID;
output  [7:0] m_axi_mem_ARLEN;
output  [2:0] m_axi_mem_ARSIZE;
output  [1:0] m_axi_mem_ARBURST;
output  [1:0] m_axi_mem_ARLOCK;
output  [3:0] m_axi_mem_ARCACHE;
output  [2:0] m_axi_mem_ARPROT;
output  [3:0] m_axi_mem_ARQOS;
output  [3:0] m_axi_mem_ARREGION;
output  [C_M_AXI_MEM_ARUSER_WIDTH - 1:0] m_axi_mem_ARUSER;
input   m_axi_mem_RVALID;
output   m_axi_mem_RREADY;
input  [C_M_AXI_MEM_DATA_WIDTH - 1:0] m_axi_mem_RDATA;
input   m_axi_mem_RLAST;
input  [C_M_AXI_MEM_ID_WIDTH - 1:0] m_axi_mem_RID;
input  [C_M_AXI_MEM_RUSER_WIDTH - 1:0] m_axi_mem_RUSER;
input  [1:0] m_axi_mem_RRESP;
input   m_axi_mem_BVALID;
output   m_axi_mem_BREADY;
input  [1:0] m_axi_mem_BRESP;
input  [C_M_AXI_MEM_ID_WIDTH - 1:0] m_axi_mem_BID;
input  [C_M_AXI_MEM_BUSER_WIDTH - 1:0] m_axi_mem_BUSER;
input   s_axi_cfg_AWVALID;
output   s_axi_cfg_AWREADY;
input  [C_S_AXI_CFG_ADDR_WIDTH - 1:0] s_axi_cfg_AWADDR;
input   s_axi_cfg_WVALID;
output   s_axi_cfg_WREADY;
input  [C_S_AXI_CFG_DATA_WIDTH - 1:0] s_axi_cfg_WDATA;
input  [C_S_AXI_CFG_WSTRB_WIDTH - 1:0] s_axi_cfg_WSTRB;
input   s_axi_cfg_ARVALID;
output   s_axi_cfg_ARREADY;
input  [C_S_AXI_CFG_ADDR_WIDTH - 1:0] s_axi_cfg_ARADDR;
output   s_axi_cfg_RVALID;
input   s_axi_cfg_RREADY;
output  [C_S_AXI_CFG_DATA_WIDTH - 1:0] s_axi_cfg_RDATA;
output  [1:0] s_axi_cfg_RRESP;
output   s_axi_cfg_BVALID;
input   s_axi_cfg_BREADY;
output  [1:0] s_axi_cfg_BRESP;
output   interrupt;

 reg    ap_rst_n_inv;
wire    ap_start;
reg    ap_done;
reg    ap_idle;
(* fsm_encoding = "none" *) reg   [106:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg    ap_ready;
wire   [31:0] n;
wire   [31:0] k;
wire   [31:0] control;
wire   [63:0] buf_ptr_node_x_coords;
wire   [63:0] buf_ptr_node_y_coords;
wire   [63:0] buf_ptr_node_cluster_assignments;
wire   [63:0] buf_ptr_centroid_x_coords;
wire   [63:0] buf_ptr_centroid_y_coords;
wire   [63:0] buf_ptr_intermediate_cluster_assignments;
wire   [63:0] buf_ptr_intermediate_centroid_x_coords;
wire   [63:0] buf_ptr_intermediate_centroid_y_coords;
wire   [63:0] max_iterations;
wire   [63:0] sub_iterations;
reg    mem_blk_n_AR;
wire    ap_CS_fsm_state2;
reg   [0:0] icmp_ln185_reg_1059;
wire    ap_CS_fsm_state11;
wire    ap_CS_fsm_state20;
wire    ap_CS_fsm_state29;
wire    ap_CS_fsm_state38;
reg    mem_blk_n_AW;
wire    ap_CS_fsm_state49;
reg    mem_blk_n_B;
wire    ap_CS_fsm_state56;
reg   [0:0] tmp_reg_1161;
reg   [0:0] icmp_ln196_reg_1165;
wire    ap_CS_fsm_state57;
wire    ap_CS_fsm_state64;
wire    ap_CS_fsm_state71;
reg   [0:0] icmp_ln188_reg_1095;
reg   [0:0] trunc_ln199_reg_1180;
reg   [0:0] icmp_ln199_reg_1184;
wire    ap_CS_fsm_state72;
wire    ap_CS_fsm_state79;
wire    ap_CS_fsm_state86;
reg   [0:0] tmp_3_reg_1152;
wire   [0:0] grp_fu_576_p3;
wire    ap_CS_fsm_state93;
reg   [0:0] tmp_4_reg_1220;
wire   [0:0] trunc_ln215_fu_943_p1;
wire    ap_CS_fsm_state100;
wire    ap_CS_fsm_state107;
reg   [0:0] trunc_ln215_reg_1229;
wire  signed [60:0] grp_fu_518_p4;
reg   [60:0] reg_590;
wire    ap_CS_fsm_state47;
wire   [0:0] icmp_ln191_fu_738_p2;
wire   [0:0] tmp_3_fu_782_p3;
wire   [0:0] ap_phi_mux_phi_ln191_phi_fu_374_p4;
wire  signed [60:0] grp_fu_527_p4;
reg   [60:0] reg_596;
wire  signed [60:0] grp_fu_536_p4;
reg   [60:0] reg_602;
wire  signed [60:0] grp_fu_545_p4;
reg   [60:0] reg_608;
wire  signed [60:0] grp_fu_554_p4;
reg   [60:0] reg_614;
reg   [63:0] buf_ptr_intermediate_centroid_y_coords_read_reg_969;
reg   [63:0] buf_ptr_intermediate_centroid_x_coords_read_reg_974;
reg   [63:0] buf_ptr_intermediate_cluster_assignments_read_reg_979;
reg   [63:0] buf_ptr_centroid_y_coords_read_reg_984;
reg   [63:0] buf_ptr_centroid_x_coords_read_reg_989;
reg   [63:0] buf_ptr_node_cluster_assignments_read_reg_994;
reg   [63:0] buf_ptr_node_y_coords_read_reg_999;
reg   [63:0] buf_ptr_node_x_coords_read_reg_1004;
reg   [31:0] grp_load_fu_510_p1;
reg   [31:0] n_assign_load_reg_1041;
wire   [0:0] icmp_ln185_fu_649_p2;
reg   [31:0] k_assign_load_reg_1063;
wire   [0:0] icmp_ln188_fu_688_p2;
wire    ap_CS_fsm_state28;
wire   [31:0] intermediate_writes_made_2_fu_728_p2;
reg   [31:0] intermediate_writes_made_2_reg_1123;
reg   [63:0] sub_iterations_assign_load_reg_1131;
reg   [31:0] n_assign_load_1_reg_1136;
reg   [31:0] k_assign_load_1_reg_1141;
wire   [28:0] mul_ln194_fu_776_p2;
reg   [28:0] mul_ln194_reg_1146;
wire   [0:0] grp_kmeans_fu_426_ap_return;
reg   [0:0] converged_reg_1156;
wire    ap_CS_fsm_state48;
wire   [0:0] grp_fu_584_p2;
reg   [60:0] p_cast9_reg_1169;
wire   [0:0] trunc_ln199_fu_826_p1;
reg   [60:0] p_cast10_reg_1188;
reg   [60:0] p_cast11_reg_1194;
reg   [12:0] node_x_coords_address0;
reg    node_x_coords_ce0;
wire   [63:0] node_x_coords_q0;
reg   [12:0] node_x_coords_address1;
reg    node_x_coords_ce1;
reg    node_x_coords_we1;
wire   [63:0] node_x_coords_q1;
reg   [12:0] node_y_coords_address0;
reg    node_y_coords_ce0;
wire   [63:0] node_y_coords_q0;
reg   [12:0] node_y_coords_address1;
reg    node_y_coords_ce1;
reg    node_y_coords_we1;
wire   [63:0] node_y_coords_q1;
reg   [12:0] node_cluster_assignments_address0;
reg    node_cluster_assignments_ce0;
wire   [63:0] node_cluster_assignments_q0;
reg   [12:0] node_cluster_assignments_address1;
reg    node_cluster_assignments_ce1;
reg    node_cluster_assignments_we1;
reg   [63:0] node_cluster_assignments_d1;
reg   [7:0] centroid_x_coords_address0;
reg    centroid_x_coords_ce0;
reg    centroid_x_coords_we0;
reg   [63:0] centroid_x_coords_d0;
wire   [63:0] centroid_x_coords_q0;
reg    centroid_x_coords_ce1;
wire   [63:0] centroid_x_coords_q1;
reg   [7:0] centroid_y_coords_address0;
reg    centroid_y_coords_ce0;
reg    centroid_y_coords_we0;
reg   [63:0] centroid_y_coords_d0;
wire   [63:0] centroid_y_coords_q0;
reg    centroid_y_coords_ce1;
wire   [63:0] centroid_y_coords_q1;
wire    grp_kmeans_top_Pipeline_1_fu_381_ap_start;
wire    grp_kmeans_top_Pipeline_1_fu_381_ap_done;
wire    grp_kmeans_top_Pipeline_1_fu_381_ap_idle;
wire    grp_kmeans_top_Pipeline_1_fu_381_ap_ready;
wire    grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_AWVALID;
wire   [63:0] grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_AWADDR;
wire   [0:0] grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_AWID;
wire   [31:0] grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_AWLEN;
wire   [2:0] grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_AWSIZE;
wire   [1:0] grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_AWBURST;
wire   [1:0] grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_AWLOCK;
wire   [3:0] grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_AWCACHE;
wire   [2:0] grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_AWPROT;
wire   [3:0] grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_AWQOS;
wire   [3:0] grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_AWREGION;
wire   [0:0] grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_AWUSER;
wire    grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_WVALID;
wire   [63:0] grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_WDATA;
wire   [7:0] grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_WSTRB;
wire    grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_WLAST;
wire   [0:0] grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_WID;
wire   [0:0] grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_WUSER;
wire    grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_ARVALID;
wire   [63:0] grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_ARADDR;
wire   [0:0] grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_ARID;
wire   [31:0] grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_ARLEN;
wire   [2:0] grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_ARSIZE;
wire   [1:0] grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_ARBURST;
wire   [1:0] grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_ARLOCK;
wire   [3:0] grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_ARCACHE;
wire   [2:0] grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_ARPROT;
wire   [3:0] grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_ARQOS;
wire   [3:0] grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_ARREGION;
wire   [0:0] grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_ARUSER;
wire    grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_RREADY;
wire    grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_BREADY;
wire   [12:0] grp_kmeans_top_Pipeline_1_fu_381_node_x_coords_address1;
wire    grp_kmeans_top_Pipeline_1_fu_381_node_x_coords_ce1;
wire    grp_kmeans_top_Pipeline_1_fu_381_node_x_coords_we1;
wire   [63:0] grp_kmeans_top_Pipeline_1_fu_381_node_x_coords_d1;
wire    grp_kmeans_top_Pipeline_2_fu_390_ap_start;
wire    grp_kmeans_top_Pipeline_2_fu_390_ap_done;
wire    grp_kmeans_top_Pipeline_2_fu_390_ap_idle;
wire    grp_kmeans_top_Pipeline_2_fu_390_ap_ready;
wire    grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_AWVALID;
wire   [63:0] grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_AWADDR;
wire   [0:0] grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_AWID;
wire   [31:0] grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_AWLEN;
wire   [2:0] grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_AWSIZE;
wire   [1:0] grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_AWBURST;
wire   [1:0] grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_AWLOCK;
wire   [3:0] grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_AWCACHE;
wire   [2:0] grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_AWPROT;
wire   [3:0] grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_AWQOS;
wire   [3:0] grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_AWREGION;
wire   [0:0] grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_AWUSER;
wire    grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_WVALID;
wire   [63:0] grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_WDATA;
wire   [7:0] grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_WSTRB;
wire    grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_WLAST;
wire   [0:0] grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_WID;
wire   [0:0] grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_WUSER;
wire    grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_ARVALID;
wire   [63:0] grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_ARADDR;
wire   [0:0] grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_ARID;
wire   [31:0] grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_ARLEN;
wire   [2:0] grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_ARSIZE;
wire   [1:0] grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_ARBURST;
wire   [1:0] grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_ARLOCK;
wire   [3:0] grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_ARCACHE;
wire   [2:0] grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_ARPROT;
wire   [3:0] grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_ARQOS;
wire   [3:0] grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_ARREGION;
wire   [0:0] grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_ARUSER;
wire    grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_RREADY;
wire    grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_BREADY;
wire   [12:0] grp_kmeans_top_Pipeline_2_fu_390_node_y_coords_address1;
wire    grp_kmeans_top_Pipeline_2_fu_390_node_y_coords_ce1;
wire    grp_kmeans_top_Pipeline_2_fu_390_node_y_coords_we1;
wire   [63:0] grp_kmeans_top_Pipeline_2_fu_390_node_y_coords_d1;
wire    grp_kmeans_top_Pipeline_3_fu_399_ap_start;
wire    grp_kmeans_top_Pipeline_3_fu_399_ap_done;
wire    grp_kmeans_top_Pipeline_3_fu_399_ap_idle;
wire    grp_kmeans_top_Pipeline_3_fu_399_ap_ready;
wire    grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_AWVALID;
wire   [63:0] grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_AWADDR;
wire   [0:0] grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_AWID;
wire   [31:0] grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_AWLEN;
wire   [2:0] grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_AWSIZE;
wire   [1:0] grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_AWBURST;
wire   [1:0] grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_AWLOCK;
wire   [3:0] grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_AWCACHE;
wire   [2:0] grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_AWPROT;
wire   [3:0] grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_AWQOS;
wire   [3:0] grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_AWREGION;
wire   [0:0] grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_AWUSER;
wire    grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_WVALID;
wire   [63:0] grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_WDATA;
wire   [7:0] grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_WSTRB;
wire    grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_WLAST;
wire   [0:0] grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_WID;
wire   [0:0] grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_WUSER;
wire    grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_ARVALID;
wire   [63:0] grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_ARADDR;
wire   [0:0] grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_ARID;
wire   [31:0] grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_ARLEN;
wire   [2:0] grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_ARSIZE;
wire   [1:0] grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_ARBURST;
wire   [1:0] grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_ARLOCK;
wire   [3:0] grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_ARCACHE;
wire   [2:0] grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_ARPROT;
wire   [3:0] grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_ARQOS;
wire   [3:0] grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_ARREGION;
wire   [0:0] grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_ARUSER;
wire    grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_RREADY;
wire    grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_BREADY;
wire   [12:0] grp_kmeans_top_Pipeline_3_fu_399_node_cluster_assignments_address1;
wire    grp_kmeans_top_Pipeline_3_fu_399_node_cluster_assignments_ce1;
wire    grp_kmeans_top_Pipeline_3_fu_399_node_cluster_assignments_we1;
wire   [63:0] grp_kmeans_top_Pipeline_3_fu_399_node_cluster_assignments_d1;
wire    grp_kmeans_top_Pipeline_4_fu_408_ap_start;
wire    grp_kmeans_top_Pipeline_4_fu_408_ap_done;
wire    grp_kmeans_top_Pipeline_4_fu_408_ap_idle;
wire    grp_kmeans_top_Pipeline_4_fu_408_ap_ready;
wire    grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_AWVALID;
wire   [63:0] grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_AWADDR;
wire   [0:0] grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_AWID;
wire   [31:0] grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_AWLEN;
wire   [2:0] grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_AWSIZE;
wire   [1:0] grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_AWBURST;
wire   [1:0] grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_AWLOCK;
wire   [3:0] grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_AWCACHE;
wire   [2:0] grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_AWPROT;
wire   [3:0] grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_AWQOS;
wire   [3:0] grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_AWREGION;
wire   [0:0] grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_AWUSER;
wire    grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_WVALID;
wire   [63:0] grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_WDATA;
wire   [7:0] grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_WSTRB;
wire    grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_WLAST;
wire   [0:0] grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_WID;
wire   [0:0] grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_WUSER;
wire    grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_ARVALID;
wire   [63:0] grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_ARADDR;
wire   [0:0] grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_ARID;
wire   [31:0] grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_ARLEN;
wire   [2:0] grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_ARSIZE;
wire   [1:0] grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_ARBURST;
wire   [1:0] grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_ARLOCK;
wire   [3:0] grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_ARCACHE;
wire   [2:0] grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_ARPROT;
wire   [3:0] grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_ARQOS;
wire   [3:0] grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_ARREGION;
wire   [0:0] grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_ARUSER;
wire    grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_RREADY;
wire    grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_BREADY;
wire   [7:0] grp_kmeans_top_Pipeline_4_fu_408_centroid_x_coords_address0;
wire    grp_kmeans_top_Pipeline_4_fu_408_centroid_x_coords_ce0;
wire    grp_kmeans_top_Pipeline_4_fu_408_centroid_x_coords_we0;
wire   [63:0] grp_kmeans_top_Pipeline_4_fu_408_centroid_x_coords_d0;
wire    grp_kmeans_top_Pipeline_5_fu_417_ap_start;
wire    grp_kmeans_top_Pipeline_5_fu_417_ap_done;
wire    grp_kmeans_top_Pipeline_5_fu_417_ap_idle;
wire    grp_kmeans_top_Pipeline_5_fu_417_ap_ready;
wire    grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_AWVALID;
wire   [63:0] grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_AWADDR;
wire   [0:0] grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_AWID;
wire   [31:0] grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_AWLEN;
wire   [2:0] grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_AWSIZE;
wire   [1:0] grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_AWBURST;
wire   [1:0] grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_AWLOCK;
wire   [3:0] grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_AWCACHE;
wire   [2:0] grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_AWPROT;
wire   [3:0] grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_AWQOS;
wire   [3:0] grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_AWREGION;
wire   [0:0] grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_AWUSER;
wire    grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_WVALID;
wire   [63:0] grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_WDATA;
wire   [7:0] grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_WSTRB;
wire    grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_WLAST;
wire   [0:0] grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_WID;
wire   [0:0] grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_WUSER;
wire    grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_ARVALID;
wire   [63:0] grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_ARADDR;
wire   [0:0] grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_ARID;
wire   [31:0] grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_ARLEN;
wire   [2:0] grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_ARSIZE;
wire   [1:0] grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_ARBURST;
wire   [1:0] grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_ARLOCK;
wire   [3:0] grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_ARCACHE;
wire   [2:0] grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_ARPROT;
wire   [3:0] grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_ARQOS;
wire   [3:0] grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_ARREGION;
wire   [0:0] grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_ARUSER;
wire    grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_RREADY;
wire    grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_BREADY;
wire   [7:0] grp_kmeans_top_Pipeline_5_fu_417_centroid_y_coords_address0;
wire    grp_kmeans_top_Pipeline_5_fu_417_centroid_y_coords_ce0;
wire    grp_kmeans_top_Pipeline_5_fu_417_centroid_y_coords_we0;
wire   [63:0] grp_kmeans_top_Pipeline_5_fu_417_centroid_y_coords_d0;
wire    grp_kmeans_fu_426_ap_start;
wire    grp_kmeans_fu_426_ap_done;
wire    grp_kmeans_fu_426_ap_idle;
wire    grp_kmeans_fu_426_ap_ready;
wire   [12:0] grp_kmeans_fu_426_node_x_coords_address0;
wire    grp_kmeans_fu_426_node_x_coords_ce0;
wire   [12:0] grp_kmeans_fu_426_node_x_coords_address1;
wire    grp_kmeans_fu_426_node_x_coords_ce1;
wire   [12:0] grp_kmeans_fu_426_node_y_coords_address0;
wire    grp_kmeans_fu_426_node_y_coords_ce0;
wire   [12:0] grp_kmeans_fu_426_node_y_coords_address1;
wire    grp_kmeans_fu_426_node_y_coords_ce1;
wire   [12:0] grp_kmeans_fu_426_node_cluster_assignments_address1;
wire    grp_kmeans_fu_426_node_cluster_assignments_ce1;
wire    grp_kmeans_fu_426_node_cluster_assignments_we1;
wire   [63:0] grp_kmeans_fu_426_node_cluster_assignments_d1;
wire   [7:0] grp_kmeans_fu_426_centroid_x_coords_address0;
wire    grp_kmeans_fu_426_centroid_x_coords_ce0;
wire    grp_kmeans_fu_426_centroid_x_coords_we0;
wire   [63:0] grp_kmeans_fu_426_centroid_x_coords_d0;
wire   [7:0] grp_kmeans_fu_426_centroid_x_coords_address1;
wire    grp_kmeans_fu_426_centroid_x_coords_ce1;
wire   [7:0] grp_kmeans_fu_426_centroid_y_coords_address0;
wire    grp_kmeans_fu_426_centroid_y_coords_ce0;
wire    grp_kmeans_fu_426_centroid_y_coords_we0;
wire   [63:0] grp_kmeans_fu_426_centroid_y_coords_d0;
wire   [7:0] grp_kmeans_fu_426_centroid_y_coords_address1;
wire    grp_kmeans_fu_426_centroid_y_coords_ce1;
wire    grp_kmeans_top_Pipeline_6_fu_438_ap_start;
wire    grp_kmeans_top_Pipeline_6_fu_438_ap_done;
wire    grp_kmeans_top_Pipeline_6_fu_438_ap_idle;
wire    grp_kmeans_top_Pipeline_6_fu_438_ap_ready;
wire    grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_AWVALID;
wire   [63:0] grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_AWADDR;
wire   [0:0] grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_AWID;
wire   [31:0] grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_AWLEN;
wire   [2:0] grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_AWSIZE;
wire   [1:0] grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_AWBURST;
wire   [1:0] grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_AWLOCK;
wire   [3:0] grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_AWCACHE;
wire   [2:0] grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_AWPROT;
wire   [3:0] grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_AWQOS;
wire   [3:0] grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_AWREGION;
wire   [0:0] grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_AWUSER;
wire    grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_WVALID;
wire   [63:0] grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_WDATA;
wire   [7:0] grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_WSTRB;
wire    grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_WLAST;
wire   [0:0] grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_WID;
wire   [0:0] grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_WUSER;
wire    grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_ARVALID;
wire   [63:0] grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_ARADDR;
wire   [0:0] grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_ARID;
wire   [31:0] grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_ARLEN;
wire   [2:0] grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_ARSIZE;
wire   [1:0] grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_ARBURST;
wire   [1:0] grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_ARLOCK;
wire   [3:0] grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_ARCACHE;
wire   [2:0] grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_ARPROT;
wire   [3:0] grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_ARQOS;
wire   [3:0] grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_ARREGION;
wire   [0:0] grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_ARUSER;
wire    grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_RREADY;
wire    grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_BREADY;
wire   [12:0] grp_kmeans_top_Pipeline_6_fu_438_node_cluster_assignments_address0;
wire    grp_kmeans_top_Pipeline_6_fu_438_node_cluster_assignments_ce0;
wire    grp_kmeans_top_Pipeline_7_fu_447_ap_start;
wire    grp_kmeans_top_Pipeline_7_fu_447_ap_done;
wire    grp_kmeans_top_Pipeline_7_fu_447_ap_idle;
wire    grp_kmeans_top_Pipeline_7_fu_447_ap_ready;
wire    grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_AWVALID;
wire   [63:0] grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_AWADDR;
wire   [0:0] grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_AWID;
wire   [31:0] grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_AWLEN;
wire   [2:0] grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_AWSIZE;
wire   [1:0] grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_AWBURST;
wire   [1:0] grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_AWLOCK;
wire   [3:0] grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_AWCACHE;
wire   [2:0] grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_AWPROT;
wire   [3:0] grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_AWQOS;
wire   [3:0] grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_AWREGION;
wire   [0:0] grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_AWUSER;
wire    grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_WVALID;
wire   [63:0] grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_WDATA;
wire   [7:0] grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_WSTRB;
wire    grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_WLAST;
wire   [0:0] grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_WID;
wire   [0:0] grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_WUSER;
wire    grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_ARVALID;
wire   [63:0] grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_ARADDR;
wire   [0:0] grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_ARID;
wire   [31:0] grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_ARLEN;
wire   [2:0] grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_ARSIZE;
wire   [1:0] grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_ARBURST;
wire   [1:0] grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_ARLOCK;
wire   [3:0] grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_ARCACHE;
wire   [2:0] grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_ARPROT;
wire   [3:0] grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_ARQOS;
wire   [3:0] grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_ARREGION;
wire   [0:0] grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_ARUSER;
wire    grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_RREADY;
wire    grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_BREADY;
wire   [7:0] grp_kmeans_top_Pipeline_7_fu_447_centroid_x_coords_address0;
wire    grp_kmeans_top_Pipeline_7_fu_447_centroid_x_coords_ce0;
wire    grp_kmeans_top_Pipeline_8_fu_456_ap_start;
wire    grp_kmeans_top_Pipeline_8_fu_456_ap_done;
wire    grp_kmeans_top_Pipeline_8_fu_456_ap_idle;
wire    grp_kmeans_top_Pipeline_8_fu_456_ap_ready;
wire    grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_AWVALID;
wire   [63:0] grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_AWADDR;
wire   [0:0] grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_AWID;
wire   [31:0] grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_AWLEN;
wire   [2:0] grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_AWSIZE;
wire   [1:0] grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_AWBURST;
wire   [1:0] grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_AWLOCK;
wire   [3:0] grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_AWCACHE;
wire   [2:0] grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_AWPROT;
wire   [3:0] grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_AWQOS;
wire   [3:0] grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_AWREGION;
wire   [0:0] grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_AWUSER;
wire    grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_WVALID;
wire   [63:0] grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_WDATA;
wire   [7:0] grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_WSTRB;
wire    grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_WLAST;
wire   [0:0] grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_WID;
wire   [0:0] grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_WUSER;
wire    grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_ARVALID;
wire   [63:0] grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_ARADDR;
wire   [0:0] grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_ARID;
wire   [31:0] grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_ARLEN;
wire   [2:0] grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_ARSIZE;
wire   [1:0] grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_ARBURST;
wire   [1:0] grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_ARLOCK;
wire   [3:0] grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_ARCACHE;
wire   [2:0] grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_ARPROT;
wire   [3:0] grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_ARQOS;
wire   [3:0] grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_ARREGION;
wire   [0:0] grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_ARUSER;
wire    grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_RREADY;
wire    grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_BREADY;
wire   [7:0] grp_kmeans_top_Pipeline_8_fu_456_centroid_y_coords_address0;
wire    grp_kmeans_top_Pipeline_8_fu_456_centroid_y_coords_ce0;
wire    grp_kmeans_top_Pipeline_9_fu_465_ap_start;
wire    grp_kmeans_top_Pipeline_9_fu_465_ap_done;
wire    grp_kmeans_top_Pipeline_9_fu_465_ap_idle;
wire    grp_kmeans_top_Pipeline_9_fu_465_ap_ready;
wire    grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_AWVALID;
wire   [63:0] grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_AWADDR;
wire   [0:0] grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_AWID;
wire   [31:0] grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_AWLEN;
wire   [2:0] grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_AWSIZE;
wire   [1:0] grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_AWBURST;
wire   [1:0] grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_AWLOCK;
wire   [3:0] grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_AWCACHE;
wire   [2:0] grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_AWPROT;
wire   [3:0] grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_AWQOS;
wire   [3:0] grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_AWREGION;
wire   [0:0] grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_AWUSER;
wire    grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_WVALID;
wire   [63:0] grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_WDATA;
wire   [7:0] grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_WSTRB;
wire    grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_WLAST;
wire   [0:0] grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_WID;
wire   [0:0] grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_WUSER;
wire    grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_ARVALID;
wire   [63:0] grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_ARADDR;
wire   [0:0] grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_ARID;
wire   [31:0] grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_ARLEN;
wire   [2:0] grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_ARSIZE;
wire   [1:0] grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_ARBURST;
wire   [1:0] grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_ARLOCK;
wire   [3:0] grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_ARCACHE;
wire   [2:0] grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_ARPROT;
wire   [3:0] grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_ARQOS;
wire   [3:0] grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_ARREGION;
wire   [0:0] grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_ARUSER;
wire    grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_RREADY;
wire    grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_BREADY;
wire   [12:0] grp_kmeans_top_Pipeline_9_fu_465_node_x_coords_address0;
wire    grp_kmeans_top_Pipeline_9_fu_465_node_x_coords_ce0;
wire    grp_kmeans_top_Pipeline_10_fu_474_ap_start;
wire    grp_kmeans_top_Pipeline_10_fu_474_ap_done;
wire    grp_kmeans_top_Pipeline_10_fu_474_ap_idle;
wire    grp_kmeans_top_Pipeline_10_fu_474_ap_ready;
wire    grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_AWVALID;
wire   [63:0] grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_AWADDR;
wire   [0:0] grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_AWID;
wire   [31:0] grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_AWLEN;
wire   [2:0] grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_AWSIZE;
wire   [1:0] grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_AWBURST;
wire   [1:0] grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_AWLOCK;
wire   [3:0] grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_AWCACHE;
wire   [2:0] grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_AWPROT;
wire   [3:0] grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_AWQOS;
wire   [3:0] grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_AWREGION;
wire   [0:0] grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_AWUSER;
wire    grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_WVALID;
wire   [63:0] grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_WDATA;
wire   [7:0] grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_WSTRB;
wire    grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_WLAST;
wire   [0:0] grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_WID;
wire   [0:0] grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_WUSER;
wire    grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_ARVALID;
wire   [63:0] grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_ARADDR;
wire   [0:0] grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_ARID;
wire   [31:0] grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_ARLEN;
wire   [2:0] grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_ARSIZE;
wire   [1:0] grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_ARBURST;
wire   [1:0] grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_ARLOCK;
wire   [3:0] grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_ARCACHE;
wire   [2:0] grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_ARPROT;
wire   [3:0] grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_ARQOS;
wire   [3:0] grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_ARREGION;
wire   [0:0] grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_ARUSER;
wire    grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_RREADY;
wire    grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_BREADY;
wire   [12:0] grp_kmeans_top_Pipeline_10_fu_474_node_y_coords_address0;
wire    grp_kmeans_top_Pipeline_10_fu_474_node_y_coords_ce0;
wire    grp_kmeans_top_Pipeline_11_fu_483_ap_start;
wire    grp_kmeans_top_Pipeline_11_fu_483_ap_done;
wire    grp_kmeans_top_Pipeline_11_fu_483_ap_idle;
wire    grp_kmeans_top_Pipeline_11_fu_483_ap_ready;
wire    grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_AWVALID;
wire   [63:0] grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_AWADDR;
wire   [0:0] grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_AWID;
wire   [31:0] grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_AWLEN;
wire   [2:0] grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_AWSIZE;
wire   [1:0] grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_AWBURST;
wire   [1:0] grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_AWLOCK;
wire   [3:0] grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_AWCACHE;
wire   [2:0] grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_AWPROT;
wire   [3:0] grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_AWQOS;
wire   [3:0] grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_AWREGION;
wire   [0:0] grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_AWUSER;
wire    grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_WVALID;
wire   [63:0] grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_WDATA;
wire   [7:0] grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_WSTRB;
wire    grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_WLAST;
wire   [0:0] grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_WID;
wire   [0:0] grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_WUSER;
wire    grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_ARVALID;
wire   [63:0] grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_ARADDR;
wire   [0:0] grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_ARID;
wire   [31:0] grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_ARLEN;
wire   [2:0] grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_ARSIZE;
wire   [1:0] grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_ARBURST;
wire   [1:0] grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_ARLOCK;
wire   [3:0] grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_ARCACHE;
wire   [2:0] grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_ARPROT;
wire   [3:0] grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_ARQOS;
wire   [3:0] grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_ARREGION;
wire   [0:0] grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_ARUSER;
wire    grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_RREADY;
wire    grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_BREADY;
wire   [12:0] grp_kmeans_top_Pipeline_11_fu_483_node_cluster_assignments_address0;
wire    grp_kmeans_top_Pipeline_11_fu_483_node_cluster_assignments_ce0;
wire    grp_kmeans_top_Pipeline_12_fu_492_ap_start;
wire    grp_kmeans_top_Pipeline_12_fu_492_ap_done;
wire    grp_kmeans_top_Pipeline_12_fu_492_ap_idle;
wire    grp_kmeans_top_Pipeline_12_fu_492_ap_ready;
wire    grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_AWVALID;
wire   [63:0] grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_AWADDR;
wire   [0:0] grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_AWID;
wire   [31:0] grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_AWLEN;
wire   [2:0] grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_AWSIZE;
wire   [1:0] grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_AWBURST;
wire   [1:0] grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_AWLOCK;
wire   [3:0] grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_AWCACHE;
wire   [2:0] grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_AWPROT;
wire   [3:0] grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_AWQOS;
wire   [3:0] grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_AWREGION;
wire   [0:0] grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_AWUSER;
wire    grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_WVALID;
wire   [63:0] grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_WDATA;
wire   [7:0] grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_WSTRB;
wire    grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_WLAST;
wire   [0:0] grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_WID;
wire   [0:0] grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_WUSER;
wire    grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_ARVALID;
wire   [63:0] grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_ARADDR;
wire   [0:0] grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_ARID;
wire   [31:0] grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_ARLEN;
wire   [2:0] grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_ARSIZE;
wire   [1:0] grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_ARBURST;
wire   [1:0] grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_ARLOCK;
wire   [3:0] grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_ARCACHE;
wire   [2:0] grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_ARPROT;
wire   [3:0] grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_ARQOS;
wire   [3:0] grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_ARREGION;
wire   [0:0] grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_ARUSER;
wire    grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_RREADY;
wire    grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_BREADY;
wire   [7:0] grp_kmeans_top_Pipeline_12_fu_492_centroid_x_coords_address0;
wire    grp_kmeans_top_Pipeline_12_fu_492_centroid_x_coords_ce0;
wire    grp_kmeans_top_Pipeline_13_fu_501_ap_start;
wire    grp_kmeans_top_Pipeline_13_fu_501_ap_done;
wire    grp_kmeans_top_Pipeline_13_fu_501_ap_idle;
wire    grp_kmeans_top_Pipeline_13_fu_501_ap_ready;
wire    grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_AWVALID;
wire   [63:0] grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_AWADDR;
wire   [0:0] grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_AWID;
wire   [31:0] grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_AWLEN;
wire   [2:0] grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_AWSIZE;
wire   [1:0] grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_AWBURST;
wire   [1:0] grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_AWLOCK;
wire   [3:0] grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_AWCACHE;
wire   [2:0] grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_AWPROT;
wire   [3:0] grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_AWQOS;
wire   [3:0] grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_AWREGION;
wire   [0:0] grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_AWUSER;
wire    grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_WVALID;
wire   [63:0] grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_WDATA;
wire   [7:0] grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_WSTRB;
wire    grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_WLAST;
wire   [0:0] grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_WID;
wire   [0:0] grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_WUSER;
wire    grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_ARVALID;
wire   [63:0] grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_ARADDR;
wire   [0:0] grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_ARID;
wire   [31:0] grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_ARLEN;
wire   [2:0] grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_ARSIZE;
wire   [1:0] grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_ARBURST;
wire   [1:0] grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_ARLOCK;
wire   [3:0] grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_ARCACHE;
wire   [2:0] grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_ARPROT;
wire   [3:0] grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_ARQOS;
wire   [3:0] grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_ARREGION;
wire   [0:0] grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_ARUSER;
wire    grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_RREADY;
wire    grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_BREADY;
wire   [7:0] grp_kmeans_top_Pipeline_13_fu_501_centroid_y_coords_address0;
wire    grp_kmeans_top_Pipeline_13_fu_501_centroid_y_coords_ce0;
reg    mem_AWVALID;
wire    mem_AWREADY;
reg   [63:0] mem_AWADDR;
reg   [31:0] mem_AWLEN;
reg    mem_WVALID;
wire    mem_WREADY;
reg   [63:0] mem_WDATA;
reg   [7:0] mem_WSTRB;
reg    mem_ARVALID;
wire    mem_ARREADY;
reg   [63:0] mem_ARADDR;
reg   [31:0] mem_ARLEN;
wire    mem_RVALID;
reg    mem_RREADY;
wire   [63:0] mem_RDATA;
wire   [8:0] mem_RFIFONUM;
wire    mem_BVALID;
reg    mem_BREADY;
reg   [0:0] phi_ln191_reg_370;
wire    ap_CS_fsm_state46;
reg    ap_block_state46_on_subcall_done;
reg    ap_predicate_op334_writeresp_state71;
reg    ap_block_state71;
reg    grp_kmeans_top_Pipeline_1_fu_381_ap_start_reg;
wire    ap_CS_fsm_state8;
reg   [106:0] ap_NS_fsm;
wire    ap_NS_fsm_state9;
wire    ap_CS_fsm_state9;
wire    ap_CS_fsm_state10;
reg    grp_kmeans_top_Pipeline_2_fu_390_ap_start_reg;
wire    ap_CS_fsm_state17;
wire    ap_NS_fsm_state18;
wire    ap_CS_fsm_state18;
wire    ap_CS_fsm_state19;
reg    grp_kmeans_top_Pipeline_3_fu_399_ap_start_reg;
wire    ap_CS_fsm_state26;
wire    ap_NS_fsm_state27;
wire    ap_CS_fsm_state27;
reg    grp_kmeans_top_Pipeline_4_fu_408_ap_start_reg;
wire    ap_CS_fsm_state35;
wire    ap_NS_fsm_state36;
wire    ap_CS_fsm_state36;
wire    ap_CS_fsm_state37;
reg    grp_kmeans_top_Pipeline_5_fu_417_ap_start_reg;
wire    ap_CS_fsm_state44;
wire    ap_NS_fsm_state45;
wire    ap_CS_fsm_state45;
reg    grp_kmeans_fu_426_ap_start_reg;
reg    grp_kmeans_top_Pipeline_6_fu_438_ap_start_reg;
wire    ap_NS_fsm_state50;
wire    ap_CS_fsm_state50;
wire    ap_CS_fsm_state51;
reg    grp_kmeans_top_Pipeline_7_fu_447_ap_start_reg;
wire    ap_NS_fsm_state58;
wire    ap_CS_fsm_state58;
wire    ap_CS_fsm_state59;
reg    grp_kmeans_top_Pipeline_8_fu_456_ap_start_reg;
wire    ap_NS_fsm_state65;
wire    ap_CS_fsm_state65;
wire    ap_CS_fsm_state66;
reg    grp_kmeans_top_Pipeline_9_fu_465_ap_start_reg;
wire    ap_NS_fsm_state73;
wire    ap_CS_fsm_state73;
wire    ap_CS_fsm_state74;
reg    grp_kmeans_top_Pipeline_10_fu_474_ap_start_reg;
wire    ap_NS_fsm_state80;
wire    ap_CS_fsm_state80;
wire    ap_CS_fsm_state81;
reg    grp_kmeans_top_Pipeline_11_fu_483_ap_start_reg;
wire    ap_NS_fsm_state87;
wire    ap_CS_fsm_state87;
wire    ap_CS_fsm_state88;
reg    grp_kmeans_top_Pipeline_12_fu_492_ap_start_reg;
wire    ap_NS_fsm_state94;
wire    ap_CS_fsm_state94;
wire    ap_CS_fsm_state95;
reg    grp_kmeans_top_Pipeline_13_fu_501_ap_start_reg;
wire    ap_NS_fsm_state101;
wire    ap_CS_fsm_state101;
wire    ap_CS_fsm_state102;
wire  signed [63:0] p_cast_cast_fu_655_p1;
wire  signed [63:0] p_cast2_cast_fu_666_p1;
wire  signed [63:0] p_cast4_cast_fu_677_p1;
wire  signed [63:0] p_cast1_cast_fu_693_p1;
wire  signed [63:0] p_cast3_cast_fu_704_p1;
wire  signed [63:0] p_cast9_cast_fu_816_p1;
wire  signed [63:0] p_cast11_cast_fu_871_p1;
wire  signed [63:0] p_cast13_cast_fu_881_p1;
wire  signed [63:0] p_cast5_cast_fu_910_p1;
wire  signed [63:0] p_cast8_cast_fu_921_p1;
wire  signed [63:0] p_cast6_cast_fu_932_p1;
wire  signed [63:0] p_cast7_cast_fu_947_p1;
wire  signed [63:0] p_cast12_cast_fu_958_p1;
reg    ap_block_state2_io;
reg    ap_predicate_op298_writeresp_state56;
reg    ap_block_state56;
reg    ap_predicate_op363_writeresp_state86;
reg    ap_block_state86;
reg    ap_predicate_op373_writereq_state86;
reg    ap_block_state86_io;
reg    ap_predicate_op380_writeresp_state93;
reg    ap_block_state93;
reg    ap_predicate_op390_writereq_state93;
reg    ap_block_state93_io;
reg    ap_predicate_op408_writeresp_state107;
reg    ap_block_state107;
reg   [31:0] n_assign_fu_158;
reg   [31:0] ap_sig_allocacmp_n_assign_load;
reg   [31:0] k_assign_fu_162;
reg   [2:0] control_assign_fu_166;
wire   [2:0] trunc_ln131_fu_620_p1;
reg   [63:0] max_iterations_assign_fu_170;
reg   [63:0] sub_iterations_assign_fu_174;
reg   [31:0] intermediate_writes_made_fu_198;
reg   [31:0] current_iteration_fu_202;
wire   [31:0] current_iteration_1_fu_895_p2;
wire  signed [31:0] sext_ln191_fu_734_p0;
wire  signed [63:0] sext_ln191_fu_734_p1;
wire   [27:0] trunc_ln194_1_fu_754_p1;
wire   [28:0] trunc_ln194_fu_747_p1;
wire   [28:0] shl_ln_fu_758_p3;
wire  signed [28:0] mul_ln194_fu_776_p0;
wire  signed [28:0] mul_ln194_fu_776_p1;
wire   [34:0] tmp_1_fu_790_p3;
wire   [63:0] p_cast14_fu_797_p1;
wire   [63:0] empty_50_fu_801_p2;
wire   [34:0] tmp_2_fu_830_p3;
wire   [63:0] p_cast15_fu_837_p1;
wire   [63:0] empty_53_fu_841_p2;
wire   [63:0] empty_56_fu_856_p2;
wire   [31:0] trunc_ln204_fu_891_p1;
reg    ap_block_state28_on_subcall_done;
reg    ap_ST_fsm_state1_blk;
reg    ap_ST_fsm_state2_blk;
wire    ap_ST_fsm_state3_blk;
wire    ap_ST_fsm_state4_blk;
wire    ap_ST_fsm_state5_blk;
wire    ap_ST_fsm_state6_blk;
wire    ap_ST_fsm_state7_blk;
wire    ap_ST_fsm_state8_blk;
wire    ap_ST_fsm_state9_blk;
reg    ap_ST_fsm_state10_blk;
reg    ap_ST_fsm_state11_blk;
wire    ap_ST_fsm_state12_blk;
wire    ap_ST_fsm_state13_blk;
wire    ap_ST_fsm_state14_blk;
wire    ap_ST_fsm_state15_blk;
wire    ap_ST_fsm_state16_blk;
wire    ap_ST_fsm_state17_blk;
wire    ap_ST_fsm_state18_blk;
reg    ap_ST_fsm_state19_blk;
reg    ap_ST_fsm_state20_blk;
wire    ap_ST_fsm_state21_blk;
wire    ap_ST_fsm_state22_blk;
wire    ap_ST_fsm_state23_blk;
wire    ap_ST_fsm_state24_blk;
wire    ap_ST_fsm_state25_blk;
wire    ap_ST_fsm_state26_blk;
wire    ap_ST_fsm_state27_blk;
reg    ap_ST_fsm_state28_blk;
reg    ap_ST_fsm_state29_blk;
wire    ap_ST_fsm_state30_blk;
wire    ap_ST_fsm_state31_blk;
wire    ap_ST_fsm_state32_blk;
wire    ap_ST_fsm_state33_blk;
wire    ap_ST_fsm_state34_blk;
wire    ap_ST_fsm_state35_blk;
wire    ap_ST_fsm_state36_blk;
reg    ap_ST_fsm_state37_blk;
reg    ap_ST_fsm_state38_blk;
wire    ap_ST_fsm_state39_blk;
wire    ap_ST_fsm_state40_blk;
wire    ap_ST_fsm_state41_blk;
wire    ap_ST_fsm_state42_blk;
wire    ap_ST_fsm_state43_blk;
wire    ap_ST_fsm_state44_blk;
wire    ap_ST_fsm_state45_blk;
reg    ap_ST_fsm_state46_blk;
wire    ap_ST_fsm_state47_blk;
reg    ap_ST_fsm_state48_blk;
reg    ap_ST_fsm_state49_blk;
wire    ap_ST_fsm_state50_blk;
reg    ap_ST_fsm_state51_blk;
wire    ap_ST_fsm_state52_blk;
wire    ap_ST_fsm_state53_blk;
wire    ap_ST_fsm_state54_blk;
wire    ap_ST_fsm_state55_blk;
reg    ap_ST_fsm_state56_blk;
reg    ap_ST_fsm_state57_blk;
wire    ap_ST_fsm_state58_blk;
reg    ap_ST_fsm_state59_blk;
wire    ap_ST_fsm_state60_blk;
wire    ap_ST_fsm_state61_blk;
wire    ap_ST_fsm_state62_blk;
wire    ap_ST_fsm_state63_blk;
reg    ap_ST_fsm_state64_blk;
wire    ap_ST_fsm_state65_blk;
reg    ap_ST_fsm_state66_blk;
wire    ap_ST_fsm_state67_blk;
wire    ap_ST_fsm_state68_blk;
wire    ap_ST_fsm_state69_blk;
wire    ap_ST_fsm_state70_blk;
reg    ap_ST_fsm_state71_blk;
reg    ap_ST_fsm_state72_blk;
wire    ap_ST_fsm_state73_blk;
reg    ap_ST_fsm_state74_blk;
wire    ap_ST_fsm_state75_blk;
wire    ap_ST_fsm_state76_blk;
wire    ap_ST_fsm_state77_blk;
wire    ap_ST_fsm_state78_blk;
reg    ap_ST_fsm_state79_blk;
wire    ap_ST_fsm_state80_blk;
reg    ap_ST_fsm_state81_blk;
wire    ap_ST_fsm_state82_blk;
wire    ap_ST_fsm_state83_blk;
wire    ap_ST_fsm_state84_blk;
wire    ap_ST_fsm_state85_blk;
reg    ap_ST_fsm_state86_blk;
wire    ap_ST_fsm_state87_blk;
reg    ap_ST_fsm_state88_blk;
wire    ap_ST_fsm_state89_blk;
wire    ap_ST_fsm_state90_blk;
wire    ap_ST_fsm_state91_blk;
wire    ap_ST_fsm_state92_blk;
reg    ap_ST_fsm_state93_blk;
wire    ap_ST_fsm_state94_blk;
reg    ap_ST_fsm_state95_blk;
wire    ap_ST_fsm_state96_blk;
wire    ap_ST_fsm_state97_blk;
wire    ap_ST_fsm_state98_blk;
wire    ap_ST_fsm_state99_blk;
reg    ap_ST_fsm_state100_blk;
wire    ap_ST_fsm_state101_blk;
reg    ap_ST_fsm_state102_blk;
wire    ap_ST_fsm_state103_blk;
wire    ap_ST_fsm_state104_blk;
wire    ap_ST_fsm_state105_blk;
wire    ap_ST_fsm_state106_blk;
reg    ap_ST_fsm_state107_blk;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_CS_fsm = 107'd1;
#0 grp_kmeans_top_Pipeline_1_fu_381_ap_start_reg = 1'b0;
#0 grp_kmeans_top_Pipeline_2_fu_390_ap_start_reg = 1'b0;
#0 grp_kmeans_top_Pipeline_3_fu_399_ap_start_reg = 1'b0;
#0 grp_kmeans_top_Pipeline_4_fu_408_ap_start_reg = 1'b0;
#0 grp_kmeans_top_Pipeline_5_fu_417_ap_start_reg = 1'b0;
#0 grp_kmeans_fu_426_ap_start_reg = 1'b0;
#0 grp_kmeans_top_Pipeline_6_fu_438_ap_start_reg = 1'b0;
#0 grp_kmeans_top_Pipeline_7_fu_447_ap_start_reg = 1'b0;
#0 grp_kmeans_top_Pipeline_8_fu_456_ap_start_reg = 1'b0;
#0 grp_kmeans_top_Pipeline_9_fu_465_ap_start_reg = 1'b0;
#0 grp_kmeans_top_Pipeline_10_fu_474_ap_start_reg = 1'b0;
#0 grp_kmeans_top_Pipeline_11_fu_483_ap_start_reg = 1'b0;
#0 grp_kmeans_top_Pipeline_12_fu_492_ap_start_reg = 1'b0;
#0 grp_kmeans_top_Pipeline_13_fu_501_ap_start_reg = 1'b0;
end

kmeans_top_node_x_coords_RAM_2P_URAM_1R1W #(
    .DataWidth( 64 ),
    .AddressRange( 8192 ),
    .AddressWidth( 13 ))
node_x_coords_U(
    .clk(ap_clk),
    .reset(ap_rst_n_inv),
    .address0(node_x_coords_address0),
    .ce0(node_x_coords_ce0),
    .q0(node_x_coords_q0),
    .address1(node_x_coords_address1),
    .ce1(node_x_coords_ce1),
    .we1(node_x_coords_we1),
    .d1(grp_kmeans_top_Pipeline_1_fu_381_node_x_coords_d1),
    .q1(node_x_coords_q1)
);

kmeans_top_node_x_coords_RAM_2P_URAM_1R1W #(
    .DataWidth( 64 ),
    .AddressRange( 8192 ),
    .AddressWidth( 13 ))
node_y_coords_U(
    .clk(ap_clk),
    .reset(ap_rst_n_inv),
    .address0(node_y_coords_address0),
    .ce0(node_y_coords_ce0),
    .q0(node_y_coords_q0),
    .address1(node_y_coords_address1),
    .ce1(node_y_coords_ce1),
    .we1(node_y_coords_we1),
    .d1(grp_kmeans_top_Pipeline_2_fu_390_node_y_coords_d1),
    .q1(node_y_coords_q1)
);

kmeans_top_node_cluster_assignments_RAM_2P_URAM_1R1W #(
    .DataWidth( 64 ),
    .AddressRange( 8192 ),
    .AddressWidth( 13 ))
node_cluster_assignments_U(
    .clk(ap_clk),
    .reset(ap_rst_n_inv),
    .address0(node_cluster_assignments_address0),
    .ce0(node_cluster_assignments_ce0),
    .q0(node_cluster_assignments_q0),
    .address1(node_cluster_assignments_address1),
    .ce1(node_cluster_assignments_ce1),
    .we1(node_cluster_assignments_we1),
    .d1(node_cluster_assignments_d1)
);

kmeans_top_centroid_x_coords_RAM_1WNR_AUTO_1R1W #(
    .DataWidth( 64 ),
    .AddressRange( 256 ),
    .AddressWidth( 8 ))
centroid_x_coords_U(
    .clk(ap_clk),
    .reset(ap_rst_n_inv),
    .address0(centroid_x_coords_address0),
    .ce0(centroid_x_coords_ce0),
    .we0(centroid_x_coords_we0),
    .d0(centroid_x_coords_d0),
    .q0(centroid_x_coords_q0),
    .address1(grp_kmeans_fu_426_centroid_x_coords_address1),
    .ce1(centroid_x_coords_ce1),
    .q1(centroid_x_coords_q1)
);

kmeans_top_centroid_x_coords_RAM_1WNR_AUTO_1R1W #(
    .DataWidth( 64 ),
    .AddressRange( 256 ),
    .AddressWidth( 8 ))
centroid_y_coords_U(
    .clk(ap_clk),
    .reset(ap_rst_n_inv),
    .address0(centroid_y_coords_address0),
    .ce0(centroid_y_coords_ce0),
    .we0(centroid_y_coords_we0),
    .d0(centroid_y_coords_d0),
    .q0(centroid_y_coords_q0),
    .address1(grp_kmeans_fu_426_centroid_y_coords_address1),
    .ce1(centroid_y_coords_ce1),
    .q1(centroid_y_coords_q1)
);

kmeans_top_kmeans_top_Pipeline_1 grp_kmeans_top_Pipeline_1_fu_381(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .ap_start(grp_kmeans_top_Pipeline_1_fu_381_ap_start),
    .ap_done(grp_kmeans_top_Pipeline_1_fu_381_ap_done),
    .ap_idle(grp_kmeans_top_Pipeline_1_fu_381_ap_idle),
    .ap_ready(grp_kmeans_top_Pipeline_1_fu_381_ap_ready),
    .m_axi_mem_AWVALID(grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_AWVALID),
    .m_axi_mem_AWREADY(1'b0),
    .m_axi_mem_AWADDR(grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_AWADDR),
    .m_axi_mem_AWID(grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_AWID),
    .m_axi_mem_AWLEN(grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_AWLEN),
    .m_axi_mem_AWSIZE(grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_AWSIZE),
    .m_axi_mem_AWBURST(grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_AWBURST),
    .m_axi_mem_AWLOCK(grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_AWLOCK),
    .m_axi_mem_AWCACHE(grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_AWCACHE),
    .m_axi_mem_AWPROT(grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_AWPROT),
    .m_axi_mem_AWQOS(grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_AWQOS),
    .m_axi_mem_AWREGION(grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_AWREGION),
    .m_axi_mem_AWUSER(grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_AWUSER),
    .m_axi_mem_WVALID(grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_WVALID),
    .m_axi_mem_WREADY(1'b0),
    .m_axi_mem_WDATA(grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_WDATA),
    .m_axi_mem_WSTRB(grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_WSTRB),
    .m_axi_mem_WLAST(grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_WLAST),
    .m_axi_mem_WID(grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_WID),
    .m_axi_mem_WUSER(grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_WUSER),
    .m_axi_mem_ARVALID(grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_ARVALID),
    .m_axi_mem_ARREADY(mem_ARREADY),
    .m_axi_mem_ARADDR(grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_ARADDR),
    .m_axi_mem_ARID(grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_ARID),
    .m_axi_mem_ARLEN(grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_ARLEN),
    .m_axi_mem_ARSIZE(grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_ARSIZE),
    .m_axi_mem_ARBURST(grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_ARBURST),
    .m_axi_mem_ARLOCK(grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_ARLOCK),
    .m_axi_mem_ARCACHE(grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_ARCACHE),
    .m_axi_mem_ARPROT(grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_ARPROT),
    .m_axi_mem_ARQOS(grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_ARQOS),
    .m_axi_mem_ARREGION(grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_ARREGION),
    .m_axi_mem_ARUSER(grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_ARUSER),
    .m_axi_mem_RVALID(mem_RVALID),
    .m_axi_mem_RREADY(grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_RREADY),
    .m_axi_mem_RDATA(mem_RDATA),
    .m_axi_mem_RLAST(1'b0),
    .m_axi_mem_RID(1'd0),
    .m_axi_mem_RFIFONUM(mem_RFIFONUM),
    .m_axi_mem_RUSER(1'd0),
    .m_axi_mem_RRESP(2'd0),
    .m_axi_mem_BVALID(1'b0),
    .m_axi_mem_BREADY(grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_BREADY),
    .m_axi_mem_BRESP(2'd0),
    .m_axi_mem_BID(1'd0),
    .m_axi_mem_BUSER(1'd0),
    .p_cast_cast(reg_590),
    .node_x_coords_address1(grp_kmeans_top_Pipeline_1_fu_381_node_x_coords_address1),
    .node_x_coords_ce1(grp_kmeans_top_Pipeline_1_fu_381_node_x_coords_ce1),
    .node_x_coords_we1(grp_kmeans_top_Pipeline_1_fu_381_node_x_coords_we1),
    .node_x_coords_d1(grp_kmeans_top_Pipeline_1_fu_381_node_x_coords_d1),
    .sext_ln182(n_assign_load_reg_1041)
);

kmeans_top_kmeans_top_Pipeline_2 grp_kmeans_top_Pipeline_2_fu_390(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .ap_start(grp_kmeans_top_Pipeline_2_fu_390_ap_start),
    .ap_done(grp_kmeans_top_Pipeline_2_fu_390_ap_done),
    .ap_idle(grp_kmeans_top_Pipeline_2_fu_390_ap_idle),
    .ap_ready(grp_kmeans_top_Pipeline_2_fu_390_ap_ready),
    .m_axi_mem_AWVALID(grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_AWVALID),
    .m_axi_mem_AWREADY(1'b0),
    .m_axi_mem_AWADDR(grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_AWADDR),
    .m_axi_mem_AWID(grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_AWID),
    .m_axi_mem_AWLEN(grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_AWLEN),
    .m_axi_mem_AWSIZE(grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_AWSIZE),
    .m_axi_mem_AWBURST(grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_AWBURST),
    .m_axi_mem_AWLOCK(grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_AWLOCK),
    .m_axi_mem_AWCACHE(grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_AWCACHE),
    .m_axi_mem_AWPROT(grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_AWPROT),
    .m_axi_mem_AWQOS(grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_AWQOS),
    .m_axi_mem_AWREGION(grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_AWREGION),
    .m_axi_mem_AWUSER(grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_AWUSER),
    .m_axi_mem_WVALID(grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_WVALID),
    .m_axi_mem_WREADY(1'b0),
    .m_axi_mem_WDATA(grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_WDATA),
    .m_axi_mem_WSTRB(grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_WSTRB),
    .m_axi_mem_WLAST(grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_WLAST),
    .m_axi_mem_WID(grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_WID),
    .m_axi_mem_WUSER(grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_WUSER),
    .m_axi_mem_ARVALID(grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_ARVALID),
    .m_axi_mem_ARREADY(mem_ARREADY),
    .m_axi_mem_ARADDR(grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_ARADDR),
    .m_axi_mem_ARID(grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_ARID),
    .m_axi_mem_ARLEN(grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_ARLEN),
    .m_axi_mem_ARSIZE(grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_ARSIZE),
    .m_axi_mem_ARBURST(grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_ARBURST),
    .m_axi_mem_ARLOCK(grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_ARLOCK),
    .m_axi_mem_ARCACHE(grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_ARCACHE),
    .m_axi_mem_ARPROT(grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_ARPROT),
    .m_axi_mem_ARQOS(grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_ARQOS),
    .m_axi_mem_ARREGION(grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_ARREGION),
    .m_axi_mem_ARUSER(grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_ARUSER),
    .m_axi_mem_RVALID(mem_RVALID),
    .m_axi_mem_RREADY(grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_RREADY),
    .m_axi_mem_RDATA(mem_RDATA),
    .m_axi_mem_RLAST(1'b0),
    .m_axi_mem_RID(1'd0),
    .m_axi_mem_RFIFONUM(mem_RFIFONUM),
    .m_axi_mem_RUSER(1'd0),
    .m_axi_mem_RRESP(2'd0),
    .m_axi_mem_BVALID(1'b0),
    .m_axi_mem_BREADY(grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_BREADY),
    .m_axi_mem_BRESP(2'd0),
    .m_axi_mem_BID(1'd0),
    .m_axi_mem_BUSER(1'd0),
    .p_cast2_cast(reg_596),
    .node_y_coords_address1(grp_kmeans_top_Pipeline_2_fu_390_node_y_coords_address1),
    .node_y_coords_ce1(grp_kmeans_top_Pipeline_2_fu_390_node_y_coords_ce1),
    .node_y_coords_we1(grp_kmeans_top_Pipeline_2_fu_390_node_y_coords_we1),
    .node_y_coords_d1(grp_kmeans_top_Pipeline_2_fu_390_node_y_coords_d1),
    .sext_ln182(n_assign_load_reg_1041)
);

kmeans_top_kmeans_top_Pipeline_3 grp_kmeans_top_Pipeline_3_fu_399(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .ap_start(grp_kmeans_top_Pipeline_3_fu_399_ap_start),
    .ap_done(grp_kmeans_top_Pipeline_3_fu_399_ap_done),
    .ap_idle(grp_kmeans_top_Pipeline_3_fu_399_ap_idle),
    .ap_ready(grp_kmeans_top_Pipeline_3_fu_399_ap_ready),
    .m_axi_mem_AWVALID(grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_AWVALID),
    .m_axi_mem_AWREADY(1'b0),
    .m_axi_mem_AWADDR(grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_AWADDR),
    .m_axi_mem_AWID(grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_AWID),
    .m_axi_mem_AWLEN(grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_AWLEN),
    .m_axi_mem_AWSIZE(grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_AWSIZE),
    .m_axi_mem_AWBURST(grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_AWBURST),
    .m_axi_mem_AWLOCK(grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_AWLOCK),
    .m_axi_mem_AWCACHE(grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_AWCACHE),
    .m_axi_mem_AWPROT(grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_AWPROT),
    .m_axi_mem_AWQOS(grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_AWQOS),
    .m_axi_mem_AWREGION(grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_AWREGION),
    .m_axi_mem_AWUSER(grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_AWUSER),
    .m_axi_mem_WVALID(grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_WVALID),
    .m_axi_mem_WREADY(1'b0),
    .m_axi_mem_WDATA(grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_WDATA),
    .m_axi_mem_WSTRB(grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_WSTRB),
    .m_axi_mem_WLAST(grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_WLAST),
    .m_axi_mem_WID(grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_WID),
    .m_axi_mem_WUSER(grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_WUSER),
    .m_axi_mem_ARVALID(grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_ARVALID),
    .m_axi_mem_ARREADY(mem_ARREADY),
    .m_axi_mem_ARADDR(grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_ARADDR),
    .m_axi_mem_ARID(grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_ARID),
    .m_axi_mem_ARLEN(grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_ARLEN),
    .m_axi_mem_ARSIZE(grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_ARSIZE),
    .m_axi_mem_ARBURST(grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_ARBURST),
    .m_axi_mem_ARLOCK(grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_ARLOCK),
    .m_axi_mem_ARCACHE(grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_ARCACHE),
    .m_axi_mem_ARPROT(grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_ARPROT),
    .m_axi_mem_ARQOS(grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_ARQOS),
    .m_axi_mem_ARREGION(grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_ARREGION),
    .m_axi_mem_ARUSER(grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_ARUSER),
    .m_axi_mem_RVALID(mem_RVALID),
    .m_axi_mem_RREADY(grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_RREADY),
    .m_axi_mem_RDATA(mem_RDATA),
    .m_axi_mem_RLAST(1'b0),
    .m_axi_mem_RID(1'd0),
    .m_axi_mem_RFIFONUM(mem_RFIFONUM),
    .m_axi_mem_RUSER(1'd0),
    .m_axi_mem_RRESP(2'd0),
    .m_axi_mem_BVALID(1'b0),
    .m_axi_mem_BREADY(grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_BREADY),
    .m_axi_mem_BRESP(2'd0),
    .m_axi_mem_BID(1'd0),
    .m_axi_mem_BUSER(1'd0),
    .p_cast4_cast(reg_602),
    .node_cluster_assignments_address1(grp_kmeans_top_Pipeline_3_fu_399_node_cluster_assignments_address1),
    .node_cluster_assignments_ce1(grp_kmeans_top_Pipeline_3_fu_399_node_cluster_assignments_ce1),
    .node_cluster_assignments_we1(grp_kmeans_top_Pipeline_3_fu_399_node_cluster_assignments_we1),
    .node_cluster_assignments_d1(grp_kmeans_top_Pipeline_3_fu_399_node_cluster_assignments_d1),
    .sext_ln182(n_assign_load_reg_1041)
);

kmeans_top_kmeans_top_Pipeline_4 grp_kmeans_top_Pipeline_4_fu_408(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .ap_start(grp_kmeans_top_Pipeline_4_fu_408_ap_start),
    .ap_done(grp_kmeans_top_Pipeline_4_fu_408_ap_done),
    .ap_idle(grp_kmeans_top_Pipeline_4_fu_408_ap_idle),
    .ap_ready(grp_kmeans_top_Pipeline_4_fu_408_ap_ready),
    .m_axi_mem_AWVALID(grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_AWVALID),
    .m_axi_mem_AWREADY(1'b0),
    .m_axi_mem_AWADDR(grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_AWADDR),
    .m_axi_mem_AWID(grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_AWID),
    .m_axi_mem_AWLEN(grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_AWLEN),
    .m_axi_mem_AWSIZE(grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_AWSIZE),
    .m_axi_mem_AWBURST(grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_AWBURST),
    .m_axi_mem_AWLOCK(grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_AWLOCK),
    .m_axi_mem_AWCACHE(grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_AWCACHE),
    .m_axi_mem_AWPROT(grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_AWPROT),
    .m_axi_mem_AWQOS(grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_AWQOS),
    .m_axi_mem_AWREGION(grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_AWREGION),
    .m_axi_mem_AWUSER(grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_AWUSER),
    .m_axi_mem_WVALID(grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_WVALID),
    .m_axi_mem_WREADY(1'b0),
    .m_axi_mem_WDATA(grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_WDATA),
    .m_axi_mem_WSTRB(grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_WSTRB),
    .m_axi_mem_WLAST(grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_WLAST),
    .m_axi_mem_WID(grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_WID),
    .m_axi_mem_WUSER(grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_WUSER),
    .m_axi_mem_ARVALID(grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_ARVALID),
    .m_axi_mem_ARREADY(mem_ARREADY),
    .m_axi_mem_ARADDR(grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_ARADDR),
    .m_axi_mem_ARID(grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_ARID),
    .m_axi_mem_ARLEN(grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_ARLEN),
    .m_axi_mem_ARSIZE(grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_ARSIZE),
    .m_axi_mem_ARBURST(grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_ARBURST),
    .m_axi_mem_ARLOCK(grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_ARLOCK),
    .m_axi_mem_ARCACHE(grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_ARCACHE),
    .m_axi_mem_ARPROT(grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_ARPROT),
    .m_axi_mem_ARQOS(grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_ARQOS),
    .m_axi_mem_ARREGION(grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_ARREGION),
    .m_axi_mem_ARUSER(grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_ARUSER),
    .m_axi_mem_RVALID(mem_RVALID),
    .m_axi_mem_RREADY(grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_RREADY),
    .m_axi_mem_RDATA(mem_RDATA),
    .m_axi_mem_RLAST(1'b0),
    .m_axi_mem_RID(1'd0),
    .m_axi_mem_RFIFONUM(mem_RFIFONUM),
    .m_axi_mem_RUSER(1'd0),
    .m_axi_mem_RRESP(2'd0),
    .m_axi_mem_BVALID(1'b0),
    .m_axi_mem_BREADY(grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_BREADY),
    .m_axi_mem_BRESP(2'd0),
    .m_axi_mem_BID(1'd0),
    .m_axi_mem_BUSER(1'd0),
    .p_cast1_cast(reg_608),
    .centroid_x_coords_address0(grp_kmeans_top_Pipeline_4_fu_408_centroid_x_coords_address0),
    .centroid_x_coords_ce0(grp_kmeans_top_Pipeline_4_fu_408_centroid_x_coords_ce0),
    .centroid_x_coords_we0(grp_kmeans_top_Pipeline_4_fu_408_centroid_x_coords_we0),
    .centroid_x_coords_d0(grp_kmeans_top_Pipeline_4_fu_408_centroid_x_coords_d0),
    .sext_ln185(k_assign_load_reg_1063)
);

kmeans_top_kmeans_top_Pipeline_5 grp_kmeans_top_Pipeline_5_fu_417(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .ap_start(grp_kmeans_top_Pipeline_5_fu_417_ap_start),
    .ap_done(grp_kmeans_top_Pipeline_5_fu_417_ap_done),
    .ap_idle(grp_kmeans_top_Pipeline_5_fu_417_ap_idle),
    .ap_ready(grp_kmeans_top_Pipeline_5_fu_417_ap_ready),
    .m_axi_mem_AWVALID(grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_AWVALID),
    .m_axi_mem_AWREADY(1'b0),
    .m_axi_mem_AWADDR(grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_AWADDR),
    .m_axi_mem_AWID(grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_AWID),
    .m_axi_mem_AWLEN(grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_AWLEN),
    .m_axi_mem_AWSIZE(grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_AWSIZE),
    .m_axi_mem_AWBURST(grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_AWBURST),
    .m_axi_mem_AWLOCK(grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_AWLOCK),
    .m_axi_mem_AWCACHE(grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_AWCACHE),
    .m_axi_mem_AWPROT(grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_AWPROT),
    .m_axi_mem_AWQOS(grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_AWQOS),
    .m_axi_mem_AWREGION(grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_AWREGION),
    .m_axi_mem_AWUSER(grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_AWUSER),
    .m_axi_mem_WVALID(grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_WVALID),
    .m_axi_mem_WREADY(1'b0),
    .m_axi_mem_WDATA(grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_WDATA),
    .m_axi_mem_WSTRB(grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_WSTRB),
    .m_axi_mem_WLAST(grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_WLAST),
    .m_axi_mem_WID(grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_WID),
    .m_axi_mem_WUSER(grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_WUSER),
    .m_axi_mem_ARVALID(grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_ARVALID),
    .m_axi_mem_ARREADY(mem_ARREADY),
    .m_axi_mem_ARADDR(grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_ARADDR),
    .m_axi_mem_ARID(grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_ARID),
    .m_axi_mem_ARLEN(grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_ARLEN),
    .m_axi_mem_ARSIZE(grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_ARSIZE),
    .m_axi_mem_ARBURST(grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_ARBURST),
    .m_axi_mem_ARLOCK(grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_ARLOCK),
    .m_axi_mem_ARCACHE(grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_ARCACHE),
    .m_axi_mem_ARPROT(grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_ARPROT),
    .m_axi_mem_ARQOS(grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_ARQOS),
    .m_axi_mem_ARREGION(grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_ARREGION),
    .m_axi_mem_ARUSER(grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_ARUSER),
    .m_axi_mem_RVALID(mem_RVALID),
    .m_axi_mem_RREADY(grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_RREADY),
    .m_axi_mem_RDATA(mem_RDATA),
    .m_axi_mem_RLAST(1'b0),
    .m_axi_mem_RID(1'd0),
    .m_axi_mem_RFIFONUM(mem_RFIFONUM),
    .m_axi_mem_RUSER(1'd0),
    .m_axi_mem_RRESP(2'd0),
    .m_axi_mem_BVALID(1'b0),
    .m_axi_mem_BREADY(grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_BREADY),
    .m_axi_mem_BRESP(2'd0),
    .m_axi_mem_BID(1'd0),
    .m_axi_mem_BUSER(1'd0),
    .p_cast3_cast(reg_614),
    .centroid_y_coords_address0(grp_kmeans_top_Pipeline_5_fu_417_centroid_y_coords_address0),
    .centroid_y_coords_ce0(grp_kmeans_top_Pipeline_5_fu_417_centroid_y_coords_ce0),
    .centroid_y_coords_we0(grp_kmeans_top_Pipeline_5_fu_417_centroid_y_coords_we0),
    .centroid_y_coords_d0(grp_kmeans_top_Pipeline_5_fu_417_centroid_y_coords_d0),
    .sext_ln185(k_assign_load_reg_1063)
);

kmeans_top_kmeans grp_kmeans_fu_426(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .ap_start(grp_kmeans_fu_426_ap_start),
    .ap_done(grp_kmeans_fu_426_ap_done),
    .ap_idle(grp_kmeans_fu_426_ap_idle),
    .ap_ready(grp_kmeans_fu_426_ap_ready),
    .node_x_coords_address0(grp_kmeans_fu_426_node_x_coords_address0),
    .node_x_coords_ce0(grp_kmeans_fu_426_node_x_coords_ce0),
    .node_x_coords_q0(node_x_coords_q0),
    .node_x_coords_address1(grp_kmeans_fu_426_node_x_coords_address1),
    .node_x_coords_ce1(grp_kmeans_fu_426_node_x_coords_ce1),
    .node_x_coords_q1(node_x_coords_q1),
    .node_y_coords_address0(grp_kmeans_fu_426_node_y_coords_address0),
    .node_y_coords_ce0(grp_kmeans_fu_426_node_y_coords_ce0),
    .node_y_coords_q0(node_y_coords_q0),
    .node_y_coords_address1(grp_kmeans_fu_426_node_y_coords_address1),
    .node_y_coords_ce1(grp_kmeans_fu_426_node_y_coords_ce1),
    .node_y_coords_q1(node_y_coords_q1),
    .node_cluster_assignments_address1(grp_kmeans_fu_426_node_cluster_assignments_address1),
    .node_cluster_assignments_ce1(grp_kmeans_fu_426_node_cluster_assignments_ce1),
    .node_cluster_assignments_we1(grp_kmeans_fu_426_node_cluster_assignments_we1),
    .node_cluster_assignments_d1(grp_kmeans_fu_426_node_cluster_assignments_d1),
    .centroid_x_coords_address0(grp_kmeans_fu_426_centroid_x_coords_address0),
    .centroid_x_coords_ce0(grp_kmeans_fu_426_centroid_x_coords_ce0),
    .centroid_x_coords_we0(grp_kmeans_fu_426_centroid_x_coords_we0),
    .centroid_x_coords_d0(grp_kmeans_fu_426_centroid_x_coords_d0),
    .centroid_x_coords_q0(centroid_x_coords_q0),
    .centroid_x_coords_address1(grp_kmeans_fu_426_centroid_x_coords_address1),
    .centroid_x_coords_ce1(grp_kmeans_fu_426_centroid_x_coords_ce1),
    .centroid_x_coords_q1(centroid_x_coords_q1),
    .centroid_y_coords_address0(grp_kmeans_fu_426_centroid_y_coords_address0),
    .centroid_y_coords_ce0(grp_kmeans_fu_426_centroid_y_coords_ce0),
    .centroid_y_coords_we0(grp_kmeans_fu_426_centroid_y_coords_we0),
    .centroid_y_coords_d0(grp_kmeans_fu_426_centroid_y_coords_d0),
    .centroid_y_coords_q0(centroid_y_coords_q0),
    .centroid_y_coords_address1(grp_kmeans_fu_426_centroid_y_coords_address1),
    .centroid_y_coords_ce1(grp_kmeans_fu_426_centroid_y_coords_ce1),
    .centroid_y_coords_q1(centroid_y_coords_q1),
    .max_iterations(sub_iterations_assign_load_reg_1131),
    .n(n_assign_load_1_reg_1136),
    .k(k_assign_load_1_reg_1141),
    .ap_return(grp_kmeans_fu_426_ap_return)
);

kmeans_top_kmeans_top_Pipeline_6 grp_kmeans_top_Pipeline_6_fu_438(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .ap_start(grp_kmeans_top_Pipeline_6_fu_438_ap_start),
    .ap_done(grp_kmeans_top_Pipeline_6_fu_438_ap_done),
    .ap_idle(grp_kmeans_top_Pipeline_6_fu_438_ap_idle),
    .ap_ready(grp_kmeans_top_Pipeline_6_fu_438_ap_ready),
    .m_axi_mem_AWVALID(grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_AWVALID),
    .m_axi_mem_AWREADY(mem_AWREADY),
    .m_axi_mem_AWADDR(grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_AWADDR),
    .m_axi_mem_AWID(grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_AWID),
    .m_axi_mem_AWLEN(grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_AWLEN),
    .m_axi_mem_AWSIZE(grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_AWSIZE),
    .m_axi_mem_AWBURST(grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_AWBURST),
    .m_axi_mem_AWLOCK(grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_AWLOCK),
    .m_axi_mem_AWCACHE(grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_AWCACHE),
    .m_axi_mem_AWPROT(grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_AWPROT),
    .m_axi_mem_AWQOS(grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_AWQOS),
    .m_axi_mem_AWREGION(grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_AWREGION),
    .m_axi_mem_AWUSER(grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_AWUSER),
    .m_axi_mem_WVALID(grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_WVALID),
    .m_axi_mem_WREADY(mem_WREADY),
    .m_axi_mem_WDATA(grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_WDATA),
    .m_axi_mem_WSTRB(grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_WSTRB),
    .m_axi_mem_WLAST(grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_WLAST),
    .m_axi_mem_WID(grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_WID),
    .m_axi_mem_WUSER(grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_WUSER),
    .m_axi_mem_ARVALID(grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_ARVALID),
    .m_axi_mem_ARREADY(1'b0),
    .m_axi_mem_ARADDR(grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_ARADDR),
    .m_axi_mem_ARID(grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_ARID),
    .m_axi_mem_ARLEN(grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_ARLEN),
    .m_axi_mem_ARSIZE(grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_ARSIZE),
    .m_axi_mem_ARBURST(grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_ARBURST),
    .m_axi_mem_ARLOCK(grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_ARLOCK),
    .m_axi_mem_ARCACHE(grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_ARCACHE),
    .m_axi_mem_ARPROT(grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_ARPROT),
    .m_axi_mem_ARQOS(grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_ARQOS),
    .m_axi_mem_ARREGION(grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_ARREGION),
    .m_axi_mem_ARUSER(grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_ARUSER),
    .m_axi_mem_RVALID(1'b0),
    .m_axi_mem_RREADY(grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_RREADY),
    .m_axi_mem_RDATA(64'd0),
    .m_axi_mem_RLAST(1'b0),
    .m_axi_mem_RID(1'd0),
    .m_axi_mem_RFIFONUM(9'd0),
    .m_axi_mem_RUSER(1'd0),
    .m_axi_mem_RRESP(2'd0),
    .m_axi_mem_BVALID(mem_BVALID),
    .m_axi_mem_BREADY(grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_BREADY),
    .m_axi_mem_BRESP(2'd0),
    .m_axi_mem_BID(1'd0),
    .m_axi_mem_BUSER(1'd0),
    .p_cast9_cast(p_cast9_reg_1169),
    .node_cluster_assignments_address0(grp_kmeans_top_Pipeline_6_fu_438_node_cluster_assignments_address0),
    .node_cluster_assignments_ce0(grp_kmeans_top_Pipeline_6_fu_438_node_cluster_assignments_ce0),
    .node_cluster_assignments_q0(node_cluster_assignments_q0),
    .sext_ln182(n_assign_load_reg_1041)
);

kmeans_top_kmeans_top_Pipeline_7 grp_kmeans_top_Pipeline_7_fu_447(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .ap_start(grp_kmeans_top_Pipeline_7_fu_447_ap_start),
    .ap_done(grp_kmeans_top_Pipeline_7_fu_447_ap_done),
    .ap_idle(grp_kmeans_top_Pipeline_7_fu_447_ap_idle),
    .ap_ready(grp_kmeans_top_Pipeline_7_fu_447_ap_ready),
    .m_axi_mem_AWVALID(grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_AWVALID),
    .m_axi_mem_AWREADY(mem_AWREADY),
    .m_axi_mem_AWADDR(grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_AWADDR),
    .m_axi_mem_AWID(grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_AWID),
    .m_axi_mem_AWLEN(grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_AWLEN),
    .m_axi_mem_AWSIZE(grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_AWSIZE),
    .m_axi_mem_AWBURST(grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_AWBURST),
    .m_axi_mem_AWLOCK(grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_AWLOCK),
    .m_axi_mem_AWCACHE(grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_AWCACHE),
    .m_axi_mem_AWPROT(grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_AWPROT),
    .m_axi_mem_AWQOS(grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_AWQOS),
    .m_axi_mem_AWREGION(grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_AWREGION),
    .m_axi_mem_AWUSER(grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_AWUSER),
    .m_axi_mem_WVALID(grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_WVALID),
    .m_axi_mem_WREADY(mem_WREADY),
    .m_axi_mem_WDATA(grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_WDATA),
    .m_axi_mem_WSTRB(grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_WSTRB),
    .m_axi_mem_WLAST(grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_WLAST),
    .m_axi_mem_WID(grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_WID),
    .m_axi_mem_WUSER(grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_WUSER),
    .m_axi_mem_ARVALID(grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_ARVALID),
    .m_axi_mem_ARREADY(1'b0),
    .m_axi_mem_ARADDR(grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_ARADDR),
    .m_axi_mem_ARID(grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_ARID),
    .m_axi_mem_ARLEN(grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_ARLEN),
    .m_axi_mem_ARSIZE(grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_ARSIZE),
    .m_axi_mem_ARBURST(grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_ARBURST),
    .m_axi_mem_ARLOCK(grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_ARLOCK),
    .m_axi_mem_ARCACHE(grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_ARCACHE),
    .m_axi_mem_ARPROT(grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_ARPROT),
    .m_axi_mem_ARQOS(grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_ARQOS),
    .m_axi_mem_ARREGION(grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_ARREGION),
    .m_axi_mem_ARUSER(grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_ARUSER),
    .m_axi_mem_RVALID(1'b0),
    .m_axi_mem_RREADY(grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_RREADY),
    .m_axi_mem_RDATA(64'd0),
    .m_axi_mem_RLAST(1'b0),
    .m_axi_mem_RID(1'd0),
    .m_axi_mem_RFIFONUM(9'd0),
    .m_axi_mem_RUSER(1'd0),
    .m_axi_mem_RRESP(2'd0),
    .m_axi_mem_BVALID(mem_BVALID),
    .m_axi_mem_BREADY(grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_BREADY),
    .m_axi_mem_BRESP(2'd0),
    .m_axi_mem_BID(1'd0),
    .m_axi_mem_BUSER(1'd0),
    .p_cast11_cast(p_cast10_reg_1188),
    .centroid_x_coords_address0(grp_kmeans_top_Pipeline_7_fu_447_centroid_x_coords_address0),
    .centroid_x_coords_ce0(grp_kmeans_top_Pipeline_7_fu_447_centroid_x_coords_ce0),
    .centroid_x_coords_q0(centroid_x_coords_q0),
    .sext_ln185(k_assign_load_reg_1063)
);

kmeans_top_kmeans_top_Pipeline_8 grp_kmeans_top_Pipeline_8_fu_456(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .ap_start(grp_kmeans_top_Pipeline_8_fu_456_ap_start),
    .ap_done(grp_kmeans_top_Pipeline_8_fu_456_ap_done),
    .ap_idle(grp_kmeans_top_Pipeline_8_fu_456_ap_idle),
    .ap_ready(grp_kmeans_top_Pipeline_8_fu_456_ap_ready),
    .m_axi_mem_AWVALID(grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_AWVALID),
    .m_axi_mem_AWREADY(mem_AWREADY),
    .m_axi_mem_AWADDR(grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_AWADDR),
    .m_axi_mem_AWID(grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_AWID),
    .m_axi_mem_AWLEN(grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_AWLEN),
    .m_axi_mem_AWSIZE(grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_AWSIZE),
    .m_axi_mem_AWBURST(grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_AWBURST),
    .m_axi_mem_AWLOCK(grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_AWLOCK),
    .m_axi_mem_AWCACHE(grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_AWCACHE),
    .m_axi_mem_AWPROT(grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_AWPROT),
    .m_axi_mem_AWQOS(grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_AWQOS),
    .m_axi_mem_AWREGION(grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_AWREGION),
    .m_axi_mem_AWUSER(grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_AWUSER),
    .m_axi_mem_WVALID(grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_WVALID),
    .m_axi_mem_WREADY(mem_WREADY),
    .m_axi_mem_WDATA(grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_WDATA),
    .m_axi_mem_WSTRB(grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_WSTRB),
    .m_axi_mem_WLAST(grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_WLAST),
    .m_axi_mem_WID(grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_WID),
    .m_axi_mem_WUSER(grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_WUSER),
    .m_axi_mem_ARVALID(grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_ARVALID),
    .m_axi_mem_ARREADY(1'b0),
    .m_axi_mem_ARADDR(grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_ARADDR),
    .m_axi_mem_ARID(grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_ARID),
    .m_axi_mem_ARLEN(grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_ARLEN),
    .m_axi_mem_ARSIZE(grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_ARSIZE),
    .m_axi_mem_ARBURST(grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_ARBURST),
    .m_axi_mem_ARLOCK(grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_ARLOCK),
    .m_axi_mem_ARCACHE(grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_ARCACHE),
    .m_axi_mem_ARPROT(grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_ARPROT),
    .m_axi_mem_ARQOS(grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_ARQOS),
    .m_axi_mem_ARREGION(grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_ARREGION),
    .m_axi_mem_ARUSER(grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_ARUSER),
    .m_axi_mem_RVALID(1'b0),
    .m_axi_mem_RREADY(grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_RREADY),
    .m_axi_mem_RDATA(64'd0),
    .m_axi_mem_RLAST(1'b0),
    .m_axi_mem_RID(1'd0),
    .m_axi_mem_RFIFONUM(9'd0),
    .m_axi_mem_RUSER(1'd0),
    .m_axi_mem_RRESP(2'd0),
    .m_axi_mem_BVALID(mem_BVALID),
    .m_axi_mem_BREADY(grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_BREADY),
    .m_axi_mem_BRESP(2'd0),
    .m_axi_mem_BID(1'd0),
    .m_axi_mem_BUSER(1'd0),
    .p_cast13_cast(p_cast11_reg_1194),
    .centroid_y_coords_address0(grp_kmeans_top_Pipeline_8_fu_456_centroid_y_coords_address0),
    .centroid_y_coords_ce0(grp_kmeans_top_Pipeline_8_fu_456_centroid_y_coords_ce0),
    .centroid_y_coords_q0(centroid_y_coords_q0),
    .sext_ln185(k_assign_load_reg_1063)
);

kmeans_top_kmeans_top_Pipeline_9 grp_kmeans_top_Pipeline_9_fu_465(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .ap_start(grp_kmeans_top_Pipeline_9_fu_465_ap_start),
    .ap_done(grp_kmeans_top_Pipeline_9_fu_465_ap_done),
    .ap_idle(grp_kmeans_top_Pipeline_9_fu_465_ap_idle),
    .ap_ready(grp_kmeans_top_Pipeline_9_fu_465_ap_ready),
    .m_axi_mem_AWVALID(grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_AWVALID),
    .m_axi_mem_AWREADY(mem_AWREADY),
    .m_axi_mem_AWADDR(grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_AWADDR),
    .m_axi_mem_AWID(grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_AWID),
    .m_axi_mem_AWLEN(grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_AWLEN),
    .m_axi_mem_AWSIZE(grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_AWSIZE),
    .m_axi_mem_AWBURST(grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_AWBURST),
    .m_axi_mem_AWLOCK(grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_AWLOCK),
    .m_axi_mem_AWCACHE(grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_AWCACHE),
    .m_axi_mem_AWPROT(grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_AWPROT),
    .m_axi_mem_AWQOS(grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_AWQOS),
    .m_axi_mem_AWREGION(grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_AWREGION),
    .m_axi_mem_AWUSER(grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_AWUSER),
    .m_axi_mem_WVALID(grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_WVALID),
    .m_axi_mem_WREADY(mem_WREADY),
    .m_axi_mem_WDATA(grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_WDATA),
    .m_axi_mem_WSTRB(grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_WSTRB),
    .m_axi_mem_WLAST(grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_WLAST),
    .m_axi_mem_WID(grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_WID),
    .m_axi_mem_WUSER(grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_WUSER),
    .m_axi_mem_ARVALID(grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_ARVALID),
    .m_axi_mem_ARREADY(1'b0),
    .m_axi_mem_ARADDR(grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_ARADDR),
    .m_axi_mem_ARID(grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_ARID),
    .m_axi_mem_ARLEN(grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_ARLEN),
    .m_axi_mem_ARSIZE(grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_ARSIZE),
    .m_axi_mem_ARBURST(grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_ARBURST),
    .m_axi_mem_ARLOCK(grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_ARLOCK),
    .m_axi_mem_ARCACHE(grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_ARCACHE),
    .m_axi_mem_ARPROT(grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_ARPROT),
    .m_axi_mem_ARQOS(grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_ARQOS),
    .m_axi_mem_ARREGION(grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_ARREGION),
    .m_axi_mem_ARUSER(grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_ARUSER),
    .m_axi_mem_RVALID(1'b0),
    .m_axi_mem_RREADY(grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_RREADY),
    .m_axi_mem_RDATA(64'd0),
    .m_axi_mem_RLAST(1'b0),
    .m_axi_mem_RID(1'd0),
    .m_axi_mem_RFIFONUM(9'd0),
    .m_axi_mem_RUSER(1'd0),
    .m_axi_mem_RRESP(2'd0),
    .m_axi_mem_BVALID(mem_BVALID),
    .m_axi_mem_BREADY(grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_BREADY),
    .m_axi_mem_BRESP(2'd0),
    .m_axi_mem_BID(1'd0),
    .m_axi_mem_BUSER(1'd0),
    .p_cast5_cast(reg_590),
    .node_x_coords_address0(grp_kmeans_top_Pipeline_9_fu_465_node_x_coords_address0),
    .node_x_coords_ce0(grp_kmeans_top_Pipeline_9_fu_465_node_x_coords_ce0),
    .node_x_coords_q0(node_x_coords_q0),
    .sext_ln182(n_assign_load_reg_1041)
);

kmeans_top_kmeans_top_Pipeline_10 grp_kmeans_top_Pipeline_10_fu_474(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .ap_start(grp_kmeans_top_Pipeline_10_fu_474_ap_start),
    .ap_done(grp_kmeans_top_Pipeline_10_fu_474_ap_done),
    .ap_idle(grp_kmeans_top_Pipeline_10_fu_474_ap_idle),
    .ap_ready(grp_kmeans_top_Pipeline_10_fu_474_ap_ready),
    .m_axi_mem_AWVALID(grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_AWVALID),
    .m_axi_mem_AWREADY(mem_AWREADY),
    .m_axi_mem_AWADDR(grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_AWADDR),
    .m_axi_mem_AWID(grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_AWID),
    .m_axi_mem_AWLEN(grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_AWLEN),
    .m_axi_mem_AWSIZE(grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_AWSIZE),
    .m_axi_mem_AWBURST(grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_AWBURST),
    .m_axi_mem_AWLOCK(grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_AWLOCK),
    .m_axi_mem_AWCACHE(grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_AWCACHE),
    .m_axi_mem_AWPROT(grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_AWPROT),
    .m_axi_mem_AWQOS(grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_AWQOS),
    .m_axi_mem_AWREGION(grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_AWREGION),
    .m_axi_mem_AWUSER(grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_AWUSER),
    .m_axi_mem_WVALID(grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_WVALID),
    .m_axi_mem_WREADY(mem_WREADY),
    .m_axi_mem_WDATA(grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_WDATA),
    .m_axi_mem_WSTRB(grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_WSTRB),
    .m_axi_mem_WLAST(grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_WLAST),
    .m_axi_mem_WID(grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_WID),
    .m_axi_mem_WUSER(grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_WUSER),
    .m_axi_mem_ARVALID(grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_ARVALID),
    .m_axi_mem_ARREADY(1'b0),
    .m_axi_mem_ARADDR(grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_ARADDR),
    .m_axi_mem_ARID(grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_ARID),
    .m_axi_mem_ARLEN(grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_ARLEN),
    .m_axi_mem_ARSIZE(grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_ARSIZE),
    .m_axi_mem_ARBURST(grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_ARBURST),
    .m_axi_mem_ARLOCK(grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_ARLOCK),
    .m_axi_mem_ARCACHE(grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_ARCACHE),
    .m_axi_mem_ARPROT(grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_ARPROT),
    .m_axi_mem_ARQOS(grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_ARQOS),
    .m_axi_mem_ARREGION(grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_ARREGION),
    .m_axi_mem_ARUSER(grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_ARUSER),
    .m_axi_mem_RVALID(1'b0),
    .m_axi_mem_RREADY(grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_RREADY),
    .m_axi_mem_RDATA(64'd0),
    .m_axi_mem_RLAST(1'b0),
    .m_axi_mem_RID(1'd0),
    .m_axi_mem_RFIFONUM(9'd0),
    .m_axi_mem_RUSER(1'd0),
    .m_axi_mem_RRESP(2'd0),
    .m_axi_mem_BVALID(mem_BVALID),
    .m_axi_mem_BREADY(grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_BREADY),
    .m_axi_mem_BRESP(2'd0),
    .m_axi_mem_BID(1'd0),
    .m_axi_mem_BUSER(1'd0),
    .p_cast8_cast(reg_596),
    .node_y_coords_address0(grp_kmeans_top_Pipeline_10_fu_474_node_y_coords_address0),
    .node_y_coords_ce0(grp_kmeans_top_Pipeline_10_fu_474_node_y_coords_ce0),
    .node_y_coords_q0(node_y_coords_q0),
    .sext_ln182(n_assign_load_reg_1041)
);

kmeans_top_kmeans_top_Pipeline_11 grp_kmeans_top_Pipeline_11_fu_483(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .ap_start(grp_kmeans_top_Pipeline_11_fu_483_ap_start),
    .ap_done(grp_kmeans_top_Pipeline_11_fu_483_ap_done),
    .ap_idle(grp_kmeans_top_Pipeline_11_fu_483_ap_idle),
    .ap_ready(grp_kmeans_top_Pipeline_11_fu_483_ap_ready),
    .m_axi_mem_AWVALID(grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_AWVALID),
    .m_axi_mem_AWREADY(mem_AWREADY),
    .m_axi_mem_AWADDR(grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_AWADDR),
    .m_axi_mem_AWID(grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_AWID),
    .m_axi_mem_AWLEN(grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_AWLEN),
    .m_axi_mem_AWSIZE(grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_AWSIZE),
    .m_axi_mem_AWBURST(grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_AWBURST),
    .m_axi_mem_AWLOCK(grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_AWLOCK),
    .m_axi_mem_AWCACHE(grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_AWCACHE),
    .m_axi_mem_AWPROT(grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_AWPROT),
    .m_axi_mem_AWQOS(grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_AWQOS),
    .m_axi_mem_AWREGION(grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_AWREGION),
    .m_axi_mem_AWUSER(grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_AWUSER),
    .m_axi_mem_WVALID(grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_WVALID),
    .m_axi_mem_WREADY(mem_WREADY),
    .m_axi_mem_WDATA(grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_WDATA),
    .m_axi_mem_WSTRB(grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_WSTRB),
    .m_axi_mem_WLAST(grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_WLAST),
    .m_axi_mem_WID(grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_WID),
    .m_axi_mem_WUSER(grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_WUSER),
    .m_axi_mem_ARVALID(grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_ARVALID),
    .m_axi_mem_ARREADY(1'b0),
    .m_axi_mem_ARADDR(grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_ARADDR),
    .m_axi_mem_ARID(grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_ARID),
    .m_axi_mem_ARLEN(grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_ARLEN),
    .m_axi_mem_ARSIZE(grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_ARSIZE),
    .m_axi_mem_ARBURST(grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_ARBURST),
    .m_axi_mem_ARLOCK(grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_ARLOCK),
    .m_axi_mem_ARCACHE(grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_ARCACHE),
    .m_axi_mem_ARPROT(grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_ARPROT),
    .m_axi_mem_ARQOS(grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_ARQOS),
    .m_axi_mem_ARREGION(grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_ARREGION),
    .m_axi_mem_ARUSER(grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_ARUSER),
    .m_axi_mem_RVALID(1'b0),
    .m_axi_mem_RREADY(grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_RREADY),
    .m_axi_mem_RDATA(64'd0),
    .m_axi_mem_RLAST(1'b0),
    .m_axi_mem_RID(1'd0),
    .m_axi_mem_RFIFONUM(9'd0),
    .m_axi_mem_RUSER(1'd0),
    .m_axi_mem_RRESP(2'd0),
    .m_axi_mem_BVALID(mem_BVALID),
    .m_axi_mem_BREADY(grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_BREADY),
    .m_axi_mem_BRESP(2'd0),
    .m_axi_mem_BID(1'd0),
    .m_axi_mem_BUSER(1'd0),
    .p_cast6_cast(reg_602),
    .node_cluster_assignments_address0(grp_kmeans_top_Pipeline_11_fu_483_node_cluster_assignments_address0),
    .node_cluster_assignments_ce0(grp_kmeans_top_Pipeline_11_fu_483_node_cluster_assignments_ce0),
    .node_cluster_assignments_q0(node_cluster_assignments_q0),
    .sext_ln182(n_assign_load_reg_1041)
);

kmeans_top_kmeans_top_Pipeline_12 grp_kmeans_top_Pipeline_12_fu_492(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .ap_start(grp_kmeans_top_Pipeline_12_fu_492_ap_start),
    .ap_done(grp_kmeans_top_Pipeline_12_fu_492_ap_done),
    .ap_idle(grp_kmeans_top_Pipeline_12_fu_492_ap_idle),
    .ap_ready(grp_kmeans_top_Pipeline_12_fu_492_ap_ready),
    .m_axi_mem_AWVALID(grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_AWVALID),
    .m_axi_mem_AWREADY(mem_AWREADY),
    .m_axi_mem_AWADDR(grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_AWADDR),
    .m_axi_mem_AWID(grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_AWID),
    .m_axi_mem_AWLEN(grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_AWLEN),
    .m_axi_mem_AWSIZE(grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_AWSIZE),
    .m_axi_mem_AWBURST(grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_AWBURST),
    .m_axi_mem_AWLOCK(grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_AWLOCK),
    .m_axi_mem_AWCACHE(grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_AWCACHE),
    .m_axi_mem_AWPROT(grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_AWPROT),
    .m_axi_mem_AWQOS(grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_AWQOS),
    .m_axi_mem_AWREGION(grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_AWREGION),
    .m_axi_mem_AWUSER(grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_AWUSER),
    .m_axi_mem_WVALID(grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_WVALID),
    .m_axi_mem_WREADY(mem_WREADY),
    .m_axi_mem_WDATA(grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_WDATA),
    .m_axi_mem_WSTRB(grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_WSTRB),
    .m_axi_mem_WLAST(grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_WLAST),
    .m_axi_mem_WID(grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_WID),
    .m_axi_mem_WUSER(grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_WUSER),
    .m_axi_mem_ARVALID(grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_ARVALID),
    .m_axi_mem_ARREADY(1'b0),
    .m_axi_mem_ARADDR(grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_ARADDR),
    .m_axi_mem_ARID(grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_ARID),
    .m_axi_mem_ARLEN(grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_ARLEN),
    .m_axi_mem_ARSIZE(grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_ARSIZE),
    .m_axi_mem_ARBURST(grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_ARBURST),
    .m_axi_mem_ARLOCK(grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_ARLOCK),
    .m_axi_mem_ARCACHE(grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_ARCACHE),
    .m_axi_mem_ARPROT(grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_ARPROT),
    .m_axi_mem_ARQOS(grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_ARQOS),
    .m_axi_mem_ARREGION(grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_ARREGION),
    .m_axi_mem_ARUSER(grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_ARUSER),
    .m_axi_mem_RVALID(1'b0),
    .m_axi_mem_RREADY(grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_RREADY),
    .m_axi_mem_RDATA(64'd0),
    .m_axi_mem_RLAST(1'b0),
    .m_axi_mem_RID(1'd0),
    .m_axi_mem_RFIFONUM(9'd0),
    .m_axi_mem_RUSER(1'd0),
    .m_axi_mem_RRESP(2'd0),
    .m_axi_mem_BVALID(mem_BVALID),
    .m_axi_mem_BREADY(grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_BREADY),
    .m_axi_mem_BRESP(2'd0),
    .m_axi_mem_BID(1'd0),
    .m_axi_mem_BUSER(1'd0),
    .p_cast7_cast(reg_608),
    .centroid_x_coords_address0(grp_kmeans_top_Pipeline_12_fu_492_centroid_x_coords_address0),
    .centroid_x_coords_ce0(grp_kmeans_top_Pipeline_12_fu_492_centroid_x_coords_ce0),
    .centroid_x_coords_q0(centroid_x_coords_q0),
    .sext_ln185(k_assign_load_reg_1063)
);

kmeans_top_kmeans_top_Pipeline_13 grp_kmeans_top_Pipeline_13_fu_501(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst_n_inv),
    .ap_start(grp_kmeans_top_Pipeline_13_fu_501_ap_start),
    .ap_done(grp_kmeans_top_Pipeline_13_fu_501_ap_done),
    .ap_idle(grp_kmeans_top_Pipeline_13_fu_501_ap_idle),
    .ap_ready(grp_kmeans_top_Pipeline_13_fu_501_ap_ready),
    .m_axi_mem_AWVALID(grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_AWVALID),
    .m_axi_mem_AWREADY(mem_AWREADY),
    .m_axi_mem_AWADDR(grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_AWADDR),
    .m_axi_mem_AWID(grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_AWID),
    .m_axi_mem_AWLEN(grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_AWLEN),
    .m_axi_mem_AWSIZE(grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_AWSIZE),
    .m_axi_mem_AWBURST(grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_AWBURST),
    .m_axi_mem_AWLOCK(grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_AWLOCK),
    .m_axi_mem_AWCACHE(grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_AWCACHE),
    .m_axi_mem_AWPROT(grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_AWPROT),
    .m_axi_mem_AWQOS(grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_AWQOS),
    .m_axi_mem_AWREGION(grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_AWREGION),
    .m_axi_mem_AWUSER(grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_AWUSER),
    .m_axi_mem_WVALID(grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_WVALID),
    .m_axi_mem_WREADY(mem_WREADY),
    .m_axi_mem_WDATA(grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_WDATA),
    .m_axi_mem_WSTRB(grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_WSTRB),
    .m_axi_mem_WLAST(grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_WLAST),
    .m_axi_mem_WID(grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_WID),
    .m_axi_mem_WUSER(grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_WUSER),
    .m_axi_mem_ARVALID(grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_ARVALID),
    .m_axi_mem_ARREADY(1'b0),
    .m_axi_mem_ARADDR(grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_ARADDR),
    .m_axi_mem_ARID(grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_ARID),
    .m_axi_mem_ARLEN(grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_ARLEN),
    .m_axi_mem_ARSIZE(grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_ARSIZE),
    .m_axi_mem_ARBURST(grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_ARBURST),
    .m_axi_mem_ARLOCK(grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_ARLOCK),
    .m_axi_mem_ARCACHE(grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_ARCACHE),
    .m_axi_mem_ARPROT(grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_ARPROT),
    .m_axi_mem_ARQOS(grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_ARQOS),
    .m_axi_mem_ARREGION(grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_ARREGION),
    .m_axi_mem_ARUSER(grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_ARUSER),
    .m_axi_mem_RVALID(1'b0),
    .m_axi_mem_RREADY(grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_RREADY),
    .m_axi_mem_RDATA(64'd0),
    .m_axi_mem_RLAST(1'b0),
    .m_axi_mem_RID(1'd0),
    .m_axi_mem_RFIFONUM(9'd0),
    .m_axi_mem_RUSER(1'd0),
    .m_axi_mem_RRESP(2'd0),
    .m_axi_mem_BVALID(mem_BVALID),
    .m_axi_mem_BREADY(grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_BREADY),
    .m_axi_mem_BRESP(2'd0),
    .m_axi_mem_BID(1'd0),
    .m_axi_mem_BUSER(1'd0),
    .p_cast12_cast(reg_614),
    .centroid_y_coords_address0(grp_kmeans_top_Pipeline_13_fu_501_centroid_y_coords_address0),
    .centroid_y_coords_ce0(grp_kmeans_top_Pipeline_13_fu_501_centroid_y_coords_ce0),
    .centroid_y_coords_q0(centroid_y_coords_q0),
    .sext_ln185(k_assign_load_reg_1063)
);

kmeans_top_cfg_s_axi #(
    .C_S_AXI_ADDR_WIDTH( C_S_AXI_CFG_ADDR_WIDTH ),
    .C_S_AXI_DATA_WIDTH( C_S_AXI_CFG_DATA_WIDTH ))
cfg_s_axi_U(
    .AWVALID(s_axi_cfg_AWVALID),
    .AWREADY(s_axi_cfg_AWREADY),
    .AWADDR(s_axi_cfg_AWADDR),
    .WVALID(s_axi_cfg_WVALID),
    .WREADY(s_axi_cfg_WREADY),
    .WDATA(s_axi_cfg_WDATA),
    .WSTRB(s_axi_cfg_WSTRB),
    .ARVALID(s_axi_cfg_ARVALID),
    .ARREADY(s_axi_cfg_ARREADY),
    .ARADDR(s_axi_cfg_ARADDR),
    .RVALID(s_axi_cfg_RVALID),
    .RREADY(s_axi_cfg_RREADY),
    .RDATA(s_axi_cfg_RDATA),
    .RRESP(s_axi_cfg_RRESP),
    .BVALID(s_axi_cfg_BVALID),
    .BREADY(s_axi_cfg_BREADY),
    .BRESP(s_axi_cfg_BRESP),
    .ACLK(ap_clk),
    .ARESET(ap_rst_n_inv),
    .ACLK_EN(1'b1),
    .n(n),
    .k(k),
    .control(control),
    .buf_ptr_node_x_coords(buf_ptr_node_x_coords),
    .buf_ptr_node_y_coords(buf_ptr_node_y_coords),
    .buf_ptr_node_cluster_assignments(buf_ptr_node_cluster_assignments),
    .buf_ptr_centroid_x_coords(buf_ptr_centroid_x_coords),
    .buf_ptr_centroid_y_coords(buf_ptr_centroid_y_coords),
    .buf_ptr_intermediate_cluster_assignments(buf_ptr_intermediate_cluster_assignments),
    .buf_ptr_intermediate_centroid_x_coords(buf_ptr_intermediate_centroid_x_coords),
    .buf_ptr_intermediate_centroid_y_coords(buf_ptr_intermediate_centroid_y_coords),
    .max_iterations(max_iterations),
    .sub_iterations(sub_iterations),
    .ap_start(ap_start),
    .interrupt(interrupt),
    .ap_ready(ap_ready),
    .ap_done(ap_done),
    .ap_idle(ap_idle)
);

kmeans_top_mem_m_axi #(
    .CONSERVATIVE( 1 ),
    .USER_MAXREQS( 5 ),
    .MAX_READ_BURST_LENGTH( 16 ),
    .MAX_WRITE_BURST_LENGTH( 16 ),
    .C_M_AXI_ID_WIDTH( C_M_AXI_MEM_ID_WIDTH ),
    .C_M_AXI_ADDR_WIDTH( C_M_AXI_MEM_ADDR_WIDTH ),
    .C_M_AXI_DATA_WIDTH( C_M_AXI_MEM_DATA_WIDTH ),
    .C_M_AXI_AWUSER_WIDTH( C_M_AXI_MEM_AWUSER_WIDTH ),
    .C_M_AXI_ARUSER_WIDTH( C_M_AXI_MEM_ARUSER_WIDTH ),
    .C_M_AXI_WUSER_WIDTH( C_M_AXI_MEM_WUSER_WIDTH ),
    .C_M_AXI_RUSER_WIDTH( C_M_AXI_MEM_RUSER_WIDTH ),
    .C_M_AXI_BUSER_WIDTH( C_M_AXI_MEM_BUSER_WIDTH ),
    .C_USER_VALUE( C_M_AXI_MEM_USER_VALUE ),
    .C_PROT_VALUE( C_M_AXI_MEM_PROT_VALUE ),
    .C_CACHE_VALUE( C_M_AXI_MEM_CACHE_VALUE ),
    .USER_RFIFONUM_WIDTH( 9 ),
    .USER_DW( 64 ),
    .USER_AW( 64 ),
    .NUM_READ_OUTSTANDING( 16 ),
    .NUM_WRITE_OUTSTANDING( 16 ))
mem_m_axi_U(
    .AWVALID(m_axi_mem_AWVALID),
    .AWREADY(m_axi_mem_AWREADY),
    .AWADDR(m_axi_mem_AWADDR),
    .AWID(m_axi_mem_AWID),
    .AWLEN(m_axi_mem_AWLEN),
    .AWSIZE(m_axi_mem_AWSIZE),
    .AWBURST(m_axi_mem_AWBURST),
    .AWLOCK(m_axi_mem_AWLOCK),
    .AWCACHE(m_axi_mem_AWCACHE),
    .AWPROT(m_axi_mem_AWPROT),
    .AWQOS(m_axi_mem_AWQOS),
    .AWREGION(m_axi_mem_AWREGION),
    .AWUSER(m_axi_mem_AWUSER),
    .WVALID(m_axi_mem_WVALID),
    .WREADY(m_axi_mem_WREADY),
    .WDATA(m_axi_mem_WDATA),
    .WSTRB(m_axi_mem_WSTRB),
    .WLAST(m_axi_mem_WLAST),
    .WID(m_axi_mem_WID),
    .WUSER(m_axi_mem_WUSER),
    .ARVALID(m_axi_mem_ARVALID),
    .ARREADY(m_axi_mem_ARREADY),
    .ARADDR(m_axi_mem_ARADDR),
    .ARID(m_axi_mem_ARID),
    .ARLEN(m_axi_mem_ARLEN),
    .ARSIZE(m_axi_mem_ARSIZE),
    .ARBURST(m_axi_mem_ARBURST),
    .ARLOCK(m_axi_mem_ARLOCK),
    .ARCACHE(m_axi_mem_ARCACHE),
    .ARPROT(m_axi_mem_ARPROT),
    .ARQOS(m_axi_mem_ARQOS),
    .ARREGION(m_axi_mem_ARREGION),
    .ARUSER(m_axi_mem_ARUSER),
    .RVALID(m_axi_mem_RVALID),
    .RREADY(m_axi_mem_RREADY),
    .RDATA(m_axi_mem_RDATA),
    .RLAST(m_axi_mem_RLAST),
    .RID(m_axi_mem_RID),
    .RUSER(m_axi_mem_RUSER),
    .RRESP(m_axi_mem_RRESP),
    .BVALID(m_axi_mem_BVALID),
    .BREADY(m_axi_mem_BREADY),
    .BRESP(m_axi_mem_BRESP),
    .BID(m_axi_mem_BID),
    .BUSER(m_axi_mem_BUSER),
    .ACLK(ap_clk),
    .ARESET(ap_rst_n_inv),
    .ACLK_EN(1'b1),
    .I_ARVALID(mem_ARVALID),
    .I_ARREADY(mem_ARREADY),
    .I_ARADDR(mem_ARADDR),
    .I_ARLEN(mem_ARLEN),
    .I_RVALID(mem_RVALID),
    .I_RREADY(mem_RREADY),
    .I_RDATA(mem_RDATA),
    .I_RFIFONUM(mem_RFIFONUM),
    .I_AWVALID(mem_AWVALID),
    .I_AWREADY(mem_AWREADY),
    .I_AWADDR(mem_AWADDR),
    .I_AWLEN(mem_AWLEN),
    .I_WVALID(mem_WVALID),
    .I_WREADY(mem_WREADY),
    .I_WDATA(mem_WDATA),
    .I_WSTRB(mem_WSTRB),
    .I_BVALID(mem_BVALID),
    .I_BREADY(mem_BREADY)
);

kmeans_top_mul_29s_29s_29_1_1 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 29 ),
    .din1_WIDTH( 29 ),
    .dout_WIDTH( 29 ))
mul_29s_29s_29_1_1_U89(
    .din0(mul_ln194_fu_776_p0),
    .din1(mul_ln194_fu_776_p1),
    .dout(mul_ln194_fu_776_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        grp_kmeans_fu_426_ap_start_reg <= 1'b0;
    end else begin
        if (((ap_phi_mux_phi_ln191_phi_fu_374_p4 == 1'd0) & (icmp_ln191_fu_738_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state47))) begin
            grp_kmeans_fu_426_ap_start_reg <= 1'b1;
        end else if ((grp_kmeans_fu_426_ap_ready == 1'b1)) begin
            grp_kmeans_fu_426_ap_start_reg <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        grp_kmeans_top_Pipeline_10_fu_474_ap_start_reg <= 1'b0;
    end else begin
        if (((1'b1 == ap_CS_fsm_state79) & (1'b1 == ap_NS_fsm_state80))) begin
            grp_kmeans_top_Pipeline_10_fu_474_ap_start_reg <= 1'b1;
        end else if ((grp_kmeans_top_Pipeline_10_fu_474_ap_ready == 1'b1)) begin
            grp_kmeans_top_Pipeline_10_fu_474_ap_start_reg <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        grp_kmeans_top_Pipeline_11_fu_483_ap_start_reg <= 1'b0;
    end else begin
        if (((1'b1 == ap_CS_fsm_state86) & (1'b1 == ap_NS_fsm_state87))) begin
            grp_kmeans_top_Pipeline_11_fu_483_ap_start_reg <= 1'b1;
        end else if ((grp_kmeans_top_Pipeline_11_fu_483_ap_ready == 1'b1)) begin
            grp_kmeans_top_Pipeline_11_fu_483_ap_start_reg <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        grp_kmeans_top_Pipeline_12_fu_492_ap_start_reg <= 1'b0;
    end else begin
        if (((1'b1 == ap_CS_fsm_state93) & (1'b1 == ap_NS_fsm_state94))) begin
            grp_kmeans_top_Pipeline_12_fu_492_ap_start_reg <= 1'b1;
        end else if ((grp_kmeans_top_Pipeline_12_fu_492_ap_ready == 1'b1)) begin
            grp_kmeans_top_Pipeline_12_fu_492_ap_start_reg <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        grp_kmeans_top_Pipeline_13_fu_501_ap_start_reg <= 1'b0;
    end else begin
        if (((1'b1 == ap_CS_fsm_state100) & (1'b1 == ap_NS_fsm_state101))) begin
            grp_kmeans_top_Pipeline_13_fu_501_ap_start_reg <= 1'b1;
        end else if ((grp_kmeans_top_Pipeline_13_fu_501_ap_ready == 1'b1)) begin
            grp_kmeans_top_Pipeline_13_fu_501_ap_start_reg <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        grp_kmeans_top_Pipeline_1_fu_381_ap_start_reg <= 1'b0;
    end else begin
        if (((1'b1 == ap_NS_fsm_state9) & (1'b1 == ap_CS_fsm_state8))) begin
            grp_kmeans_top_Pipeline_1_fu_381_ap_start_reg <= 1'b1;
        end else if ((grp_kmeans_top_Pipeline_1_fu_381_ap_ready == 1'b1)) begin
            grp_kmeans_top_Pipeline_1_fu_381_ap_start_reg <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        grp_kmeans_top_Pipeline_2_fu_390_ap_start_reg <= 1'b0;
    end else begin
        if (((1'b1 == ap_NS_fsm_state18) & (1'b1 == ap_CS_fsm_state17))) begin
            grp_kmeans_top_Pipeline_2_fu_390_ap_start_reg <= 1'b1;
        end else if ((grp_kmeans_top_Pipeline_2_fu_390_ap_ready == 1'b1)) begin
            grp_kmeans_top_Pipeline_2_fu_390_ap_start_reg <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        grp_kmeans_top_Pipeline_3_fu_399_ap_start_reg <= 1'b0;
    end else begin
        if (((1'b1 == ap_NS_fsm_state27) & (1'b1 == ap_CS_fsm_state26))) begin
            grp_kmeans_top_Pipeline_3_fu_399_ap_start_reg <= 1'b1;
        end else if ((grp_kmeans_top_Pipeline_3_fu_399_ap_ready == 1'b1)) begin
            grp_kmeans_top_Pipeline_3_fu_399_ap_start_reg <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        grp_kmeans_top_Pipeline_4_fu_408_ap_start_reg <= 1'b0;
    end else begin
        if (((1'b1 == ap_NS_fsm_state36) & (1'b1 == ap_CS_fsm_state35))) begin
            grp_kmeans_top_Pipeline_4_fu_408_ap_start_reg <= 1'b1;
        end else if ((grp_kmeans_top_Pipeline_4_fu_408_ap_ready == 1'b1)) begin
            grp_kmeans_top_Pipeline_4_fu_408_ap_start_reg <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        grp_kmeans_top_Pipeline_5_fu_417_ap_start_reg <= 1'b0;
    end else begin
        if (((1'b1 == ap_NS_fsm_state45) & (1'b1 == ap_CS_fsm_state44))) begin
            grp_kmeans_top_Pipeline_5_fu_417_ap_start_reg <= 1'b1;
        end else if ((grp_kmeans_top_Pipeline_5_fu_417_ap_ready == 1'b1)) begin
            grp_kmeans_top_Pipeline_5_fu_417_ap_start_reg <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        grp_kmeans_top_Pipeline_6_fu_438_ap_start_reg <= 1'b0;
    end else begin
        if (((1'b1 == ap_CS_fsm_state49) & (1'b1 == ap_NS_fsm_state50))) begin
            grp_kmeans_top_Pipeline_6_fu_438_ap_start_reg <= 1'b1;
        end else if ((grp_kmeans_top_Pipeline_6_fu_438_ap_ready == 1'b1)) begin
            grp_kmeans_top_Pipeline_6_fu_438_ap_start_reg <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        grp_kmeans_top_Pipeline_7_fu_447_ap_start_reg <= 1'b0;
    end else begin
        if (((1'b1 == ap_CS_fsm_state57) & (1'b1 == ap_NS_fsm_state58))) begin
            grp_kmeans_top_Pipeline_7_fu_447_ap_start_reg <= 1'b1;
        end else if ((grp_kmeans_top_Pipeline_7_fu_447_ap_ready == 1'b1)) begin
            grp_kmeans_top_Pipeline_7_fu_447_ap_start_reg <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        grp_kmeans_top_Pipeline_8_fu_456_ap_start_reg <= 1'b0;
    end else begin
        if (((1'b1 == ap_CS_fsm_state64) & (1'b1 == ap_NS_fsm_state65))) begin
            grp_kmeans_top_Pipeline_8_fu_456_ap_start_reg <= 1'b1;
        end else if ((grp_kmeans_top_Pipeline_8_fu_456_ap_ready == 1'b1)) begin
            grp_kmeans_top_Pipeline_8_fu_456_ap_start_reg <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst_n_inv == 1'b1) begin
        grp_kmeans_top_Pipeline_9_fu_465_ap_start_reg <= 1'b0;
    end else begin
        if (((1'b1 == ap_CS_fsm_state72) & (1'b1 == ap_NS_fsm_state73))) begin
            grp_kmeans_top_Pipeline_9_fu_465_ap_start_reg <= 1'b1;
        end else if ((grp_kmeans_top_Pipeline_9_fu_465_ap_ready == 1'b1)) begin
            grp_kmeans_top_Pipeline_9_fu_465_ap_start_reg <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_state46) & (1'b0 == ap_block_state46_on_subcall_done))) begin
        current_iteration_fu_202 <= 32'd0;
    end else if ((~((ap_predicate_op334_writeresp_state71 == 1'b1) & (mem_BVALID == 1'b0)) & (1'b1 == ap_CS_fsm_state71))) begin
        current_iteration_fu_202 <= current_iteration_1_fu_895_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_state46) & (1'b0 == ap_block_state46_on_subcall_done))) begin
        intermediate_writes_made_fu_198 <= 32'd0;
    end else if ((~((ap_predicate_op334_writeresp_state71 == 1'b1) & (mem_BVALID == 1'b0)) & (1'b1 == ap_CS_fsm_state71))) begin
        intermediate_writes_made_fu_198 <= intermediate_writes_made_2_reg_1123;
    end
end

always @ (posedge ap_clk) begin
    if ((~((ap_predicate_op334_writeresp_state71 == 1'b1) & (mem_BVALID == 1'b0)) & (1'b1 == ap_CS_fsm_state71))) begin
        phi_ln191_reg_370 <= converged_reg_1156;
    end else if (((1'b1 == ap_CS_fsm_state46) & (1'b0 == ap_block_state46_on_subcall_done))) begin
        phi_ln191_reg_370 <= 1'd0;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        buf_ptr_centroid_x_coords_read_reg_989 <= buf_ptr_centroid_x_coords;
        buf_ptr_centroid_y_coords_read_reg_984 <= buf_ptr_centroid_y_coords;
        buf_ptr_intermediate_centroid_x_coords_read_reg_974 <= buf_ptr_intermediate_centroid_x_coords;
        buf_ptr_intermediate_centroid_y_coords_read_reg_969 <= buf_ptr_intermediate_centroid_y_coords;
        buf_ptr_intermediate_cluster_assignments_read_reg_979 <= buf_ptr_intermediate_cluster_assignments;
        buf_ptr_node_cluster_assignments_read_reg_994 <= buf_ptr_node_cluster_assignments;
        buf_ptr_node_x_coords_read_reg_1004 <= buf_ptr_node_x_coords;
        buf_ptr_node_y_coords_read_reg_999 <= buf_ptr_node_y_coords;
        icmp_ln185_reg_1059 <= icmp_ln185_fu_649_p2;
        n_assign_load_reg_1041 <= grp_load_fu_510_p1;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
        control_assign_fu_166 <= trunc_ln131_fu_620_p1;
        k_assign_fu_162 <= k;
        max_iterations_assign_fu_170 <= max_iterations;
        n_assign_fu_158 <= n;
        sub_iterations_assign_fu_174 <= sub_iterations;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state48)) begin
        converged_reg_1156 <= grp_kmeans_fu_426_ap_return;
        tmp_reg_1161 <= control_assign_fu_166[32'd1];
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state28)) begin
        icmp_ln188_reg_1095 <= icmp_ln188_fu_688_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((grp_fu_576_p3 == 1'd1) & (1'b1 == ap_CS_fsm_state48))) begin
        icmp_ln196_reg_1165 <= grp_fu_584_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln199_fu_826_p1 == 1'd1) & (1'b1 == ap_CS_fsm_state56))) begin
        icmp_ln199_reg_1184 <= grp_fu_584_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state47)) begin
        intermediate_writes_made_2_reg_1123 <= intermediate_writes_made_2_fu_728_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_phi_mux_phi_ln191_phi_fu_374_p4 == 1'd0) & (icmp_ln191_fu_738_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state47))) begin
        k_assign_load_1_reg_1141 <= k_assign_fu_162;
        mul_ln194_reg_1146 <= mul_ln194_fu_776_p2;
        n_assign_load_1_reg_1136 <= grp_load_fu_510_p1;
        sub_iterations_assign_load_reg_1131 <= sub_iterations_assign_fu_174;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        k_assign_load_reg_1063 <= k_assign_fu_162;
    end
end

always @ (posedge ap_clk) begin
    if (((trunc_ln199_fu_826_p1 == 1'd1) & (grp_fu_584_p2 == 1'd1) & (icmp_ln188_reg_1095 == 1'd1) & (1'b1 == ap_CS_fsm_state56))) begin
        p_cast10_reg_1188 <= {{empty_53_fu_841_p2[63:3]}};
        p_cast11_reg_1194 <= {{empty_56_fu_856_p2[63:3]}};
    end
end

always @ (posedge ap_clk) begin
    if (((grp_fu_584_p2 == 1'd1) & (grp_fu_576_p3 == 1'd1) & (1'b1 == ap_CS_fsm_state48) & (icmp_ln185_reg_1059 == 1'd1))) begin
        p_cast9_reg_1169 <= {{empty_50_fu_801_p2[63:3]}};
    end
end

always @ (posedge ap_clk) begin
    if ((((1'b1 == ap_CS_fsm_state47) & (((ap_phi_mux_phi_ln191_phi_fu_374_p4 == 1'd1) & (tmp_3_fu_782_p3 == 1'd1) & (icmp_ln185_reg_1059 == 1'd1)) | ((tmp_3_fu_782_p3 == 1'd1) & (icmp_ln191_fu_738_p2 == 1'd0) & (icmp_ln185_reg_1059 == 1'd1)))) | ((1'b1 == ap_CS_fsm_state2) & (icmp_ln185_reg_1059 == 1'd1)))) begin
        reg_590 <= {{buf_ptr_node_x_coords_read_reg_1004[63:3]}};
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_state11) | ((1'b1 == ap_CS_fsm_state47) & (((ap_phi_mux_phi_ln191_phi_fu_374_p4 == 1'd1) & (tmp_3_fu_782_p3 == 1'd1) & (icmp_ln185_reg_1059 == 1'd1)) | ((tmp_3_fu_782_p3 == 1'd1) & (icmp_ln191_fu_738_p2 == 1'd0) & (icmp_ln185_reg_1059 == 1'd1)))))) begin
        reg_596 <= {{buf_ptr_node_y_coords_read_reg_999[63:3]}};
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_state20) | ((grp_fu_576_p3 == 1'd1) & (1'b1 == ap_CS_fsm_state86) & (icmp_ln185_reg_1059 == 1'd1)))) begin
        reg_602 <= {{buf_ptr_node_cluster_assignments_read_reg_994[63:3]}};
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_state29) | ((trunc_ln215_fu_943_p1 == 1'd1) & (icmp_ln188_reg_1095 == 1'd1) & (1'b1 == ap_CS_fsm_state93)))) begin
        reg_608 <= {{buf_ptr_centroid_x_coords_read_reg_989[63:3]}};
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_state38) | ((trunc_ln215_fu_943_p1 == 1'd1) & (icmp_ln188_reg_1095 == 1'd1) & (1'b1 == ap_CS_fsm_state93)))) begin
        reg_614 <= {{buf_ptr_centroid_y_coords_read_reg_984[63:3]}};
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_state47) & ((ap_phi_mux_phi_ln191_phi_fu_374_p4 == 1'd1) | (icmp_ln191_fu_738_p2 == 1'd0)))) begin
        tmp_3_reg_1152 <= control_assign_fu_166[32'd2];
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state86)) begin
        tmp_4_reg_1220 <= control_assign_fu_166[32'd1];
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state56)) begin
        trunc_ln199_reg_1180 <= trunc_ln199_fu_826_p1;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state93)) begin
        trunc_ln215_reg_1229 <= trunc_ln215_fu_943_p1;
    end
end

always @ (*) begin
    if (((mem_BVALID == 1'b0) | (mem_AWREADY == 1'b0))) begin
        ap_ST_fsm_state100_blk = 1'b1;
    end else begin
        ap_ST_fsm_state100_blk = 1'b0;
    end
end

assign ap_ST_fsm_state101_blk = 1'b0;

always @ (*) begin
    if ((grp_kmeans_top_Pipeline_13_fu_501_ap_done == 1'b0)) begin
        ap_ST_fsm_state102_blk = 1'b1;
    end else begin
        ap_ST_fsm_state102_blk = 1'b0;
    end
end

assign ap_ST_fsm_state103_blk = 1'b0;

assign ap_ST_fsm_state104_blk = 1'b0;

assign ap_ST_fsm_state105_blk = 1'b0;

assign ap_ST_fsm_state106_blk = 1'b0;

always @ (*) begin
    if (((ap_predicate_op408_writeresp_state107 == 1'b1) & (mem_BVALID == 1'b0))) begin
        ap_ST_fsm_state107_blk = 1'b1;
    end else begin
        ap_ST_fsm_state107_blk = 1'b0;
    end
end

always @ (*) begin
    if ((grp_kmeans_top_Pipeline_1_fu_381_ap_done == 1'b0)) begin
        ap_ST_fsm_state10_blk = 1'b1;
    end else begin
        ap_ST_fsm_state10_blk = 1'b0;
    end
end

always @ (*) begin
    if ((mem_ARREADY == 1'b0)) begin
        ap_ST_fsm_state11_blk = 1'b1;
    end else begin
        ap_ST_fsm_state11_blk = 1'b0;
    end
end

assign ap_ST_fsm_state12_blk = 1'b0;

assign ap_ST_fsm_state13_blk = 1'b0;

assign ap_ST_fsm_state14_blk = 1'b0;

assign ap_ST_fsm_state15_blk = 1'b0;

assign ap_ST_fsm_state16_blk = 1'b0;

assign ap_ST_fsm_state17_blk = 1'b0;

assign ap_ST_fsm_state18_blk = 1'b0;

always @ (*) begin
    if ((grp_kmeans_top_Pipeline_2_fu_390_ap_done == 1'b0)) begin
        ap_ST_fsm_state19_blk = 1'b1;
    end else begin
        ap_ST_fsm_state19_blk = 1'b0;
    end
end

always @ (*) begin
    if ((ap_start == 1'b0)) begin
        ap_ST_fsm_state1_blk = 1'b1;
    end else begin
        ap_ST_fsm_state1_blk = 1'b0;
    end
end

always @ (*) begin
    if ((mem_ARREADY == 1'b0)) begin
        ap_ST_fsm_state20_blk = 1'b1;
    end else begin
        ap_ST_fsm_state20_blk = 1'b0;
    end
end

assign ap_ST_fsm_state21_blk = 1'b0;

assign ap_ST_fsm_state22_blk = 1'b0;

assign ap_ST_fsm_state23_blk = 1'b0;

assign ap_ST_fsm_state24_blk = 1'b0;

assign ap_ST_fsm_state25_blk = 1'b0;

assign ap_ST_fsm_state26_blk = 1'b0;

assign ap_ST_fsm_state27_blk = 1'b0;

always @ (*) begin
    if ((1'b1 == ap_block_state28_on_subcall_done)) begin
        ap_ST_fsm_state28_blk = 1'b1;
    end else begin
        ap_ST_fsm_state28_blk = 1'b0;
    end
end

always @ (*) begin
    if ((mem_ARREADY == 1'b0)) begin
        ap_ST_fsm_state29_blk = 1'b1;
    end else begin
        ap_ST_fsm_state29_blk = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_block_state2_io)) begin
        ap_ST_fsm_state2_blk = 1'b1;
    end else begin
        ap_ST_fsm_state2_blk = 1'b0;
    end
end

assign ap_ST_fsm_state30_blk = 1'b0;

assign ap_ST_fsm_state31_blk = 1'b0;

assign ap_ST_fsm_state32_blk = 1'b0;

assign ap_ST_fsm_state33_blk = 1'b0;

assign ap_ST_fsm_state34_blk = 1'b0;

assign ap_ST_fsm_state35_blk = 1'b0;

assign ap_ST_fsm_state36_blk = 1'b0;

always @ (*) begin
    if ((grp_kmeans_top_Pipeline_4_fu_408_ap_done == 1'b0)) begin
        ap_ST_fsm_state37_blk = 1'b1;
    end else begin
        ap_ST_fsm_state37_blk = 1'b0;
    end
end

always @ (*) begin
    if ((mem_ARREADY == 1'b0)) begin
        ap_ST_fsm_state38_blk = 1'b1;
    end else begin
        ap_ST_fsm_state38_blk = 1'b0;
    end
end

assign ap_ST_fsm_state39_blk = 1'b0;

assign ap_ST_fsm_state3_blk = 1'b0;

assign ap_ST_fsm_state40_blk = 1'b0;

assign ap_ST_fsm_state41_blk = 1'b0;

assign ap_ST_fsm_state42_blk = 1'b0;

assign ap_ST_fsm_state43_blk = 1'b0;

assign ap_ST_fsm_state44_blk = 1'b0;

assign ap_ST_fsm_state45_blk = 1'b0;

always @ (*) begin
    if ((1'b1 == ap_block_state46_on_subcall_done)) begin
        ap_ST_fsm_state46_blk = 1'b1;
    end else begin
        ap_ST_fsm_state46_blk = 1'b0;
    end
end

assign ap_ST_fsm_state47_blk = 1'b0;

always @ (*) begin
    if ((grp_kmeans_fu_426_ap_done == 1'b0)) begin
        ap_ST_fsm_state48_blk = 1'b1;
    end else begin
        ap_ST_fsm_state48_blk = 1'b0;
    end
end

always @ (*) begin
    if ((mem_AWREADY == 1'b0)) begin
        ap_ST_fsm_state49_blk = 1'b1;
    end else begin
        ap_ST_fsm_state49_blk = 1'b0;
    end
end

assign ap_ST_fsm_state4_blk = 1'b0;

assign ap_ST_fsm_state50_blk = 1'b0;

always @ (*) begin
    if ((grp_kmeans_top_Pipeline_6_fu_438_ap_done == 1'b0)) begin
        ap_ST_fsm_state51_blk = 1'b1;
    end else begin
        ap_ST_fsm_state51_blk = 1'b0;
    end
end

assign ap_ST_fsm_state52_blk = 1'b0;

assign ap_ST_fsm_state53_blk = 1'b0;

assign ap_ST_fsm_state54_blk = 1'b0;

assign ap_ST_fsm_state55_blk = 1'b0;

always @ (*) begin
    if (((ap_predicate_op298_writeresp_state56 == 1'b1) & (mem_BVALID == 1'b0))) begin
        ap_ST_fsm_state56_blk = 1'b1;
    end else begin
        ap_ST_fsm_state56_blk = 1'b0;
    end
end

always @ (*) begin
    if ((mem_AWREADY == 1'b0)) begin
        ap_ST_fsm_state57_blk = 1'b1;
    end else begin
        ap_ST_fsm_state57_blk = 1'b0;
    end
end

assign ap_ST_fsm_state58_blk = 1'b0;

always @ (*) begin
    if ((grp_kmeans_top_Pipeline_7_fu_447_ap_done == 1'b0)) begin
        ap_ST_fsm_state59_blk = 1'b1;
    end else begin
        ap_ST_fsm_state59_blk = 1'b0;
    end
end

assign ap_ST_fsm_state5_blk = 1'b0;

assign ap_ST_fsm_state60_blk = 1'b0;

assign ap_ST_fsm_state61_blk = 1'b0;

assign ap_ST_fsm_state62_blk = 1'b0;

assign ap_ST_fsm_state63_blk = 1'b0;

always @ (*) begin
    if (((mem_BVALID == 1'b0) | (mem_AWREADY == 1'b0))) begin
        ap_ST_fsm_state64_blk = 1'b1;
    end else begin
        ap_ST_fsm_state64_blk = 1'b0;
    end
end

assign ap_ST_fsm_state65_blk = 1'b0;

always @ (*) begin
    if ((grp_kmeans_top_Pipeline_8_fu_456_ap_done == 1'b0)) begin
        ap_ST_fsm_state66_blk = 1'b1;
    end else begin
        ap_ST_fsm_state66_blk = 1'b0;
    end
end

assign ap_ST_fsm_state67_blk = 1'b0;

assign ap_ST_fsm_state68_blk = 1'b0;

assign ap_ST_fsm_state69_blk = 1'b0;

assign ap_ST_fsm_state6_blk = 1'b0;

assign ap_ST_fsm_state70_blk = 1'b0;

always @ (*) begin
    if (((ap_predicate_op334_writeresp_state71 == 1'b1) & (mem_BVALID == 1'b0))) begin
        ap_ST_fsm_state71_blk = 1'b1;
    end else begin
        ap_ST_fsm_state71_blk = 1'b0;
    end
end

always @ (*) begin
    if ((mem_AWREADY == 1'b0)) begin
        ap_ST_fsm_state72_blk = 1'b1;
    end else begin
        ap_ST_fsm_state72_blk = 1'b0;
    end
end

assign ap_ST_fsm_state73_blk = 1'b0;

always @ (*) begin
    if ((grp_kmeans_top_Pipeline_9_fu_465_ap_done == 1'b0)) begin
        ap_ST_fsm_state74_blk = 1'b1;
    end else begin
        ap_ST_fsm_state74_blk = 1'b0;
    end
end

assign ap_ST_fsm_state75_blk = 1'b0;

assign ap_ST_fsm_state76_blk = 1'b0;

assign ap_ST_fsm_state77_blk = 1'b0;

assign ap_ST_fsm_state78_blk = 1'b0;

always @ (*) begin
    if (((mem_BVALID == 1'b0) | (mem_AWREADY == 1'b0))) begin
        ap_ST_fsm_state79_blk = 1'b1;
    end else begin
        ap_ST_fsm_state79_blk = 1'b0;
    end
end

assign ap_ST_fsm_state7_blk = 1'b0;

assign ap_ST_fsm_state80_blk = 1'b0;

always @ (*) begin
    if ((grp_kmeans_top_Pipeline_10_fu_474_ap_done == 1'b0)) begin
        ap_ST_fsm_state81_blk = 1'b1;
    end else begin
        ap_ST_fsm_state81_blk = 1'b0;
    end
end

assign ap_ST_fsm_state82_blk = 1'b0;

assign ap_ST_fsm_state83_blk = 1'b0;

assign ap_ST_fsm_state84_blk = 1'b0;

assign ap_ST_fsm_state85_blk = 1'b0;

always @ (*) begin
    if (((1'b1 == ap_block_state86_io) | ((ap_predicate_op363_writeresp_state86 == 1'b1) & (mem_BVALID == 1'b0)))) begin
        ap_ST_fsm_state86_blk = 1'b1;
    end else begin
        ap_ST_fsm_state86_blk = 1'b0;
    end
end

assign ap_ST_fsm_state87_blk = 1'b0;

always @ (*) begin
    if ((grp_kmeans_top_Pipeline_11_fu_483_ap_done == 1'b0)) begin
        ap_ST_fsm_state88_blk = 1'b1;
    end else begin
        ap_ST_fsm_state88_blk = 1'b0;
    end
end

assign ap_ST_fsm_state89_blk = 1'b0;

assign ap_ST_fsm_state8_blk = 1'b0;

assign ap_ST_fsm_state90_blk = 1'b0;

assign ap_ST_fsm_state91_blk = 1'b0;

assign ap_ST_fsm_state92_blk = 1'b0;

always @ (*) begin
    if (((1'b1 == ap_block_state93_io) | ((ap_predicate_op380_writeresp_state93 == 1'b1) & (mem_BVALID == 1'b0)))) begin
        ap_ST_fsm_state93_blk = 1'b1;
    end else begin
        ap_ST_fsm_state93_blk = 1'b0;
    end
end

assign ap_ST_fsm_state94_blk = 1'b0;

always @ (*) begin
    if ((grp_kmeans_top_Pipeline_12_fu_492_ap_done == 1'b0)) begin
        ap_ST_fsm_state95_blk = 1'b1;
    end else begin
        ap_ST_fsm_state95_blk = 1'b0;
    end
end

assign ap_ST_fsm_state96_blk = 1'b0;

assign ap_ST_fsm_state97_blk = 1'b0;

assign ap_ST_fsm_state98_blk = 1'b0;

assign ap_ST_fsm_state99_blk = 1'b0;

assign ap_ST_fsm_state9_blk = 1'b0;

always @ (*) begin
    if ((~((ap_predicate_op408_writeresp_state107 == 1'b1) & (mem_BVALID == 1'b0)) & (1'b1 == ap_CS_fsm_state107))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_predicate_op408_writeresp_state107 == 1'b1) & (mem_BVALID == 1'b0)) & (1'b1 == ap_CS_fsm_state107))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        ap_sig_allocacmp_n_assign_load = n;
    end else begin
        ap_sig_allocacmp_n_assign_load = n_assign_fu_158;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state95)) begin
        centroid_x_coords_address0 = grp_kmeans_top_Pipeline_12_fu_492_centroid_x_coords_address0;
    end else if ((1'b1 == ap_CS_fsm_state59)) begin
        centroid_x_coords_address0 = grp_kmeans_top_Pipeline_7_fu_447_centroid_x_coords_address0;
    end else if ((1'b1 == ap_CS_fsm_state48)) begin
        centroid_x_coords_address0 = grp_kmeans_fu_426_centroid_x_coords_address0;
    end else if ((1'b1 == ap_CS_fsm_state37)) begin
        centroid_x_coords_address0 = grp_kmeans_top_Pipeline_4_fu_408_centroid_x_coords_address0;
    end else begin
        centroid_x_coords_address0 = 'bx;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state95)) begin
        centroid_x_coords_ce0 = grp_kmeans_top_Pipeline_12_fu_492_centroid_x_coords_ce0;
    end else if ((1'b1 == ap_CS_fsm_state59)) begin
        centroid_x_coords_ce0 = grp_kmeans_top_Pipeline_7_fu_447_centroid_x_coords_ce0;
    end else if ((1'b1 == ap_CS_fsm_state48)) begin
        centroid_x_coords_ce0 = grp_kmeans_fu_426_centroid_x_coords_ce0;
    end else if ((1'b1 == ap_CS_fsm_state37)) begin
        centroid_x_coords_ce0 = grp_kmeans_top_Pipeline_4_fu_408_centroid_x_coords_ce0;
    end else begin
        centroid_x_coords_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state48)) begin
        centroid_x_coords_ce1 = grp_kmeans_fu_426_centroid_x_coords_ce1;
    end else begin
        centroid_x_coords_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state48)) begin
        centroid_x_coords_d0 = grp_kmeans_fu_426_centroid_x_coords_d0;
    end else if ((1'b1 == ap_CS_fsm_state37)) begin
        centroid_x_coords_d0 = grp_kmeans_top_Pipeline_4_fu_408_centroid_x_coords_d0;
    end else begin
        centroid_x_coords_d0 = 'bx;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state48)) begin
        centroid_x_coords_we0 = grp_kmeans_fu_426_centroid_x_coords_we0;
    end else if ((1'b1 == ap_CS_fsm_state37)) begin
        centroid_x_coords_we0 = grp_kmeans_top_Pipeline_4_fu_408_centroid_x_coords_we0;
    end else begin
        centroid_x_coords_we0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state102)) begin
        centroid_y_coords_address0 = grp_kmeans_top_Pipeline_13_fu_501_centroid_y_coords_address0;
    end else if ((1'b1 == ap_CS_fsm_state66)) begin
        centroid_y_coords_address0 = grp_kmeans_top_Pipeline_8_fu_456_centroid_y_coords_address0;
    end else if ((1'b1 == ap_CS_fsm_state48)) begin
        centroid_y_coords_address0 = grp_kmeans_fu_426_centroid_y_coords_address0;
    end else if (((icmp_ln188_reg_1095 == 1'd1) & (1'b1 == ap_CS_fsm_state46))) begin
        centroid_y_coords_address0 = grp_kmeans_top_Pipeline_5_fu_417_centroid_y_coords_address0;
    end else begin
        centroid_y_coords_address0 = 'bx;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state102)) begin
        centroid_y_coords_ce0 = grp_kmeans_top_Pipeline_13_fu_501_centroid_y_coords_ce0;
    end else if ((1'b1 == ap_CS_fsm_state66)) begin
        centroid_y_coords_ce0 = grp_kmeans_top_Pipeline_8_fu_456_centroid_y_coords_ce0;
    end else if ((1'b1 == ap_CS_fsm_state48)) begin
        centroid_y_coords_ce0 = grp_kmeans_fu_426_centroid_y_coords_ce0;
    end else if (((icmp_ln188_reg_1095 == 1'd1) & (1'b1 == ap_CS_fsm_state46))) begin
        centroid_y_coords_ce0 = grp_kmeans_top_Pipeline_5_fu_417_centroid_y_coords_ce0;
    end else begin
        centroid_y_coords_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state48)) begin
        centroid_y_coords_ce1 = grp_kmeans_fu_426_centroid_y_coords_ce1;
    end else begin
        centroid_y_coords_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state48)) begin
        centroid_y_coords_d0 = grp_kmeans_fu_426_centroid_y_coords_d0;
    end else if (((icmp_ln188_reg_1095 == 1'd1) & (1'b1 == ap_CS_fsm_state46))) begin
        centroid_y_coords_d0 = grp_kmeans_top_Pipeline_5_fu_417_centroid_y_coords_d0;
    end else begin
        centroid_y_coords_d0 = 'bx;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state48)) begin
        centroid_y_coords_we0 = grp_kmeans_fu_426_centroid_y_coords_we0;
    end else if (((icmp_ln188_reg_1095 == 1'd1) & (1'b1 == ap_CS_fsm_state46))) begin
        centroid_y_coords_we0 = grp_kmeans_top_Pipeline_5_fu_417_centroid_y_coords_we0;
    end else begin
        centroid_y_coords_we0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_phi_mux_phi_ln191_phi_fu_374_p4 == 1'd0) & (icmp_ln191_fu_738_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state47))) begin
        grp_load_fu_510_p1 = n_assign_fu_158;
    end else if ((1'b1 == ap_CS_fsm_state1)) begin
        grp_load_fu_510_p1 = ap_sig_allocacmp_n_assign_load;
    end else begin
        grp_load_fu_510_p1 = 'bx;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state38) & (mem_ARREADY == 1'b1))) begin
        mem_ARADDR = p_cast3_cast_fu_704_p1;
    end else if (((1'b1 == ap_CS_fsm_state29) & (mem_ARREADY == 1'b1))) begin
        mem_ARADDR = p_cast1_cast_fu_693_p1;
    end else if (((1'b1 == ap_CS_fsm_state20) & (mem_ARREADY == 1'b1))) begin
        mem_ARADDR = p_cast4_cast_fu_677_p1;
    end else if (((1'b1 == ap_CS_fsm_state11) & (mem_ARREADY == 1'b1))) begin
        mem_ARADDR = p_cast2_cast_fu_666_p1;
    end else if (((1'b1 == ap_CS_fsm_state2) & (icmp_ln185_reg_1059 == 1'd1) & (1'b0 == ap_block_state2_io))) begin
        mem_ARADDR = p_cast_cast_fu_655_p1;
    end else if (((1'b1 == ap_CS_fsm_state45) | ((icmp_ln188_reg_1095 == 1'd1) & (1'b1 == ap_CS_fsm_state46)))) begin
        mem_ARADDR = grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_ARADDR;
    end else if (((1'b1 == ap_CS_fsm_state37) | (1'b1 == ap_CS_fsm_state36))) begin
        mem_ARADDR = grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_ARADDR;
    end else if (((1'b1 == ap_CS_fsm_state27) | ((1'b1 == ap_CS_fsm_state28) & (icmp_ln185_reg_1059 == 1'd1)))) begin
        mem_ARADDR = grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_ARADDR;
    end else if (((1'b1 == ap_CS_fsm_state19) | (1'b1 == ap_CS_fsm_state18))) begin
        mem_ARADDR = grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_ARADDR;
    end else if (((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state9))) begin
        mem_ARADDR = grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_ARADDR;
    end else begin
        mem_ARADDR = 'bx;
    end
end

always @ (*) begin
    if ((((1'b1 == ap_CS_fsm_state38) & (mem_ARREADY == 1'b1)) | ((1'b1 == ap_CS_fsm_state29) & (mem_ARREADY == 1'b1)))) begin
        mem_ARLEN = k_assign_load_reg_1063;
    end else if ((((1'b1 == ap_CS_fsm_state20) & (mem_ARREADY == 1'b1)) | ((1'b1 == ap_CS_fsm_state11) & (mem_ARREADY == 1'b1)) | ((1'b1 == ap_CS_fsm_state2) & (icmp_ln185_reg_1059 == 1'd1) & (1'b0 == ap_block_state2_io)))) begin
        mem_ARLEN = n_assign_load_reg_1041;
    end else if (((1'b1 == ap_CS_fsm_state45) | ((icmp_ln188_reg_1095 == 1'd1) & (1'b1 == ap_CS_fsm_state46)))) begin
        mem_ARLEN = grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_ARLEN;
    end else if (((1'b1 == ap_CS_fsm_state37) | (1'b1 == ap_CS_fsm_state36))) begin
        mem_ARLEN = grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_ARLEN;
    end else if (((1'b1 == ap_CS_fsm_state27) | ((1'b1 == ap_CS_fsm_state28) & (icmp_ln185_reg_1059 == 1'd1)))) begin
        mem_ARLEN = grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_ARLEN;
    end else if (((1'b1 == ap_CS_fsm_state19) | (1'b1 == ap_CS_fsm_state18))) begin
        mem_ARLEN = grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_ARLEN;
    end else if (((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state9))) begin
        mem_ARLEN = grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_ARLEN;
    end else begin
        mem_ARLEN = 'bx;
    end
end

always @ (*) begin
    if ((((1'b1 == ap_CS_fsm_state38) & (mem_ARREADY == 1'b1)) | ((1'b1 == ap_CS_fsm_state29) & (mem_ARREADY == 1'b1)) | ((1'b1 == ap_CS_fsm_state20) & (mem_ARREADY == 1'b1)) | ((1'b1 == ap_CS_fsm_state11) & (mem_ARREADY == 1'b1)) | ((1'b1 == ap_CS_fsm_state2) & (icmp_ln185_reg_1059 == 1'd1) & (1'b0 == ap_block_state2_io)))) begin
        mem_ARVALID = 1'b1;
    end else if (((1'b1 == ap_CS_fsm_state45) | ((icmp_ln188_reg_1095 == 1'd1) & (1'b1 == ap_CS_fsm_state46)))) begin
        mem_ARVALID = grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_ARVALID;
    end else if (((1'b1 == ap_CS_fsm_state37) | (1'b1 == ap_CS_fsm_state36))) begin
        mem_ARVALID = grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_ARVALID;
    end else if (((1'b1 == ap_CS_fsm_state27) | ((1'b1 == ap_CS_fsm_state28) & (icmp_ln185_reg_1059 == 1'd1)))) begin
        mem_ARVALID = grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_ARVALID;
    end else if (((1'b1 == ap_CS_fsm_state19) | (1'b1 == ap_CS_fsm_state18))) begin
        mem_ARVALID = grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_ARVALID;
    end else if (((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state9))) begin
        mem_ARVALID = grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_ARVALID;
    end else begin
        mem_ARVALID = 1'b0;
    end
end

always @ (*) begin
    if ((~((mem_BVALID == 1'b0) | (mem_AWREADY == 1'b0)) & (1'b1 == ap_CS_fsm_state100))) begin
        mem_AWADDR = p_cast12_cast_fu_958_p1;
    end else if ((~((1'b1 == ap_block_state93_io) | ((ap_predicate_op380_writeresp_state93 == 1'b1) & (mem_BVALID == 1'b0))) & (1'b1 == ap_CS_fsm_state93) & (ap_predicate_op390_writereq_state93 == 1'b1))) begin
        mem_AWADDR = p_cast7_cast_fu_947_p1;
    end else if ((~((1'b1 == ap_block_state86_io) | ((ap_predicate_op363_writeresp_state86 == 1'b1) & (mem_BVALID == 1'b0))) & (1'b1 == ap_CS_fsm_state86) & (ap_predicate_op373_writereq_state86 == 1'b1))) begin
        mem_AWADDR = p_cast6_cast_fu_932_p1;
    end else if ((~((mem_BVALID == 1'b0) | (mem_AWREADY == 1'b0)) & (1'b1 == ap_CS_fsm_state79))) begin
        mem_AWADDR = p_cast8_cast_fu_921_p1;
    end else if (((1'b1 == ap_CS_fsm_state72) & (mem_AWREADY == 1'b1))) begin
        mem_AWADDR = p_cast5_cast_fu_910_p1;
    end else if ((~((mem_BVALID == 1'b0) | (mem_AWREADY == 1'b0)) & (1'b1 == ap_CS_fsm_state64))) begin
        mem_AWADDR = p_cast13_cast_fu_881_p1;
    end else if (((1'b1 == ap_CS_fsm_state57) & (mem_AWREADY == 1'b1))) begin
        mem_AWADDR = p_cast11_cast_fu_871_p1;
    end else if (((1'b1 == ap_CS_fsm_state49) & (mem_AWREADY == 1'b1))) begin
        mem_AWADDR = p_cast9_cast_fu_816_p1;
    end else if (((1'b1 == ap_CS_fsm_state102) | (1'b1 == ap_CS_fsm_state101))) begin
        mem_AWADDR = grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_AWADDR;
    end else if (((1'b1 == ap_CS_fsm_state95) | (1'b1 == ap_CS_fsm_state94))) begin
        mem_AWADDR = grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_AWADDR;
    end else if (((1'b1 == ap_CS_fsm_state88) | (1'b1 == ap_CS_fsm_state87))) begin
        mem_AWADDR = grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_AWADDR;
    end else if (((1'b1 == ap_CS_fsm_state81) | (1'b1 == ap_CS_fsm_state80))) begin
        mem_AWADDR = grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_AWADDR;
    end else if (((1'b1 == ap_CS_fsm_state74) | (1'b1 == ap_CS_fsm_state73))) begin
        mem_AWADDR = grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_AWADDR;
    end else if (((1'b1 == ap_CS_fsm_state66) | (1'b1 == ap_CS_fsm_state65))) begin
        mem_AWADDR = grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_AWADDR;
    end else if (((1'b1 == ap_CS_fsm_state59) | (1'b1 == ap_CS_fsm_state58))) begin
        mem_AWADDR = grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_AWADDR;
    end else if (((1'b1 == ap_CS_fsm_state51) | (1'b1 == ap_CS_fsm_state50))) begin
        mem_AWADDR = grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_AWADDR;
    end else begin
        mem_AWADDR = 'bx;
    end
end

always @ (*) begin
    if ((((1'b1 == ap_CS_fsm_state57) & (mem_AWREADY == 1'b1)) | (~((1'b1 == ap_block_state93_io) | ((ap_predicate_op380_writeresp_state93 == 1'b1) & (mem_BVALID == 1'b0))) & (1'b1 == ap_CS_fsm_state93) & (ap_predicate_op390_writereq_state93 == 1'b1)) | (~((mem_BVALID == 1'b0) | (mem_AWREADY == 1'b0)) & (1'b1 == ap_CS_fsm_state100)) | (~((mem_BVALID == 1'b0) | (mem_AWREADY == 1'b0)) & (1'b1 == ap_CS_fsm_state64)))) begin
        mem_AWLEN = k_assign_load_reg_1063;
    end else if ((((1'b1 == ap_CS_fsm_state72) & (mem_AWREADY == 1'b1)) | ((1'b1 == ap_CS_fsm_state49) & (mem_AWREADY == 1'b1)) | (~((1'b1 == ap_block_state86_io) | ((ap_predicate_op363_writeresp_state86 == 1'b1) & (mem_BVALID == 1'b0))) & (1'b1 == ap_CS_fsm_state86) & (ap_predicate_op373_writereq_state86 == 1'b1)) | (~((mem_BVALID == 1'b0) | (mem_AWREADY == 1'b0)) & (1'b1 == ap_CS_fsm_state79)))) begin
        mem_AWLEN = n_assign_load_reg_1041;
    end else if (((1'b1 == ap_CS_fsm_state102) | (1'b1 == ap_CS_fsm_state101))) begin
        mem_AWLEN = grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_AWLEN;
    end else if (((1'b1 == ap_CS_fsm_state95) | (1'b1 == ap_CS_fsm_state94))) begin
        mem_AWLEN = grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_AWLEN;
    end else if (((1'b1 == ap_CS_fsm_state88) | (1'b1 == ap_CS_fsm_state87))) begin
        mem_AWLEN = grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_AWLEN;
    end else if (((1'b1 == ap_CS_fsm_state81) | (1'b1 == ap_CS_fsm_state80))) begin
        mem_AWLEN = grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_AWLEN;
    end else if (((1'b1 == ap_CS_fsm_state74) | (1'b1 == ap_CS_fsm_state73))) begin
        mem_AWLEN = grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_AWLEN;
    end else if (((1'b1 == ap_CS_fsm_state66) | (1'b1 == ap_CS_fsm_state65))) begin
        mem_AWLEN = grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_AWLEN;
    end else if (((1'b1 == ap_CS_fsm_state59) | (1'b1 == ap_CS_fsm_state58))) begin
        mem_AWLEN = grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_AWLEN;
    end else if (((1'b1 == ap_CS_fsm_state51) | (1'b1 == ap_CS_fsm_state50))) begin
        mem_AWLEN = grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_AWLEN;
    end else begin
        mem_AWLEN = 'bx;
    end
end

always @ (*) begin
    if ((((1'b1 == ap_CS_fsm_state72) & (mem_AWREADY == 1'b1)) | ((1'b1 == ap_CS_fsm_state57) & (mem_AWREADY == 1'b1)) | ((1'b1 == ap_CS_fsm_state49) & (mem_AWREADY == 1'b1)) | (~((1'b1 == ap_block_state93_io) | ((ap_predicate_op380_writeresp_state93 == 1'b1) & (mem_BVALID == 1'b0))) & (1'b1 == ap_CS_fsm_state93) & (ap_predicate_op390_writereq_state93 == 1'b1)) | (~((1'b1 == ap_block_state86_io) | ((ap_predicate_op363_writeresp_state86 == 1'b1) & (mem_BVALID == 1'b0))) & (1'b1 == ap_CS_fsm_state86) & (ap_predicate_op373_writereq_state86 == 1'b1)) | (~((mem_BVALID == 1'b0) | (mem_AWREADY == 1'b0)) & (1'b1 == ap_CS_fsm_state100)) | (~((mem_BVALID == 1'b0) | (mem_AWREADY == 1'b0)) & (1'b1 == ap_CS_fsm_state79)) | (~((mem_BVALID == 1'b0) | (mem_AWREADY == 1'b0)) & (1'b1 == ap_CS_fsm_state64)))) begin
        mem_AWVALID = 1'b1;
    end else if (((1'b1 == ap_CS_fsm_state102) | (1'b1 == ap_CS_fsm_state101))) begin
        mem_AWVALID = grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_AWVALID;
    end else if (((1'b1 == ap_CS_fsm_state95) | (1'b1 == ap_CS_fsm_state94))) begin
        mem_AWVALID = grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_AWVALID;
    end else if (((1'b1 == ap_CS_fsm_state88) | (1'b1 == ap_CS_fsm_state87))) begin
        mem_AWVALID = grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_AWVALID;
    end else if (((1'b1 == ap_CS_fsm_state81) | (1'b1 == ap_CS_fsm_state80))) begin
        mem_AWVALID = grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_AWVALID;
    end else if (((1'b1 == ap_CS_fsm_state74) | (1'b1 == ap_CS_fsm_state73))) begin
        mem_AWVALID = grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_AWVALID;
    end else if (((1'b1 == ap_CS_fsm_state66) | (1'b1 == ap_CS_fsm_state65))) begin
        mem_AWVALID = grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_AWVALID;
    end else if (((1'b1 == ap_CS_fsm_state59) | (1'b1 == ap_CS_fsm_state58))) begin
        mem_AWVALID = grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_AWVALID;
    end else if (((1'b1 == ap_CS_fsm_state51) | (1'b1 == ap_CS_fsm_state50))) begin
        mem_AWVALID = grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_AWVALID;
    end else begin
        mem_AWVALID = 1'b0;
    end
end

always @ (*) begin
    if (((~((ap_predicate_op408_writeresp_state107 == 1'b1) & (mem_BVALID == 1'b0)) & (1'b1 == ap_CS_fsm_state107) & (ap_predicate_op408_writeresp_state107 == 1'b1)) | (~((1'b1 == ap_block_state93_io) | ((ap_predicate_op380_writeresp_state93 == 1'b1) & (mem_BVALID == 1'b0))) & (1'b1 == ap_CS_fsm_state93) & (ap_predicate_op380_writeresp_state93 == 1'b1)) | (~((1'b1 == ap_block_state86_io) | ((ap_predicate_op363_writeresp_state86 == 1'b1) & (mem_BVALID == 1'b0))) & (1'b1 == ap_CS_fsm_state86) & (ap_predicate_op363_writeresp_state86 == 1'b1)) | (~((mem_BVALID == 1'b0) | (mem_AWREADY == 1'b0)) & (1'b1 == ap_CS_fsm_state100)) | (~((mem_BVALID == 1'b0) | (mem_AWREADY == 1'b0)) & (1'b1 == ap_CS_fsm_state79)) | (~((mem_BVALID == 1'b0) | (mem_AWREADY == 1'b0)) & (1'b1 == ap_CS_fsm_state64)) | (~((ap_predicate_op298_writeresp_state56 == 1'b1) & (mem_BVALID == 1'b0)) & (1'b1 == ap_CS_fsm_state56) & (ap_predicate_op298_writeresp_state56 == 1'b1)) | (~((ap_predicate_op334_writeresp_state71 == 1'b1) & (mem_BVALID == 1'b0)) & (1'b1 == ap_CS_fsm_state71) & (ap_predicate_op334_writeresp_state71 == 1'b1)))) begin
        mem_BREADY = 1'b1;
    end else if (((1'b1 == ap_CS_fsm_state102) | (1'b1 == ap_CS_fsm_state101))) begin
        mem_BREADY = grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_BREADY;
    end else if (((1'b1 == ap_CS_fsm_state95) | (1'b1 == ap_CS_fsm_state94))) begin
        mem_BREADY = grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_BREADY;
    end else if (((1'b1 == ap_CS_fsm_state88) | (1'b1 == ap_CS_fsm_state87))) begin
        mem_BREADY = grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_BREADY;
    end else if (((1'b1 == ap_CS_fsm_state81) | (1'b1 == ap_CS_fsm_state80))) begin
        mem_BREADY = grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_BREADY;
    end else if (((1'b1 == ap_CS_fsm_state74) | (1'b1 == ap_CS_fsm_state73))) begin
        mem_BREADY = grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_BREADY;
    end else if (((1'b1 == ap_CS_fsm_state66) | (1'b1 == ap_CS_fsm_state65))) begin
        mem_BREADY = grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_BREADY;
    end else if (((1'b1 == ap_CS_fsm_state59) | (1'b1 == ap_CS_fsm_state58))) begin
        mem_BREADY = grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_BREADY;
    end else if (((1'b1 == ap_CS_fsm_state51) | (1'b1 == ap_CS_fsm_state50))) begin
        mem_BREADY = grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_BREADY;
    end else begin
        mem_BREADY = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state45) | ((icmp_ln188_reg_1095 == 1'd1) & (1'b1 == ap_CS_fsm_state46)))) begin
        mem_RREADY = grp_kmeans_top_Pipeline_5_fu_417_m_axi_mem_RREADY;
    end else if (((1'b1 == ap_CS_fsm_state37) | (1'b1 == ap_CS_fsm_state36))) begin
        mem_RREADY = grp_kmeans_top_Pipeline_4_fu_408_m_axi_mem_RREADY;
    end else if (((1'b1 == ap_CS_fsm_state27) | ((1'b1 == ap_CS_fsm_state28) & (icmp_ln185_reg_1059 == 1'd1)))) begin
        mem_RREADY = grp_kmeans_top_Pipeline_3_fu_399_m_axi_mem_RREADY;
    end else if (((1'b1 == ap_CS_fsm_state19) | (1'b1 == ap_CS_fsm_state18))) begin
        mem_RREADY = grp_kmeans_top_Pipeline_2_fu_390_m_axi_mem_RREADY;
    end else if (((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state9))) begin
        mem_RREADY = grp_kmeans_top_Pipeline_1_fu_381_m_axi_mem_RREADY;
    end else begin
        mem_RREADY = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state102) | (1'b1 == ap_CS_fsm_state101))) begin
        mem_WDATA = grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_WDATA;
    end else if (((1'b1 == ap_CS_fsm_state95) | (1'b1 == ap_CS_fsm_state94))) begin
        mem_WDATA = grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_WDATA;
    end else if (((1'b1 == ap_CS_fsm_state88) | (1'b1 == ap_CS_fsm_state87))) begin
        mem_WDATA = grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_WDATA;
    end else if (((1'b1 == ap_CS_fsm_state81) | (1'b1 == ap_CS_fsm_state80))) begin
        mem_WDATA = grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_WDATA;
    end else if (((1'b1 == ap_CS_fsm_state74) | (1'b1 == ap_CS_fsm_state73))) begin
        mem_WDATA = grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_WDATA;
    end else if (((1'b1 == ap_CS_fsm_state66) | (1'b1 == ap_CS_fsm_state65))) begin
        mem_WDATA = grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_WDATA;
    end else if (((1'b1 == ap_CS_fsm_state59) | (1'b1 == ap_CS_fsm_state58))) begin
        mem_WDATA = grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_WDATA;
    end else if (((1'b1 == ap_CS_fsm_state51) | (1'b1 == ap_CS_fsm_state50))) begin
        mem_WDATA = grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_WDATA;
    end else begin
        mem_WDATA = 'bx;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state102) | (1'b1 == ap_CS_fsm_state101))) begin
        mem_WSTRB = grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_WSTRB;
    end else if (((1'b1 == ap_CS_fsm_state95) | (1'b1 == ap_CS_fsm_state94))) begin
        mem_WSTRB = grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_WSTRB;
    end else if (((1'b1 == ap_CS_fsm_state88) | (1'b1 == ap_CS_fsm_state87))) begin
        mem_WSTRB = grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_WSTRB;
    end else if (((1'b1 == ap_CS_fsm_state81) | (1'b1 == ap_CS_fsm_state80))) begin
        mem_WSTRB = grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_WSTRB;
    end else if (((1'b1 == ap_CS_fsm_state74) | (1'b1 == ap_CS_fsm_state73))) begin
        mem_WSTRB = grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_WSTRB;
    end else if (((1'b1 == ap_CS_fsm_state66) | (1'b1 == ap_CS_fsm_state65))) begin
        mem_WSTRB = grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_WSTRB;
    end else if (((1'b1 == ap_CS_fsm_state59) | (1'b1 == ap_CS_fsm_state58))) begin
        mem_WSTRB = grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_WSTRB;
    end else if (((1'b1 == ap_CS_fsm_state51) | (1'b1 == ap_CS_fsm_state50))) begin
        mem_WSTRB = grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_WSTRB;
    end else begin
        mem_WSTRB = 'bx;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state102) | (1'b1 == ap_CS_fsm_state101))) begin
        mem_WVALID = grp_kmeans_top_Pipeline_13_fu_501_m_axi_mem_WVALID;
    end else if (((1'b1 == ap_CS_fsm_state95) | (1'b1 == ap_CS_fsm_state94))) begin
        mem_WVALID = grp_kmeans_top_Pipeline_12_fu_492_m_axi_mem_WVALID;
    end else if (((1'b1 == ap_CS_fsm_state88) | (1'b1 == ap_CS_fsm_state87))) begin
        mem_WVALID = grp_kmeans_top_Pipeline_11_fu_483_m_axi_mem_WVALID;
    end else if (((1'b1 == ap_CS_fsm_state81) | (1'b1 == ap_CS_fsm_state80))) begin
        mem_WVALID = grp_kmeans_top_Pipeline_10_fu_474_m_axi_mem_WVALID;
    end else if (((1'b1 == ap_CS_fsm_state74) | (1'b1 == ap_CS_fsm_state73))) begin
        mem_WVALID = grp_kmeans_top_Pipeline_9_fu_465_m_axi_mem_WVALID;
    end else if (((1'b1 == ap_CS_fsm_state66) | (1'b1 == ap_CS_fsm_state65))) begin
        mem_WVALID = grp_kmeans_top_Pipeline_8_fu_456_m_axi_mem_WVALID;
    end else if (((1'b1 == ap_CS_fsm_state59) | (1'b1 == ap_CS_fsm_state58))) begin
        mem_WVALID = grp_kmeans_top_Pipeline_7_fu_447_m_axi_mem_WVALID;
    end else if (((1'b1 == ap_CS_fsm_state51) | (1'b1 == ap_CS_fsm_state50))) begin
        mem_WVALID = grp_kmeans_top_Pipeline_6_fu_438_m_axi_mem_WVALID;
    end else begin
        mem_WVALID = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state38) | (1'b1 == ap_CS_fsm_state29) | (1'b1 == ap_CS_fsm_state20) | (1'b1 == ap_CS_fsm_state11) | ((1'b1 == ap_CS_fsm_state2) & (icmp_ln185_reg_1059 == 1'd1)))) begin
        mem_blk_n_AR = m_axi_mem_ARREADY;
    end else begin
        mem_blk_n_AR = 1'b1;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state100) | (1'b1 == ap_CS_fsm_state79) | (1'b1 == ap_CS_fsm_state72) | (1'b1 == ap_CS_fsm_state64) | (1'b1 == ap_CS_fsm_state57) | (1'b1 == ap_CS_fsm_state49) | ((trunc_ln215_fu_943_p1 == 1'd1) & (icmp_ln188_reg_1095 == 1'd1) & (1'b1 == ap_CS_fsm_state93)) | ((grp_fu_576_p3 == 1'd1) & (1'b1 == ap_CS_fsm_state86) & (icmp_ln185_reg_1059 == 1'd1)))) begin
        mem_blk_n_AW = m_axi_mem_AWREADY;
    end else begin
        mem_blk_n_AW = 1'b1;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state100) | (1'b1 == ap_CS_fsm_state79) | (1'b1 == ap_CS_fsm_state64) | ((trunc_ln215_reg_1229 == 1'd1) & (icmp_ln188_reg_1095 == 1'd1) & (1'b1 == ap_CS_fsm_state107)) | ((tmp_4_reg_1220 == 1'd1) & (1'b1 == ap_CS_fsm_state93) & (icmp_ln185_reg_1059 == 1'd1)) | ((tmp_3_reg_1152 == 1'd1) & (1'b1 == ap_CS_fsm_state86) & (icmp_ln185_reg_1059 == 1'd1)) | ((icmp_ln199_reg_1184 == 1'd1) & (trunc_ln199_reg_1180 == 1'd1) & (icmp_ln188_reg_1095 == 1'd1) & (1'b1 == ap_CS_fsm_state71)) | ((icmp_ln196_reg_1165 == 1'd1) & (tmp_reg_1161 == 1'd1) & (1'b1 == ap_CS_fsm_state56) & (icmp_ln185_reg_1059 == 1'd1)))) begin
        mem_blk_n_B = m_axi_mem_BVALID;
    end else begin
        mem_blk_n_B = 1'b1;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state88)) begin
        node_cluster_assignments_address0 = grp_kmeans_top_Pipeline_11_fu_483_node_cluster_assignments_address0;
    end else if ((1'b1 == ap_CS_fsm_state51)) begin
        node_cluster_assignments_address0 = grp_kmeans_top_Pipeline_6_fu_438_node_cluster_assignments_address0;
    end else begin
        node_cluster_assignments_address0 = 'bx;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state48)) begin
        node_cluster_assignments_address1 = grp_kmeans_fu_426_node_cluster_assignments_address1;
    end else if (((1'b1 == ap_CS_fsm_state28) & (icmp_ln185_reg_1059 == 1'd1))) begin
        node_cluster_assignments_address1 = grp_kmeans_top_Pipeline_3_fu_399_node_cluster_assignments_address1;
    end else begin
        node_cluster_assignments_address1 = 'bx;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state88)) begin
        node_cluster_assignments_ce0 = grp_kmeans_top_Pipeline_11_fu_483_node_cluster_assignments_ce0;
    end else if ((1'b1 == ap_CS_fsm_state51)) begin
        node_cluster_assignments_ce0 = grp_kmeans_top_Pipeline_6_fu_438_node_cluster_assignments_ce0;
    end else begin
        node_cluster_assignments_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state48)) begin
        node_cluster_assignments_ce1 = grp_kmeans_fu_426_node_cluster_assignments_ce1;
    end else if (((1'b1 == ap_CS_fsm_state28) & (icmp_ln185_reg_1059 == 1'd1))) begin
        node_cluster_assignments_ce1 = grp_kmeans_top_Pipeline_3_fu_399_node_cluster_assignments_ce1;
    end else begin
        node_cluster_assignments_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state48)) begin
        node_cluster_assignments_d1 = grp_kmeans_fu_426_node_cluster_assignments_d1;
    end else if (((1'b1 == ap_CS_fsm_state28) & (icmp_ln185_reg_1059 == 1'd1))) begin
        node_cluster_assignments_d1 = grp_kmeans_top_Pipeline_3_fu_399_node_cluster_assignments_d1;
    end else begin
        node_cluster_assignments_d1 = 'bx;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state48)) begin
        node_cluster_assignments_we1 = grp_kmeans_fu_426_node_cluster_assignments_we1;
    end else if (((1'b1 == ap_CS_fsm_state28) & (icmp_ln185_reg_1059 == 1'd1))) begin
        node_cluster_assignments_we1 = grp_kmeans_top_Pipeline_3_fu_399_node_cluster_assignments_we1;
    end else begin
        node_cluster_assignments_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state74)) begin
        node_x_coords_address0 = grp_kmeans_top_Pipeline_9_fu_465_node_x_coords_address0;
    end else if ((1'b1 == ap_CS_fsm_state48)) begin
        node_x_coords_address0 = grp_kmeans_fu_426_node_x_coords_address0;
    end else begin
        node_x_coords_address0 = 'bx;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state48)) begin
        node_x_coords_address1 = grp_kmeans_fu_426_node_x_coords_address1;
    end else if ((1'b1 == ap_CS_fsm_state10)) begin
        node_x_coords_address1 = grp_kmeans_top_Pipeline_1_fu_381_node_x_coords_address1;
    end else begin
        node_x_coords_address1 = 'bx;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state74)) begin
        node_x_coords_ce0 = grp_kmeans_top_Pipeline_9_fu_465_node_x_coords_ce0;
    end else if ((1'b1 == ap_CS_fsm_state48)) begin
        node_x_coords_ce0 = grp_kmeans_fu_426_node_x_coords_ce0;
    end else begin
        node_x_coords_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state48)) begin
        node_x_coords_ce1 = grp_kmeans_fu_426_node_x_coords_ce1;
    end else if ((1'b1 == ap_CS_fsm_state10)) begin
        node_x_coords_ce1 = grp_kmeans_top_Pipeline_1_fu_381_node_x_coords_ce1;
    end else begin
        node_x_coords_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state10)) begin
        node_x_coords_we1 = grp_kmeans_top_Pipeline_1_fu_381_node_x_coords_we1;
    end else begin
        node_x_coords_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state81)) begin
        node_y_coords_address0 = grp_kmeans_top_Pipeline_10_fu_474_node_y_coords_address0;
    end else if ((1'b1 == ap_CS_fsm_state48)) begin
        node_y_coords_address0 = grp_kmeans_fu_426_node_y_coords_address0;
    end else begin
        node_y_coords_address0 = 'bx;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state48)) begin
        node_y_coords_address1 = grp_kmeans_fu_426_node_y_coords_address1;
    end else if ((1'b1 == ap_CS_fsm_state19)) begin
        node_y_coords_address1 = grp_kmeans_top_Pipeline_2_fu_390_node_y_coords_address1;
    end else begin
        node_y_coords_address1 = 'bx;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state81)) begin
        node_y_coords_ce0 = grp_kmeans_top_Pipeline_10_fu_474_node_y_coords_ce0;
    end else if ((1'b1 == ap_CS_fsm_state48)) begin
        node_y_coords_ce0 = grp_kmeans_fu_426_node_y_coords_ce0;
    end else begin
        node_y_coords_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state48)) begin
        node_y_coords_ce1 = grp_kmeans_fu_426_node_y_coords_ce1;
    end else if ((1'b1 == ap_CS_fsm_state19)) begin
        node_y_coords_ce1 = grp_kmeans_top_Pipeline_2_fu_390_node_y_coords_ce1;
    end else begin
        node_y_coords_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state19)) begin
        node_y_coords_we1 = grp_kmeans_top_Pipeline_2_fu_390_node_y_coords_we1;
    end else begin
        node_y_coords_we1 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            if (((1'b1 == ap_CS_fsm_state2) & (icmp_ln185_reg_1059 == 1'd0) & (1'b0 == ap_block_state2_io))) begin
                ap_NS_fsm = ap_ST_fsm_state28;
            end else if (((1'b1 == ap_CS_fsm_state2) & (icmp_ln185_reg_1059 == 1'd1) & (1'b0 == ap_block_state2_io))) begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end
        end
        ap_ST_fsm_state3 : begin
            ap_NS_fsm = ap_ST_fsm_state4;
        end
        ap_ST_fsm_state4 : begin
            ap_NS_fsm = ap_ST_fsm_state5;
        end
        ap_ST_fsm_state5 : begin
            ap_NS_fsm = ap_ST_fsm_state6;
        end
        ap_ST_fsm_state6 : begin
            ap_NS_fsm = ap_ST_fsm_state7;
        end
        ap_ST_fsm_state7 : begin
            ap_NS_fsm = ap_ST_fsm_state8;
        end
        ap_ST_fsm_state8 : begin
            ap_NS_fsm = ap_ST_fsm_state9;
        end
        ap_ST_fsm_state9 : begin
            ap_NS_fsm = ap_ST_fsm_state10;
        end
        ap_ST_fsm_state10 : begin
            if (((grp_kmeans_top_Pipeline_1_fu_381_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state10))) begin
                ap_NS_fsm = ap_ST_fsm_state11;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state10;
            end
        end
        ap_ST_fsm_state11 : begin
            if (((1'b1 == ap_CS_fsm_state11) & (mem_ARREADY == 1'b1))) begin
                ap_NS_fsm = ap_ST_fsm_state12;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state11;
            end
        end
        ap_ST_fsm_state12 : begin
            ap_NS_fsm = ap_ST_fsm_state13;
        end
        ap_ST_fsm_state13 : begin
            ap_NS_fsm = ap_ST_fsm_state14;
        end
        ap_ST_fsm_state14 : begin
            ap_NS_fsm = ap_ST_fsm_state15;
        end
        ap_ST_fsm_state15 : begin
            ap_NS_fsm = ap_ST_fsm_state16;
        end
        ap_ST_fsm_state16 : begin
            ap_NS_fsm = ap_ST_fsm_state17;
        end
        ap_ST_fsm_state17 : begin
            ap_NS_fsm = ap_ST_fsm_state18;
        end
        ap_ST_fsm_state18 : begin
            ap_NS_fsm = ap_ST_fsm_state19;
        end
        ap_ST_fsm_state19 : begin
            if (((grp_kmeans_top_Pipeline_2_fu_390_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state19))) begin
                ap_NS_fsm = ap_ST_fsm_state20;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state19;
            end
        end
        ap_ST_fsm_state20 : begin
            if (((1'b1 == ap_CS_fsm_state20) & (mem_ARREADY == 1'b1))) begin
                ap_NS_fsm = ap_ST_fsm_state21;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state20;
            end
        end
        ap_ST_fsm_state21 : begin
            ap_NS_fsm = ap_ST_fsm_state22;
        end
        ap_ST_fsm_state22 : begin
            ap_NS_fsm = ap_ST_fsm_state23;
        end
        ap_ST_fsm_state23 : begin
            ap_NS_fsm = ap_ST_fsm_state24;
        end
        ap_ST_fsm_state24 : begin
            ap_NS_fsm = ap_ST_fsm_state25;
        end
        ap_ST_fsm_state25 : begin
            ap_NS_fsm = ap_ST_fsm_state26;
        end
        ap_ST_fsm_state26 : begin
            ap_NS_fsm = ap_ST_fsm_state27;
        end
        ap_ST_fsm_state27 : begin
            ap_NS_fsm = ap_ST_fsm_state28;
        end
        ap_ST_fsm_state28 : begin
            if (((icmp_ln188_fu_688_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state28) & (1'b0 == ap_block_state28_on_subcall_done))) begin
                ap_NS_fsm = ap_ST_fsm_state46;
            end else if (((icmp_ln188_fu_688_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state28) & (1'b0 == ap_block_state28_on_subcall_done))) begin
                ap_NS_fsm = ap_ST_fsm_state29;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state28;
            end
        end
        ap_ST_fsm_state29 : begin
            if (((1'b1 == ap_CS_fsm_state29) & (mem_ARREADY == 1'b1))) begin
                ap_NS_fsm = ap_ST_fsm_state30;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state29;
            end
        end
        ap_ST_fsm_state30 : begin
            ap_NS_fsm = ap_ST_fsm_state31;
        end
        ap_ST_fsm_state31 : begin
            ap_NS_fsm = ap_ST_fsm_state32;
        end
        ap_ST_fsm_state32 : begin
            ap_NS_fsm = ap_ST_fsm_state33;
        end
        ap_ST_fsm_state33 : begin
            ap_NS_fsm = ap_ST_fsm_state34;
        end
        ap_ST_fsm_state34 : begin
            ap_NS_fsm = ap_ST_fsm_state35;
        end
        ap_ST_fsm_state35 : begin
            ap_NS_fsm = ap_ST_fsm_state36;
        end
        ap_ST_fsm_state36 : begin
            ap_NS_fsm = ap_ST_fsm_state37;
        end
        ap_ST_fsm_state37 : begin
            if (((grp_kmeans_top_Pipeline_4_fu_408_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state37))) begin
                ap_NS_fsm = ap_ST_fsm_state38;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state37;
            end
        end
        ap_ST_fsm_state38 : begin
            if (((1'b1 == ap_CS_fsm_state38) & (mem_ARREADY == 1'b1))) begin
                ap_NS_fsm = ap_ST_fsm_state39;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state38;
            end
        end
        ap_ST_fsm_state39 : begin
            ap_NS_fsm = ap_ST_fsm_state40;
        end
        ap_ST_fsm_state40 : begin
            ap_NS_fsm = ap_ST_fsm_state41;
        end
        ap_ST_fsm_state41 : begin
            ap_NS_fsm = ap_ST_fsm_state42;
        end
        ap_ST_fsm_state42 : begin
            ap_NS_fsm = ap_ST_fsm_state43;
        end
        ap_ST_fsm_state43 : begin
            ap_NS_fsm = ap_ST_fsm_state44;
        end
        ap_ST_fsm_state44 : begin
            ap_NS_fsm = ap_ST_fsm_state45;
        end
        ap_ST_fsm_state45 : begin
            ap_NS_fsm = ap_ST_fsm_state46;
        end
        ap_ST_fsm_state46 : begin
            if (((1'b1 == ap_CS_fsm_state46) & (1'b0 == ap_block_state46_on_subcall_done))) begin
                ap_NS_fsm = ap_ST_fsm_state47;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state46;
            end
        end
        ap_ST_fsm_state47 : begin
            if (((1'b1 == ap_CS_fsm_state47) & (((ap_phi_mux_phi_ln191_phi_fu_374_p4 == 1'd1) & (tmp_3_fu_782_p3 == 1'd1) & (icmp_ln185_reg_1059 == 1'd1)) | ((tmp_3_fu_782_p3 == 1'd1) & (icmp_ln191_fu_738_p2 == 1'd0) & (icmp_ln185_reg_1059 == 1'd1))))) begin
                ap_NS_fsm = ap_ST_fsm_state72;
            end else if (((1'b1 == ap_CS_fsm_state47) & (((((ap_phi_mux_phi_ln191_phi_fu_374_p4 == 1'd1) & (tmp_3_fu_782_p3 == 1'd0)) | ((tmp_3_fu_782_p3 == 1'd0) & (icmp_ln191_fu_738_p2 == 1'd0))) | ((icmp_ln191_fu_738_p2 == 1'd0) & (icmp_ln185_reg_1059 == 1'd0))) | ((ap_phi_mux_phi_ln191_phi_fu_374_p4 == 1'd1) & (icmp_ln185_reg_1059 == 1'd0))))) begin
                ap_NS_fsm = ap_ST_fsm_state86;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state48;
            end
        end
        ap_ST_fsm_state48 : begin
            if (((grp_kmeans_fu_426_ap_done == 1'b1) & (grp_fu_584_p2 == 1'd1) & (grp_fu_576_p3 == 1'd1) & (1'b1 == ap_CS_fsm_state48) & (icmp_ln185_reg_1059 == 1'd1))) begin
                ap_NS_fsm = ap_ST_fsm_state49;
            end else if (((grp_kmeans_fu_426_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state48) & ((icmp_ln185_reg_1059 == 1'd0) | ((grp_fu_584_p2 == 1'd0) | (grp_fu_576_p3 == 1'd0))))) begin
                ap_NS_fsm = ap_ST_fsm_state56;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state48;
            end
        end
        ap_ST_fsm_state49 : begin
            if (((1'b1 == ap_CS_fsm_state49) & (mem_AWREADY == 1'b1))) begin
                ap_NS_fsm = ap_ST_fsm_state50;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state49;
            end
        end
        ap_ST_fsm_state50 : begin
            ap_NS_fsm = ap_ST_fsm_state51;
        end
        ap_ST_fsm_state51 : begin
            if (((grp_kmeans_top_Pipeline_6_fu_438_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state51))) begin
                ap_NS_fsm = ap_ST_fsm_state52;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state51;
            end
        end
        ap_ST_fsm_state52 : begin
            ap_NS_fsm = ap_ST_fsm_state53;
        end
        ap_ST_fsm_state53 : begin
            ap_NS_fsm = ap_ST_fsm_state54;
        end
        ap_ST_fsm_state54 : begin
            ap_NS_fsm = ap_ST_fsm_state55;
        end
        ap_ST_fsm_state55 : begin
            ap_NS_fsm = ap_ST_fsm_state56;
        end
        ap_ST_fsm_state56 : begin
            if ((~((ap_predicate_op298_writeresp_state56 == 1'b1) & (mem_BVALID == 1'b0)) & (trunc_ln199_fu_826_p1 == 1'd1) & (grp_fu_584_p2 == 1'd1) & (icmp_ln188_reg_1095 == 1'd1) & (1'b1 == ap_CS_fsm_state56))) begin
                ap_NS_fsm = ap_ST_fsm_state57;
            end else if ((~((ap_predicate_op298_writeresp_state56 == 1'b1) & (mem_BVALID == 1'b0)) & (1'b1 == ap_CS_fsm_state56) & ((icmp_ln188_reg_1095 == 1'd0) | ((trunc_ln199_fu_826_p1 == 1'd0) | (grp_fu_584_p2 == 1'd0))))) begin
                ap_NS_fsm = ap_ST_fsm_state71;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state56;
            end
        end
        ap_ST_fsm_state57 : begin
            if (((1'b1 == ap_CS_fsm_state57) & (mem_AWREADY == 1'b1))) begin
                ap_NS_fsm = ap_ST_fsm_state58;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state57;
            end
        end
        ap_ST_fsm_state58 : begin
            ap_NS_fsm = ap_ST_fsm_state59;
        end
        ap_ST_fsm_state59 : begin
            if (((grp_kmeans_top_Pipeline_7_fu_447_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state59))) begin
                ap_NS_fsm = ap_ST_fsm_state60;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state59;
            end
        end
        ap_ST_fsm_state60 : begin
            ap_NS_fsm = ap_ST_fsm_state61;
        end
        ap_ST_fsm_state61 : begin
            ap_NS_fsm = ap_ST_fsm_state62;
        end
        ap_ST_fsm_state62 : begin
            ap_NS_fsm = ap_ST_fsm_state63;
        end
        ap_ST_fsm_state63 : begin
            ap_NS_fsm = ap_ST_fsm_state64;
        end
        ap_ST_fsm_state64 : begin
            if ((~((mem_BVALID == 1'b0) | (mem_AWREADY == 1'b0)) & (1'b1 == ap_CS_fsm_state64))) begin
                ap_NS_fsm = ap_ST_fsm_state65;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state64;
            end
        end
        ap_ST_fsm_state65 : begin
            ap_NS_fsm = ap_ST_fsm_state66;
        end
        ap_ST_fsm_state66 : begin
            if (((grp_kmeans_top_Pipeline_8_fu_456_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state66))) begin
                ap_NS_fsm = ap_ST_fsm_state67;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state66;
            end
        end
        ap_ST_fsm_state67 : begin
            ap_NS_fsm = ap_ST_fsm_state68;
        end
        ap_ST_fsm_state68 : begin
            ap_NS_fsm = ap_ST_fsm_state69;
        end
        ap_ST_fsm_state69 : begin
            ap_NS_fsm = ap_ST_fsm_state70;
        end
        ap_ST_fsm_state70 : begin
            ap_NS_fsm = ap_ST_fsm_state71;
        end
        ap_ST_fsm_state71 : begin
            if ((~((ap_predicate_op334_writeresp_state71 == 1'b1) & (mem_BVALID == 1'b0)) & (1'b1 == ap_CS_fsm_state71))) begin
                ap_NS_fsm = ap_ST_fsm_state47;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state71;
            end
        end
        ap_ST_fsm_state72 : begin
            if (((1'b1 == ap_CS_fsm_state72) & (mem_AWREADY == 1'b1))) begin
                ap_NS_fsm = ap_ST_fsm_state73;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state72;
            end
        end
        ap_ST_fsm_state73 : begin
            ap_NS_fsm = ap_ST_fsm_state74;
        end
        ap_ST_fsm_state74 : begin
            if (((1'b1 == ap_CS_fsm_state74) & (grp_kmeans_top_Pipeline_9_fu_465_ap_done == 1'b1))) begin
                ap_NS_fsm = ap_ST_fsm_state75;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state74;
            end
        end
        ap_ST_fsm_state75 : begin
            ap_NS_fsm = ap_ST_fsm_state76;
        end
        ap_ST_fsm_state76 : begin
            ap_NS_fsm = ap_ST_fsm_state77;
        end
        ap_ST_fsm_state77 : begin
            ap_NS_fsm = ap_ST_fsm_state78;
        end
        ap_ST_fsm_state78 : begin
            ap_NS_fsm = ap_ST_fsm_state79;
        end
        ap_ST_fsm_state79 : begin
            if ((~((mem_BVALID == 1'b0) | (mem_AWREADY == 1'b0)) & (1'b1 == ap_CS_fsm_state79))) begin
                ap_NS_fsm = ap_ST_fsm_state80;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state79;
            end
        end
        ap_ST_fsm_state80 : begin
            ap_NS_fsm = ap_ST_fsm_state81;
        end
        ap_ST_fsm_state81 : begin
            if (((1'b1 == ap_CS_fsm_state81) & (grp_kmeans_top_Pipeline_10_fu_474_ap_done == 1'b1))) begin
                ap_NS_fsm = ap_ST_fsm_state82;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state81;
            end
        end
        ap_ST_fsm_state82 : begin
            ap_NS_fsm = ap_ST_fsm_state83;
        end
        ap_ST_fsm_state83 : begin
            ap_NS_fsm = ap_ST_fsm_state84;
        end
        ap_ST_fsm_state84 : begin
            ap_NS_fsm = ap_ST_fsm_state85;
        end
        ap_ST_fsm_state85 : begin
            ap_NS_fsm = ap_ST_fsm_state86;
        end
        ap_ST_fsm_state86 : begin
            if ((~((1'b1 == ap_block_state86_io) | ((ap_predicate_op363_writeresp_state86 == 1'b1) & (mem_BVALID == 1'b0))) & (grp_fu_576_p3 == 1'd1) & (1'b1 == ap_CS_fsm_state86) & (icmp_ln185_reg_1059 == 1'd1))) begin
                ap_NS_fsm = ap_ST_fsm_state87;
            end else if ((~((1'b1 == ap_block_state86_io) | ((ap_predicate_op363_writeresp_state86 == 1'b1) & (mem_BVALID == 1'b0))) & (1'b1 == ap_CS_fsm_state86) & ((grp_fu_576_p3 == 1'd0) | (icmp_ln185_reg_1059 == 1'd0)))) begin
                ap_NS_fsm = ap_ST_fsm_state93;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state86;
            end
        end
        ap_ST_fsm_state87 : begin
            ap_NS_fsm = ap_ST_fsm_state88;
        end
        ap_ST_fsm_state88 : begin
            if (((1'b1 == ap_CS_fsm_state88) & (grp_kmeans_top_Pipeline_11_fu_483_ap_done == 1'b1))) begin
                ap_NS_fsm = ap_ST_fsm_state89;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state88;
            end
        end
        ap_ST_fsm_state89 : begin
            ap_NS_fsm = ap_ST_fsm_state90;
        end
        ap_ST_fsm_state90 : begin
            ap_NS_fsm = ap_ST_fsm_state91;
        end
        ap_ST_fsm_state91 : begin
            ap_NS_fsm = ap_ST_fsm_state92;
        end
        ap_ST_fsm_state92 : begin
            ap_NS_fsm = ap_ST_fsm_state93;
        end
        ap_ST_fsm_state93 : begin
            if ((~((1'b1 == ap_block_state93_io) | ((ap_predicate_op380_writeresp_state93 == 1'b1) & (mem_BVALID == 1'b0))) & (trunc_ln215_fu_943_p1 == 1'd1) & (icmp_ln188_reg_1095 == 1'd1) & (1'b1 == ap_CS_fsm_state93))) begin
                ap_NS_fsm = ap_ST_fsm_state94;
            end else if ((~((1'b1 == ap_block_state93_io) | ((ap_predicate_op380_writeresp_state93 == 1'b1) & (mem_BVALID == 1'b0))) & (1'b1 == ap_CS_fsm_state93) & ((trunc_ln215_fu_943_p1 == 1'd0) | (icmp_ln188_reg_1095 == 1'd0)))) begin
                ap_NS_fsm = ap_ST_fsm_state107;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state93;
            end
        end
        ap_ST_fsm_state94 : begin
            ap_NS_fsm = ap_ST_fsm_state95;
        end
        ap_ST_fsm_state95 : begin
            if (((1'b1 == ap_CS_fsm_state95) & (grp_kmeans_top_Pipeline_12_fu_492_ap_done == 1'b1))) begin
                ap_NS_fsm = ap_ST_fsm_state96;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state95;
            end
        end
        ap_ST_fsm_state96 : begin
            ap_NS_fsm = ap_ST_fsm_state97;
        end
        ap_ST_fsm_state97 : begin
            ap_NS_fsm = ap_ST_fsm_state98;
        end
        ap_ST_fsm_state98 : begin
            ap_NS_fsm = ap_ST_fsm_state99;
        end
        ap_ST_fsm_state99 : begin
            ap_NS_fsm = ap_ST_fsm_state100;
        end
        ap_ST_fsm_state100 : begin
            if ((~((mem_BVALID == 1'b0) | (mem_AWREADY == 1'b0)) & (1'b1 == ap_CS_fsm_state100))) begin
                ap_NS_fsm = ap_ST_fsm_state101;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state100;
            end
        end
        ap_ST_fsm_state101 : begin
            ap_NS_fsm = ap_ST_fsm_state102;
        end
        ap_ST_fsm_state102 : begin
            if (((1'b1 == ap_CS_fsm_state102) & (grp_kmeans_top_Pipeline_13_fu_501_ap_done == 1'b1))) begin
                ap_NS_fsm = ap_ST_fsm_state103;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state102;
            end
        end
        ap_ST_fsm_state103 : begin
            ap_NS_fsm = ap_ST_fsm_state104;
        end
        ap_ST_fsm_state104 : begin
            ap_NS_fsm = ap_ST_fsm_state105;
        end
        ap_ST_fsm_state105 : begin
            ap_NS_fsm = ap_ST_fsm_state106;
        end
        ap_ST_fsm_state106 : begin
            ap_NS_fsm = ap_ST_fsm_state107;
        end
        ap_ST_fsm_state107 : begin
            if ((~((ap_predicate_op408_writeresp_state107 == 1'b1) & (mem_BVALID == 1'b0)) & (1'b1 == ap_CS_fsm_state107))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state107;
            end
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state10 = ap_CS_fsm[32'd9];

assign ap_CS_fsm_state100 = ap_CS_fsm[32'd99];

assign ap_CS_fsm_state101 = ap_CS_fsm[32'd100];

assign ap_CS_fsm_state102 = ap_CS_fsm[32'd101];

assign ap_CS_fsm_state107 = ap_CS_fsm[32'd106];

assign ap_CS_fsm_state11 = ap_CS_fsm[32'd10];

assign ap_CS_fsm_state17 = ap_CS_fsm[32'd16];

assign ap_CS_fsm_state18 = ap_CS_fsm[32'd17];

assign ap_CS_fsm_state19 = ap_CS_fsm[32'd18];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state20 = ap_CS_fsm[32'd19];

assign ap_CS_fsm_state26 = ap_CS_fsm[32'd25];

assign ap_CS_fsm_state27 = ap_CS_fsm[32'd26];

assign ap_CS_fsm_state28 = ap_CS_fsm[32'd27];

assign ap_CS_fsm_state29 = ap_CS_fsm[32'd28];

assign ap_CS_fsm_state35 = ap_CS_fsm[32'd34];

assign ap_CS_fsm_state36 = ap_CS_fsm[32'd35];

assign ap_CS_fsm_state37 = ap_CS_fsm[32'd36];

assign ap_CS_fsm_state38 = ap_CS_fsm[32'd37];

assign ap_CS_fsm_state44 = ap_CS_fsm[32'd43];

assign ap_CS_fsm_state45 = ap_CS_fsm[32'd44];

assign ap_CS_fsm_state46 = ap_CS_fsm[32'd45];

assign ap_CS_fsm_state47 = ap_CS_fsm[32'd46];

assign ap_CS_fsm_state48 = ap_CS_fsm[32'd47];

assign ap_CS_fsm_state49 = ap_CS_fsm[32'd48];

assign ap_CS_fsm_state50 = ap_CS_fsm[32'd49];

assign ap_CS_fsm_state51 = ap_CS_fsm[32'd50];

assign ap_CS_fsm_state56 = ap_CS_fsm[32'd55];

assign ap_CS_fsm_state57 = ap_CS_fsm[32'd56];

assign ap_CS_fsm_state58 = ap_CS_fsm[32'd57];

assign ap_CS_fsm_state59 = ap_CS_fsm[32'd58];

assign ap_CS_fsm_state64 = ap_CS_fsm[32'd63];

assign ap_CS_fsm_state65 = ap_CS_fsm[32'd64];

assign ap_CS_fsm_state66 = ap_CS_fsm[32'd65];

assign ap_CS_fsm_state71 = ap_CS_fsm[32'd70];

assign ap_CS_fsm_state72 = ap_CS_fsm[32'd71];

assign ap_CS_fsm_state73 = ap_CS_fsm[32'd72];

assign ap_CS_fsm_state74 = ap_CS_fsm[32'd73];

assign ap_CS_fsm_state79 = ap_CS_fsm[32'd78];

assign ap_CS_fsm_state8 = ap_CS_fsm[32'd7];

assign ap_CS_fsm_state80 = ap_CS_fsm[32'd79];

assign ap_CS_fsm_state81 = ap_CS_fsm[32'd80];

assign ap_CS_fsm_state86 = ap_CS_fsm[32'd85];

assign ap_CS_fsm_state87 = ap_CS_fsm[32'd86];

assign ap_CS_fsm_state88 = ap_CS_fsm[32'd87];

assign ap_CS_fsm_state9 = ap_CS_fsm[32'd8];

assign ap_CS_fsm_state93 = ap_CS_fsm[32'd92];

assign ap_CS_fsm_state94 = ap_CS_fsm[32'd93];

assign ap_CS_fsm_state95 = ap_CS_fsm[32'd94];

assign ap_NS_fsm_state101 = ap_NS_fsm[32'd100];

assign ap_NS_fsm_state18 = ap_NS_fsm[32'd17];

assign ap_NS_fsm_state27 = ap_NS_fsm[32'd26];

assign ap_NS_fsm_state36 = ap_NS_fsm[32'd35];

assign ap_NS_fsm_state45 = ap_NS_fsm[32'd44];

assign ap_NS_fsm_state50 = ap_NS_fsm[32'd49];

assign ap_NS_fsm_state58 = ap_NS_fsm[32'd57];

assign ap_NS_fsm_state65 = ap_NS_fsm[32'd64];

assign ap_NS_fsm_state73 = ap_NS_fsm[32'd72];

assign ap_NS_fsm_state80 = ap_NS_fsm[32'd79];

assign ap_NS_fsm_state87 = ap_NS_fsm[32'd86];

assign ap_NS_fsm_state9 = ap_NS_fsm[32'd8];

assign ap_NS_fsm_state94 = ap_NS_fsm[32'd93];

always @ (*) begin
    ap_block_state107 = ((ap_predicate_op408_writeresp_state107 == 1'b1) & (mem_BVALID == 1'b0));
end

always @ (*) begin
    ap_block_state28_on_subcall_done = ((grp_kmeans_top_Pipeline_3_fu_399_ap_done == 1'b0) & (icmp_ln185_reg_1059 == 1'd1));
end

always @ (*) begin
    ap_block_state2_io = ((icmp_ln185_reg_1059 == 1'd1) & (mem_ARREADY == 1'b0));
end

always @ (*) begin
    ap_block_state46_on_subcall_done = ((grp_kmeans_top_Pipeline_5_fu_417_ap_done == 1'b0) & (icmp_ln188_reg_1095 == 1'd1));
end

always @ (*) begin
    ap_block_state56 = ((ap_predicate_op298_writeresp_state56 == 1'b1) & (mem_BVALID == 1'b0));
end

always @ (*) begin
    ap_block_state71 = ((ap_predicate_op334_writeresp_state71 == 1'b1) & (mem_BVALID == 1'b0));
end

always @ (*) begin
    ap_block_state86 = ((ap_predicate_op363_writeresp_state86 == 1'b1) & (mem_BVALID == 1'b0));
end

always @ (*) begin
    ap_block_state86_io = ((ap_predicate_op373_writereq_state86 == 1'b1) & (mem_AWREADY == 1'b0));
end

always @ (*) begin
    ap_block_state93 = ((ap_predicate_op380_writeresp_state93 == 1'b1) & (mem_BVALID == 1'b0));
end

always @ (*) begin
    ap_block_state93_io = ((ap_predicate_op390_writereq_state93 == 1'b1) & (mem_AWREADY == 1'b0));
end

assign ap_phi_mux_phi_ln191_phi_fu_374_p4 = phi_ln191_reg_370;

always @ (*) begin
    ap_predicate_op298_writeresp_state56 = ((icmp_ln196_reg_1165 == 1'd1) & (tmp_reg_1161 == 1'd1) & (icmp_ln185_reg_1059 == 1'd1));
end

always @ (*) begin
    ap_predicate_op334_writeresp_state71 = ((icmp_ln199_reg_1184 == 1'd1) & (trunc_ln199_reg_1180 == 1'd1) & (icmp_ln188_reg_1095 == 1'd1));
end

always @ (*) begin
    ap_predicate_op363_writeresp_state86 = ((tmp_3_reg_1152 == 1'd1) & (icmp_ln185_reg_1059 == 1'd1));
end

always @ (*) begin
    ap_predicate_op373_writereq_state86 = ((grp_fu_576_p3 == 1'd1) & (icmp_ln185_reg_1059 == 1'd1));
end

always @ (*) begin
    ap_predicate_op380_writeresp_state93 = ((tmp_4_reg_1220 == 1'd1) & (icmp_ln185_reg_1059 == 1'd1));
end

always @ (*) begin
    ap_predicate_op390_writereq_state93 = ((trunc_ln215_fu_943_p1 == 1'd1) & (icmp_ln188_reg_1095 == 1'd1));
end

always @ (*) begin
    ap_predicate_op408_writeresp_state107 = ((trunc_ln215_reg_1229 == 1'd1) & (icmp_ln188_reg_1095 == 1'd1));
end

always @ (*) begin
    ap_rst_n_inv = ~ap_rst_n;
end

assign current_iteration_1_fu_895_p2 = (trunc_ln204_fu_891_p1 + current_iteration_fu_202);

assign empty_50_fu_801_p2 = (p_cast14_fu_797_p1 + buf_ptr_intermediate_cluster_assignments_read_reg_979);

assign empty_53_fu_841_p2 = (p_cast15_fu_837_p1 + buf_ptr_intermediate_centroid_x_coords_read_reg_974);

assign empty_56_fu_856_p2 = (p_cast15_fu_837_p1 + buf_ptr_intermediate_centroid_y_coords_read_reg_969);

assign grp_fu_518_p4 = {{buf_ptr_node_x_coords_read_reg_1004[63:3]}};

assign grp_fu_527_p4 = {{buf_ptr_node_y_coords_read_reg_999[63:3]}};

assign grp_fu_536_p4 = {{buf_ptr_node_cluster_assignments_read_reg_994[63:3]}};

assign grp_fu_545_p4 = {{buf_ptr_centroid_x_coords_read_reg_989[63:3]}};

assign grp_fu_554_p4 = {{buf_ptr_centroid_y_coords_read_reg_984[63:3]}};

assign grp_fu_576_p3 = control_assign_fu_166[32'd1];

assign grp_fu_584_p2 = ((sub_iterations_assign_fu_174 < max_iterations_assign_fu_170) ? 1'b1 : 1'b0);

assign grp_kmeans_fu_426_ap_start = grp_kmeans_fu_426_ap_start_reg;

assign grp_kmeans_top_Pipeline_10_fu_474_ap_start = grp_kmeans_top_Pipeline_10_fu_474_ap_start_reg;

assign grp_kmeans_top_Pipeline_11_fu_483_ap_start = grp_kmeans_top_Pipeline_11_fu_483_ap_start_reg;

assign grp_kmeans_top_Pipeline_12_fu_492_ap_start = grp_kmeans_top_Pipeline_12_fu_492_ap_start_reg;

assign grp_kmeans_top_Pipeline_13_fu_501_ap_start = grp_kmeans_top_Pipeline_13_fu_501_ap_start_reg;

assign grp_kmeans_top_Pipeline_1_fu_381_ap_start = grp_kmeans_top_Pipeline_1_fu_381_ap_start_reg;

assign grp_kmeans_top_Pipeline_2_fu_390_ap_start = grp_kmeans_top_Pipeline_2_fu_390_ap_start_reg;

assign grp_kmeans_top_Pipeline_3_fu_399_ap_start = grp_kmeans_top_Pipeline_3_fu_399_ap_start_reg;

assign grp_kmeans_top_Pipeline_4_fu_408_ap_start = grp_kmeans_top_Pipeline_4_fu_408_ap_start_reg;

assign grp_kmeans_top_Pipeline_5_fu_417_ap_start = grp_kmeans_top_Pipeline_5_fu_417_ap_start_reg;

assign grp_kmeans_top_Pipeline_6_fu_438_ap_start = grp_kmeans_top_Pipeline_6_fu_438_ap_start_reg;

assign grp_kmeans_top_Pipeline_7_fu_447_ap_start = grp_kmeans_top_Pipeline_7_fu_447_ap_start_reg;

assign grp_kmeans_top_Pipeline_8_fu_456_ap_start = grp_kmeans_top_Pipeline_8_fu_456_ap_start_reg;

assign grp_kmeans_top_Pipeline_9_fu_465_ap_start = grp_kmeans_top_Pipeline_9_fu_465_ap_start_reg;

assign icmp_ln185_fu_649_p2 = ((grp_load_fu_510_p1 != 32'd0) ? 1'b1 : 1'b0);

assign icmp_ln188_fu_688_p2 = ((k_assign_load_reg_1063 != 32'd0) ? 1'b1 : 1'b0);

assign icmp_ln191_fu_738_p2 = ((max_iterations_assign_fu_170 > sext_ln191_fu_734_p1) ? 1'b1 : 1'b0);

assign intermediate_writes_made_2_fu_728_p2 = (intermediate_writes_made_fu_198 + 32'd1);

assign mul_ln194_fu_776_p0 = intermediate_writes_made_fu_198[28:0];

assign mul_ln194_fu_776_p1 = (trunc_ln194_fu_747_p1 + shl_ln_fu_758_p3);

assign p_cast11_cast_fu_871_p1 = $signed(p_cast10_reg_1188);

assign p_cast12_cast_fu_958_p1 = $signed(reg_614);

assign p_cast13_cast_fu_881_p1 = $signed(p_cast11_reg_1194);

assign p_cast14_fu_797_p1 = tmp_1_fu_790_p3;

assign p_cast15_fu_837_p1 = tmp_2_fu_830_p3;

assign p_cast1_cast_fu_693_p1 = grp_fu_545_p4;

assign p_cast2_cast_fu_666_p1 = grp_fu_527_p4;

assign p_cast3_cast_fu_704_p1 = grp_fu_554_p4;

assign p_cast4_cast_fu_677_p1 = grp_fu_536_p4;

assign p_cast5_cast_fu_910_p1 = $signed(reg_590);

assign p_cast6_cast_fu_932_p1 = grp_fu_536_p4;

assign p_cast7_cast_fu_947_p1 = grp_fu_545_p4;

assign p_cast8_cast_fu_921_p1 = $signed(reg_596);

assign p_cast9_cast_fu_816_p1 = $signed(p_cast9_reg_1169);

assign p_cast_cast_fu_655_p1 = grp_fu_518_p4;

assign sext_ln191_fu_734_p0 = current_iteration_fu_202;

assign sext_ln191_fu_734_p1 = sext_ln191_fu_734_p0;

assign shl_ln_fu_758_p3 = {{trunc_ln194_1_fu_754_p1}, {1'd0}};

assign tmp_1_fu_790_p3 = {{mul_ln194_reg_1146}, {6'd0}};

assign tmp_2_fu_830_p3 = {{mul_ln194_reg_1146}, {6'd0}};

assign tmp_3_fu_782_p3 = control_assign_fu_166[32'd2];

assign trunc_ln131_fu_620_p1 = control[2:0];

assign trunc_ln194_1_fu_754_p1 = k_assign_fu_162[27:0];

assign trunc_ln194_fu_747_p1 = n_assign_fu_158[28:0];

assign trunc_ln199_fu_826_p1 = control_assign_fu_166[0:0];

assign trunc_ln204_fu_891_p1 = sub_iterations_assign_fu_174[31:0];

assign trunc_ln215_fu_943_p1 = control_assign_fu_166[0:0];

endmodule //kmeans_top


// Content from kmeans_top_kmeans.v
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2022.2 (64-bit)
// Version: 2022.2
// Copyright (C) Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module kmeans_top_kmeans (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        node_x_coords_address0,
        node_x_coords_ce0,
        node_x_coords_q0,
        node_x_coords_address1,
        node_x_coords_ce1,
        node_x_coords_q1,
        node_y_coords_address0,
        node_y_coords_ce0,
        node_y_coords_q0,
        node_y_coords_address1,
        node_y_coords_ce1,
        node_y_coords_q1,
        node_cluster_assignments_address1,
        node_cluster_assignments_ce1,
        node_cluster_assignments_we1,
        node_cluster_assignments_d1,
        centroid_x_coords_address0,
        centroid_x_coords_ce0,
        centroid_x_coords_we0,
        centroid_x_coords_d0,
        centroid_x_coords_q0,
        centroid_x_coords_address1,
        centroid_x_coords_ce1,
        centroid_x_coords_q1,
        centroid_y_coords_address0,
        centroid_y_coords_ce0,
        centroid_y_coords_we0,
        centroid_y_coords_d0,
        centroid_y_coords_q0,
        centroid_y_coords_address1,
        centroid_y_coords_ce1,
        centroid_y_coords_q1,
        max_iterations,
        n,
        k,
        ap_return
);

parameter    ap_ST_fsm_state1 = 150'd1;
parameter    ap_ST_fsm_state2 = 150'd2;
parameter    ap_ST_fsm_state3 = 150'd4;
parameter    ap_ST_fsm_state4 = 150'd8;
parameter    ap_ST_fsm_state5 = 150'd16;
parameter    ap_ST_fsm_state6 = 150'd32;
parameter    ap_ST_fsm_state7 = 150'd64;
parameter    ap_ST_fsm_state8 = 150'd128;
parameter    ap_ST_fsm_state9 = 150'd256;
parameter    ap_ST_fsm_state10 = 150'd512;
parameter    ap_ST_fsm_state11 = 150'd1024;
parameter    ap_ST_fsm_state12 = 150'd2048;
parameter    ap_ST_fsm_state13 = 150'd4096;
parameter    ap_ST_fsm_state14 = 150'd8192;
parameter    ap_ST_fsm_state15 = 150'd16384;
parameter    ap_ST_fsm_state16 = 150'd32768;
parameter    ap_ST_fsm_state17 = 150'd65536;
parameter    ap_ST_fsm_state18 = 150'd131072;
parameter    ap_ST_fsm_state19 = 150'd262144;
parameter    ap_ST_fsm_state20 = 150'd524288;
parameter    ap_ST_fsm_state21 = 150'd1048576;
parameter    ap_ST_fsm_state22 = 150'd2097152;
parameter    ap_ST_fsm_state23 = 150'd4194304;
parameter    ap_ST_fsm_state24 = 150'd8388608;
parameter    ap_ST_fsm_state25 = 150'd16777216;
parameter    ap_ST_fsm_state26 = 150'd33554432;
parameter    ap_ST_fsm_state27 = 150'd67108864;
parameter    ap_ST_fsm_state28 = 150'd134217728;
parameter    ap_ST_fsm_state29 = 150'd268435456;
parameter    ap_ST_fsm_state30 = 150'd536870912;
parameter    ap_ST_fsm_state31 = 150'd1073741824;
parameter    ap_ST_fsm_state32 = 150'd2147483648;
parameter    ap_ST_fsm_state33 = 150'd4294967296;
parameter    ap_ST_fsm_state34 = 150'd8589934592;
parameter    ap_ST_fsm_state35 = 150'd17179869184;
parameter    ap_ST_fsm_state36 = 150'd34359738368;
parameter    ap_ST_fsm_state37 = 150'd68719476736;
parameter    ap_ST_fsm_state38 = 150'd137438953472;
parameter    ap_ST_fsm_state39 = 150'd274877906944;
parameter    ap_ST_fsm_state40 = 150'd549755813888;
parameter    ap_ST_fsm_state41 = 150'd1099511627776;
parameter    ap_ST_fsm_state42 = 150'd2199023255552;
parameter    ap_ST_fsm_state43 = 150'd4398046511104;
parameter    ap_ST_fsm_state44 = 150'd8796093022208;
parameter    ap_ST_fsm_state45 = 150'd17592186044416;
parameter    ap_ST_fsm_state46 = 150'd35184372088832;
parameter    ap_ST_fsm_state47 = 150'd70368744177664;
parameter    ap_ST_fsm_state48 = 150'd140737488355328;
parameter    ap_ST_fsm_state49 = 150'd281474976710656;
parameter    ap_ST_fsm_state50 = 150'd562949953421312;
parameter    ap_ST_fsm_state51 = 150'd1125899906842624;
parameter    ap_ST_fsm_state52 = 150'd2251799813685248;
parameter    ap_ST_fsm_state53 = 150'd4503599627370496;
parameter    ap_ST_fsm_state54 = 150'd9007199254740992;
parameter    ap_ST_fsm_state55 = 150'd18014398509481984;
parameter    ap_ST_fsm_state56 = 150'd36028797018963968;
parameter    ap_ST_fsm_state57 = 150'd72057594037927936;
parameter    ap_ST_fsm_state58 = 150'd144115188075855872;
parameter    ap_ST_fsm_state59 = 150'd288230376151711744;
parameter    ap_ST_fsm_state60 = 150'd576460752303423488;
parameter    ap_ST_fsm_state61 = 150'd1152921504606846976;
parameter    ap_ST_fsm_state62 = 150'd2305843009213693952;
parameter    ap_ST_fsm_state63 = 150'd4611686018427387904;
parameter    ap_ST_fsm_state64 = 150'd9223372036854775808;
parameter    ap_ST_fsm_state65 = 150'd18446744073709551616;
parameter    ap_ST_fsm_state66 = 150'd36893488147419103232;
parameter    ap_ST_fsm_state67 = 150'd73786976294838206464;
parameter    ap_ST_fsm_state68 = 150'd147573952589676412928;
parameter    ap_ST_fsm_state69 = 150'd295147905179352825856;
parameter    ap_ST_fsm_state70 = 150'd590295810358705651712;
parameter    ap_ST_fsm_state71 = 150'd1180591620717411303424;
parameter    ap_ST_fsm_state72 = 150'd2361183241434822606848;
parameter    ap_ST_fsm_state73 = 150'd4722366482869645213696;
parameter    ap_ST_fsm_state74 = 150'd9444732965739290427392;
parameter    ap_ST_fsm_state75 = 150'd18889465931478580854784;
parameter    ap_ST_fsm_state76 = 150'd37778931862957161709568;
parameter    ap_ST_fsm_state77 = 150'd75557863725914323419136;
parameter    ap_ST_fsm_state78 = 150'd151115727451828646838272;
parameter    ap_ST_fsm_state79 = 150'd302231454903657293676544;
parameter    ap_ST_fsm_state80 = 150'd604462909807314587353088;
parameter    ap_ST_fsm_state81 = 150'd1208925819614629174706176;
parameter    ap_ST_fsm_state82 = 150'd2417851639229258349412352;
parameter    ap_ST_fsm_state83 = 150'd4835703278458516698824704;
parameter    ap_ST_fsm_state84 = 150'd9671406556917033397649408;
parameter    ap_ST_fsm_state85 = 150'd19342813113834066795298816;
parameter    ap_ST_fsm_state86 = 150'd38685626227668133590597632;
parameter    ap_ST_fsm_state87 = 150'd77371252455336267181195264;
parameter    ap_ST_fsm_state88 = 150'd154742504910672534362390528;
parameter    ap_ST_fsm_state89 = 150'd309485009821345068724781056;
parameter    ap_ST_fsm_state90 = 150'd618970019642690137449562112;
parameter    ap_ST_fsm_state91 = 150'd1237940039285380274899124224;
parameter    ap_ST_fsm_state92 = 150'd2475880078570760549798248448;
parameter    ap_ST_fsm_state93 = 150'd4951760157141521099596496896;
parameter    ap_ST_fsm_state94 = 150'd9903520314283042199192993792;
parameter    ap_ST_fsm_state95 = 150'd19807040628566084398385987584;
parameter    ap_ST_fsm_state96 = 150'd39614081257132168796771975168;
parameter    ap_ST_fsm_state97 = 150'd79228162514264337593543950336;
parameter    ap_ST_fsm_state98 = 150'd158456325028528675187087900672;
parameter    ap_ST_fsm_state99 = 150'd316912650057057350374175801344;
parameter    ap_ST_fsm_state100 = 150'd633825300114114700748351602688;
parameter    ap_ST_fsm_state101 = 150'd1267650600228229401496703205376;
parameter    ap_ST_fsm_state102 = 150'd2535301200456458802993406410752;
parameter    ap_ST_fsm_state103 = 150'd5070602400912917605986812821504;
parameter    ap_ST_fsm_state104 = 150'd10141204801825835211973625643008;
parameter    ap_ST_fsm_state105 = 150'd20282409603651670423947251286016;
parameter    ap_ST_fsm_state106 = 150'd40564819207303340847894502572032;
parameter    ap_ST_fsm_state107 = 150'd81129638414606681695789005144064;
parameter    ap_ST_fsm_state108 = 150'd162259276829213363391578010288128;
parameter    ap_ST_fsm_state109 = 150'd324518553658426726783156020576256;
parameter    ap_ST_fsm_state110 = 150'd649037107316853453566312041152512;
parameter    ap_ST_fsm_state111 = 150'd1298074214633706907132624082305024;
parameter    ap_ST_fsm_state112 = 150'd2596148429267413814265248164610048;
parameter    ap_ST_fsm_state113 = 150'd5192296858534827628530496329220096;
parameter    ap_ST_fsm_state114 = 150'd10384593717069655257060992658440192;
parameter    ap_ST_fsm_state115 = 150'd20769187434139310514121985316880384;
parameter    ap_ST_fsm_state116 = 150'd41538374868278621028243970633760768;
parameter    ap_ST_fsm_state117 = 150'd83076749736557242056487941267521536;
parameter    ap_ST_fsm_state118 = 150'd166153499473114484112975882535043072;
parameter    ap_ST_fsm_state119 = 150'd332306998946228968225951765070086144;
parameter    ap_ST_fsm_state120 = 150'd664613997892457936451903530140172288;
parameter    ap_ST_fsm_state121 = 150'd1329227995784915872903807060280344576;
parameter    ap_ST_fsm_state122 = 150'd2658455991569831745807614120560689152;
parameter    ap_ST_fsm_state123 = 150'd5316911983139663491615228241121378304;
parameter    ap_ST_fsm_state124 = 150'd10633823966279326983230456482242756608;
parameter    ap_ST_fsm_state125 = 150'd21267647932558653966460912964485513216;
parameter    ap_ST_fsm_state126 = 150'd42535295865117307932921825928971026432;
parameter    ap_ST_fsm_state127 = 150'd85070591730234615865843651857942052864;
parameter    ap_ST_fsm_state128 = 150'd170141183460469231731687303715884105728;
parameter    ap_ST_fsm_state129 = 150'd340282366920938463463374607431768211456;
parameter    ap_ST_fsm_state130 = 150'd680564733841876926926749214863536422912;
parameter    ap_ST_fsm_state131 = 150'd1361129467683753853853498429727072845824;
parameter    ap_ST_fsm_state132 = 150'd2722258935367507707706996859454145691648;
parameter    ap_ST_fsm_state133 = 150'd5444517870735015415413993718908291383296;
parameter    ap_ST_fsm_state134 = 150'd10889035741470030830827987437816582766592;
parameter    ap_ST_fsm_state135 = 150'd21778071482940061661655974875633165533184;
parameter    ap_ST_fsm_state136 = 150'd43556142965880123323311949751266331066368;
parameter    ap_ST_fsm_state137 = 150'd87112285931760246646623899502532662132736;
parameter    ap_ST_fsm_state138 = 150'd174224571863520493293247799005065324265472;
parameter    ap_ST_fsm_state139 = 150'd348449143727040986586495598010130648530944;
parameter    ap_ST_fsm_state140 = 150'd696898287454081973172991196020261297061888;
parameter    ap_ST_fsm_state141 = 150'd1393796574908163946345982392040522594123776;
parameter    ap_ST_fsm_state142 = 150'd2787593149816327892691964784081045188247552;
parameter    ap_ST_fsm_state143 = 150'd5575186299632655785383929568162090376495104;
parameter    ap_ST_fsm_state144 = 150'd11150372599265311570767859136324180752990208;
parameter    ap_ST_fsm_state145 = 150'd22300745198530623141535718272648361505980416;
parameter    ap_ST_fsm_state146 = 150'd44601490397061246283071436545296723011960832;
parameter    ap_ST_fsm_state147 = 150'd89202980794122492566142873090593446023921664;
parameter    ap_ST_fsm_state148 = 150'd178405961588244985132285746181186892047843328;
parameter    ap_ST_fsm_state149 = 150'd356811923176489970264571492362373784095686656;
parameter    ap_ST_fsm_state150 = 150'd713623846352979940529142984724747568191373312;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
output  [12:0] node_x_coords_address0;
output   node_x_coords_ce0;
input  [63:0] node_x_coords_q0;
output  [12:0] node_x_coords_address1;
output   node_x_coords_ce1;
input  [63:0] node_x_coords_q1;
output  [12:0] node_y_coords_address0;
output   node_y_coords_ce0;
input  [63:0] node_y_coords_q0;
output  [12:0] node_y_coords_address1;
output   node_y_coords_ce1;
input  [63:0] node_y_coords_q1;
output  [12:0] node_cluster_assignments_address1;
output   node_cluster_assignments_ce1;
output   node_cluster_assignments_we1;
output  [63:0] node_cluster_assignments_d1;
output  [7:0] centroid_x_coords_address0;
output   centroid_x_coords_ce0;
output   centroid_x_coords_we0;
output  [63:0] centroid_x_coords_d0;
input  [63:0] centroid_x_coords_q0;
output  [7:0] centroid_x_coords_address1;
output   centroid_x_coords_ce1;
input  [63:0] centroid_x_coords_q1;
output  [7:0] centroid_y_coords_address0;
output   centroid_y_coords_ce0;
output   centroid_y_coords_we0;
output  [63:0] centroid_y_coords_d0;
input  [63:0] centroid_y_coords_q0;
output  [7:0] centroid_y_coords_address1;
output   centroid_y_coords_ce1;
input  [63:0] centroid_y_coords_q1;
input  [63:0] max_iterations;
input  [31:0] n;
input  [31:0] k;
output  [0:0] ap_return;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg[12:0] node_x_coords_address0;
reg node_x_coords_ce0;
reg node_x_coords_ce1;
reg[12:0] node_y_coords_address0;
reg node_y_coords_ce0;
reg node_y_coords_ce1;
reg node_cluster_assignments_ce1;
reg node_cluster_assignments_we1;
reg[7:0] centroid_x_coords_address0;
reg centroid_x_coords_ce0;
reg centroid_x_coords_we0;
reg centroid_x_coords_ce1;
reg[7:0] centroid_y_coords_address0;
reg centroid_y_coords_ce0;
reg centroid_y_coords_we0;
reg centroid_y_coords_ce1;
reg[0:0] ap_return;

(* fsm_encoding = "none" *) reg   [149:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
wire   [15:0] cluster_cardinality_next_q0;
reg   [15:0] reg_389;
wire    ap_CS_fsm_state9;
wire    ap_CS_fsm_state79;
wire   [30:0] empty_fu_393_p1;
reg   [30:0] empty_reg_602;
wire   [0:0] empty_76_fu_402_p2;
reg   [0:0] empty_76_reg_619;
wire   [33:0] tmp_fu_408_p3;
reg   [33:0] tmp_reg_623;
wire   [0:0] cmp165_fu_416_p2;
reg   [0:0] cmp165_reg_628;
wire   [31:0] current_iteration_3_fu_430_p2;
reg   [31:0] current_iteration_3_reg_632;
wire    ap_CS_fsm_state2;
wire   [13:0] add_ln69_fu_449_p2;
reg   [13:0] add_ln69_reg_640;
wire    ap_CS_fsm_state4;
wire   [12:0] trunc_ln37_fu_464_p1;
reg   [12:0] trunc_ln37_reg_648;
wire   [0:0] icmp_ln69_fu_459_p2;
wire    ap_CS_fsm_state6;
reg   [7:0] centroid_x_coords_next_addr_reg_663;
reg   [7:0] centroid_y_coords_next_addr_reg_668;
reg   [7:0] cluster_cardinality_next_addr_reg_673;
wire   [30:0] add_ln101_fu_508_p2;
reg   [30:0] add_ln101_reg_678;
wire    ap_CS_fsm_state8;
wire   [63:0] zext_ln101_fu_514_p1;
reg   [63:0] zext_ln101_reg_683;
wire   [0:0] icmp_ln101_fu_523_p2;
wire   [0:0] grp_fu_383_p2;
reg   [0:0] icmp_ln103_reg_697;
wire   [63:0] centroid_x_coords_next_q0;
wire    ap_CS_fsm_state10;
wire   [30:0] add_ln107_fu_539_p2;
reg   [30:0] add_ln107_reg_716;
wire    ap_CS_fsm_state78;
wire   [63:0] zext_ln107_fu_545_p1;
reg   [63:0] zext_ln107_reg_721;
wire   [0:0] icmp_ln107_fu_554_p2;
reg   [0:0] icmp_ln109_reg_735;
wire   [63:0] centroid_y_coords_next_q0;
wire    ap_CS_fsm_state80;
reg   [7:0] centroid_x_coords_next_address0;
reg    centroid_x_coords_next_ce0;
reg    centroid_x_coords_next_we0;
reg   [63:0] centroid_x_coords_next_d0;
reg   [7:0] centroid_y_coords_next_address0;
reg    centroid_y_coords_next_ce0;
reg    centroid_y_coords_next_we0;
reg   [63:0] centroid_y_coords_next_d0;
reg   [7:0] cluster_cardinality_next_address0;
reg    cluster_cardinality_next_ce0;
reg    cluster_cardinality_next_we0;
reg   [15:0] cluster_cardinality_next_d0;
reg   [7:0] centroid_x_coords_prev_address0;
reg    centroid_x_coords_prev_ce0;
reg    centroid_x_coords_prev_we0;
wire   [63:0] centroid_x_coords_prev_q0;
wire    grp_kmeans_Pipeline_1_fu_332_ap_start;
wire    grp_kmeans_Pipeline_1_fu_332_ap_done;
wire    grp_kmeans_Pipeline_1_fu_332_ap_idle;
wire    grp_kmeans_Pipeline_1_fu_332_ap_ready;
wire   [7:0] grp_kmeans_Pipeline_1_fu_332_centroid_x_coords_address0;
wire    grp_kmeans_Pipeline_1_fu_332_centroid_x_coords_ce0;
wire   [7:0] grp_kmeans_Pipeline_1_fu_332_centroid_x_coords_prev_address0;
wire    grp_kmeans_Pipeline_1_fu_332_centroid_x_coords_prev_ce0;
wire    grp_kmeans_Pipeline_1_fu_332_centroid_x_coords_prev_we0;
wire   [63:0] grp_kmeans_Pipeline_1_fu_332_centroid_x_coords_prev_d0;
wire    grp_kmeans_Pipeline_2_fu_340_ap_start;
wire    grp_kmeans_Pipeline_2_fu_340_ap_done;
wire    grp_kmeans_Pipeline_2_fu_340_ap_idle;
wire    grp_kmeans_Pipeline_2_fu_340_ap_ready;
wire   [7:0] grp_kmeans_Pipeline_2_fu_340_cluster_cardinality_next_address0;
wire    grp_kmeans_Pipeline_2_fu_340_cluster_cardinality_next_ce0;
wire    grp_kmeans_Pipeline_2_fu_340_cluster_cardinality_next_we0;
wire   [15:0] grp_kmeans_Pipeline_2_fu_340_cluster_cardinality_next_d0;
wire    grp_kmeans_Pipeline_3_fu_346_ap_start;
wire    grp_kmeans_Pipeline_3_fu_346_ap_done;
wire    grp_kmeans_Pipeline_3_fu_346_ap_idle;
wire    grp_kmeans_Pipeline_3_fu_346_ap_ready;
wire   [7:0] grp_kmeans_Pipeline_3_fu_346_centroid_x_coords_next_address0;
wire    grp_kmeans_Pipeline_3_fu_346_centroid_x_coords_next_ce0;
wire    grp_kmeans_Pipeline_3_fu_346_centroid_x_coords_next_we0;
wire   [63:0] grp_kmeans_Pipeline_3_fu_346_centroid_x_coords_next_d0;
wire    grp_kmeans_Pipeline_4_fu_352_ap_start;
wire    grp_kmeans_Pipeline_4_fu_352_ap_done;
wire    grp_kmeans_Pipeline_4_fu_352_ap_idle;
wire    grp_kmeans_Pipeline_4_fu_352_ap_ready;
wire   [7:0] grp_kmeans_Pipeline_4_fu_352_centroid_y_coords_next_address0;
wire    grp_kmeans_Pipeline_4_fu_352_centroid_y_coords_next_ce0;
wire    grp_kmeans_Pipeline_4_fu_352_centroid_y_coords_next_we0;
wire   [63:0] grp_kmeans_Pipeline_4_fu_352_centroid_y_coords_next_d0;
wire    grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_ap_start;
wire    grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_ap_done;
wire    grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_ap_idle;
wire    grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_ap_ready;
wire   [12:0] grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_node_x_coords_address0;
wire    grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_node_x_coords_ce0;
wire   [12:0] grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_node_x_coords_address1;
wire    grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_node_x_coords_ce1;
wire   [12:0] grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_node_y_coords_address0;
wire    grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_node_y_coords_ce0;
wire   [12:0] grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_node_y_coords_address1;
wire    grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_node_y_coords_ce1;
wire   [7:0] grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_centroid_y_coords_address0;
wire    grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_centroid_y_coords_ce0;
wire   [7:0] grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_centroid_y_coords_address1;
wire    grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_centroid_y_coords_ce1;
wire   [7:0] grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_centroid_x_coords_address0;
wire    grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_centroid_x_coords_ce0;
wire   [7:0] grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_centroid_x_coords_address1;
wire    grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_centroid_x_coords_ce1;
wire   [31:0] grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_min_dist_index_out;
wire    grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_min_dist_index_out_ap_vld;
wire    grp_kmeans_Pipeline_VITIS_LOOP_116_6_fu_373_ap_start;
wire    grp_kmeans_Pipeline_VITIS_LOOP_116_6_fu_373_ap_done;
wire    grp_kmeans_Pipeline_VITIS_LOOP_116_6_fu_373_ap_idle;
wire    grp_kmeans_Pipeline_VITIS_LOOP_116_6_fu_373_ap_ready;
wire   [7:0] grp_kmeans_Pipeline_VITIS_LOOP_116_6_fu_373_centroid_y_coords_address0;
wire    grp_kmeans_Pipeline_VITIS_LOOP_116_6_fu_373_centroid_y_coords_ce0;
wire   [7:0] grp_kmeans_Pipeline_VITIS_LOOP_116_6_fu_373_centroid_x_coords_prev_address0;
wire    grp_kmeans_Pipeline_VITIS_LOOP_116_6_fu_373_centroid_x_coords_prev_ce0;
wire   [7:0] grp_kmeans_Pipeline_VITIS_LOOP_116_6_fu_373_centroid_x_coords_address0;
wire    grp_kmeans_Pipeline_VITIS_LOOP_116_6_fu_373_centroid_x_coords_ce0;
wire   [1:0] grp_kmeans_Pipeline_VITIS_LOOP_116_6_fu_373_ap_return;
wire   [0:0] ap_phi_mux_converged_phi_fu_263_p4;
reg   [0:0] converged_reg_259;
wire    ap_CS_fsm_state149;
reg   [13:0] i_reg_270;
wire    ap_CS_fsm_state7;
wire    ap_CS_fsm_state3;
reg    ap_block_state3_on_subcall_done;
reg   [30:0] i_1_reg_282;
wire    ap_CS_fsm_state77;
reg   [30:0] i_2_reg_293;
wire    ap_CS_fsm_state147;
reg   [0:0] converged_1_reg_304;
wire    ap_CS_fsm_state148;
reg    ap_block_state148_on_subcall_done;
wire   [0:0] cond_fu_570_p2;
reg   [0:0] converged_0_lcssa_reg_319;
wire   [0:0] icmp_ln53_fu_443_p2;
reg    grp_kmeans_Pipeline_1_fu_332_ap_start_reg;
reg    grp_kmeans_Pipeline_2_fu_340_ap_start_reg;
reg    grp_kmeans_Pipeline_3_fu_346_ap_start_reg;
reg    grp_kmeans_Pipeline_4_fu_352_ap_start_reg;
reg    grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_ap_start_reg;
wire    ap_CS_fsm_state5;
reg    grp_kmeans_Pipeline_VITIS_LOOP_116_6_fu_373_ap_start_reg;
wire   [63:0] zext_ln69_fu_469_p1;
wire  signed [63:0] sext_ln94_fu_479_p1;
reg   [31:0] current_iteration_fu_80;
reg   [63:0] max_iterations_assign_fu_88;
wire   [63:0] add_ln95_fu_487_p2;
wire   [63:0] add_ln96_fu_494_p2;
wire   [15:0] add_ln97_fu_501_p2;
wire   [63:0] grp_fu_532_p2;
wire   [63:0] grp_fu_563_p2;
wire   [63:0] zext_ln53_fu_436_p1;
wire   [31:0] zext_ln69_1_fu_455_p1;
wire   [31:0] zext_ln101_1_fu_519_p1;
wire   [15:0] grp_fu_532_p1;
wire   [31:0] zext_ln107_1_fu_550_p1;
wire   [15:0] grp_fu_563_p1;
reg    grp_fu_532_ap_start;
wire    grp_fu_532_ap_done;
reg    grp_fu_563_ap_start;
wire    grp_fu_563_ap_done;
reg   [0:0] ap_return_preg;
wire    ap_CS_fsm_state150;
reg   [149:0] ap_NS_fsm;
reg    ap_ST_fsm_state1_blk;
wire    ap_ST_fsm_state2_blk;
reg    ap_ST_fsm_state3_blk;
wire    ap_ST_fsm_state4_blk;
reg    ap_ST_fsm_state5_blk;
wire    ap_ST_fsm_state6_blk;
wire    ap_ST_fsm_state7_blk;
wire    ap_ST_fsm_state8_blk;
wire    ap_ST_fsm_state9_blk;
wire    ap_ST_fsm_state10_blk;
wire    ap_ST_fsm_state11_blk;
wire    ap_ST_fsm_state12_blk;
wire    ap_ST_fsm_state13_blk;
wire    ap_ST_fsm_state14_blk;
wire    ap_ST_fsm_state15_blk;
wire    ap_ST_fsm_state16_blk;
wire    ap_ST_fsm_state17_blk;
wire    ap_ST_fsm_state18_blk;
wire    ap_ST_fsm_state19_blk;
wire    ap_ST_fsm_state20_blk;
wire    ap_ST_fsm_state21_blk;
wire    ap_ST_fsm_state22_blk;
wire    ap_ST_fsm_state23_blk;
wire    ap_ST_fsm_state24_blk;
wire    ap_ST_fsm_state25_blk;
wire    ap_ST_fsm_state26_blk;
wire    ap_ST_fsm_state27_blk;
wire    ap_ST_fsm_state28_blk;
wire    ap_ST_fsm_state29_blk;
wire    ap_ST_fsm_state30_blk;
wire    ap_ST_fsm_state31_blk;
wire    ap_ST_fsm_state32_blk;
wire    ap_ST_fsm_state33_blk;
wire    ap_ST_fsm_state34_blk;
wire    ap_ST_fsm_state35_blk;
wire    ap_ST_fsm_state36_blk;
wire    ap_ST_fsm_state37_blk;
wire    ap_ST_fsm_state38_blk;
wire    ap_ST_fsm_state39_blk;
wire    ap_ST_fsm_state40_blk;
wire    ap_ST_fsm_state41_blk;
wire    ap_ST_fsm_state42_blk;
wire    ap_ST_fsm_state43_blk;
wire    ap_ST_fsm_state44_blk;
wire    ap_ST_fsm_state45_blk;
wire    ap_ST_fsm_state46_blk;
wire    ap_ST_fsm_state47_blk;
wire    ap_ST_fsm_state48_blk;
wire    ap_ST_fsm_state49_blk;
wire    ap_ST_fsm_state50_blk;
wire    ap_ST_fsm_state51_blk;
wire    ap_ST_fsm_state52_blk;
wire    ap_ST_fsm_state53_blk;
wire    ap_ST_fsm_state54_blk;
wire    ap_ST_fsm_state55_blk;
wire    ap_ST_fsm_state56_blk;
wire    ap_ST_fsm_state57_blk;
wire    ap_ST_fsm_state58_blk;
wire    ap_ST_fsm_state59_blk;
wire    ap_ST_fsm_state60_blk;
wire    ap_ST_fsm_state61_blk;
wire    ap_ST_fsm_state62_blk;
wire    ap_ST_fsm_state63_blk;
wire    ap_ST_fsm_state64_blk;
wire    ap_ST_fsm_state65_blk;
wire    ap_ST_fsm_state66_blk;
wire    ap_ST_fsm_state67_blk;
wire    ap_ST_fsm_state68_blk;
wire    ap_ST_fsm_state69_blk;
wire    ap_ST_fsm_state70_blk;
wire    ap_ST_fsm_state71_blk;
wire    ap_ST_fsm_state72_blk;
wire    ap_ST_fsm_state73_blk;
wire    ap_ST_fsm_state74_blk;
wire    ap_ST_fsm_state75_blk;
wire    ap_ST_fsm_state76_blk;
wire    ap_ST_fsm_state77_blk;
wire    ap_ST_fsm_state78_blk;
wire    ap_ST_fsm_state79_blk;
wire    ap_ST_fsm_state80_blk;
wire    ap_ST_fsm_state81_blk;
wire    ap_ST_fsm_state82_blk;
wire    ap_ST_fsm_state83_blk;
wire    ap_ST_fsm_state84_blk;
wire    ap_ST_fsm_state85_blk;
wire    ap_ST_fsm_state86_blk;
wire    ap_ST_fsm_state87_blk;
wire    ap_ST_fsm_state88_blk;
wire    ap_ST_fsm_state89_blk;
wire    ap_ST_fsm_state90_blk;
wire    ap_ST_fsm_state91_blk;
wire    ap_ST_fsm_state92_blk;
wire    ap_ST_fsm_state93_blk;
wire    ap_ST_fsm_state94_blk;
wire    ap_ST_fsm_state95_blk;
wire    ap_ST_fsm_state96_blk;
wire    ap_ST_fsm_state97_blk;
wire    ap_ST_fsm_state98_blk;
wire    ap_ST_fsm_state99_blk;
wire    ap_ST_fsm_state100_blk;
wire    ap_ST_fsm_state101_blk;
wire    ap_ST_fsm_state102_blk;
wire    ap_ST_fsm_state103_blk;
wire    ap_ST_fsm_state104_blk;
wire    ap_ST_fsm_state105_blk;
wire    ap_ST_fsm_state106_blk;
wire    ap_ST_fsm_state107_blk;
wire    ap_ST_fsm_state108_blk;
wire    ap_ST_fsm_state109_blk;
wire    ap_ST_fsm_state110_blk;
wire    ap_ST_fsm_state111_blk;
wire    ap_ST_fsm_state112_blk;
wire    ap_ST_fsm_state113_blk;
wire    ap_ST_fsm_state114_blk;
wire    ap_ST_fsm_state115_blk;
wire    ap_ST_fsm_state116_blk;
wire    ap_ST_fsm_state117_blk;
wire    ap_ST_fsm_state118_blk;
wire    ap_ST_fsm_state119_blk;
wire    ap_ST_fsm_state120_blk;
wire    ap_ST_fsm_state121_blk;
wire    ap_ST_fsm_state122_blk;
wire    ap_ST_fsm_state123_blk;
wire    ap_ST_fsm_state124_blk;
wire    ap_ST_fsm_state125_blk;
wire    ap_ST_fsm_state126_blk;
wire    ap_ST_fsm_state127_blk;
wire    ap_ST_fsm_state128_blk;
wire    ap_ST_fsm_state129_blk;
wire    ap_ST_fsm_state130_blk;
wire    ap_ST_fsm_state131_blk;
wire    ap_ST_fsm_state132_blk;
wire    ap_ST_fsm_state133_blk;
wire    ap_ST_fsm_state134_blk;
wire    ap_ST_fsm_state135_blk;
wire    ap_ST_fsm_state136_blk;
wire    ap_ST_fsm_state137_blk;
wire    ap_ST_fsm_state138_blk;
wire    ap_ST_fsm_state139_blk;
wire    ap_ST_fsm_state140_blk;
wire    ap_ST_fsm_state141_blk;
wire    ap_ST_fsm_state142_blk;
wire    ap_ST_fsm_state143_blk;
wire    ap_ST_fsm_state144_blk;
wire    ap_ST_fsm_state145_blk;
wire    ap_ST_fsm_state146_blk;
wire    ap_ST_fsm_state147_blk;
reg    ap_ST_fsm_state148_blk;
wire    ap_ST_fsm_state149_blk;
wire    ap_ST_fsm_state150_blk;
wire   [63:0] grp_fu_532_p10;
wire   [63:0] grp_fu_563_p10;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_CS_fsm = 150'd1;
#0 grp_kmeans_Pipeline_1_fu_332_ap_start_reg = 1'b0;
#0 grp_kmeans_Pipeline_2_fu_340_ap_start_reg = 1'b0;
#0 grp_kmeans_Pipeline_3_fu_346_ap_start_reg = 1'b0;
#0 grp_kmeans_Pipeline_4_fu_352_ap_start_reg = 1'b0;
#0 grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_ap_start_reg = 1'b0;
#0 grp_kmeans_Pipeline_VITIS_LOOP_116_6_fu_373_ap_start_reg = 1'b0;
#0 ap_return_preg = 1'd0;
end

kmeans_top_kmeans_centroid_x_coords_next_RAM_AUTO_1R1W #(
    .DataWidth( 64 ),
    .AddressRange( 256 ),
    .AddressWidth( 8 ))
centroid_x_coords_next_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(centroid_x_coords_next_address0),
    .ce0(centroid_x_coords_next_ce0),
    .we0(centroid_x_coords_next_we0),
    .d0(centroid_x_coords_next_d0),
    .q0(centroid_x_coords_next_q0)
);

kmeans_top_kmeans_centroid_x_coords_next_RAM_AUTO_1R1W #(
    .DataWidth( 64 ),
    .AddressRange( 256 ),
    .AddressWidth( 8 ))
centroid_y_coords_next_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(centroid_y_coords_next_address0),
    .ce0(centroid_y_coords_next_ce0),
    .we0(centroid_y_coords_next_we0),
    .d0(centroid_y_coords_next_d0),
    .q0(centroid_y_coords_next_q0)
);

kmeans_top_kmeans_cluster_cardinality_next_RAM_AUTO_1R1W #(
    .DataWidth( 16 ),
    .AddressRange( 256 ),
    .AddressWidth( 8 ))
cluster_cardinality_next_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(cluster_cardinality_next_address0),
    .ce0(cluster_cardinality_next_ce0),
    .we0(cluster_cardinality_next_we0),
    .d0(cluster_cardinality_next_d0),
    .q0(cluster_cardinality_next_q0)
);

kmeans_top_kmeans_centroid_x_coords_next_RAM_AUTO_1R1W #(
    .DataWidth( 64 ),
    .AddressRange( 256 ),
    .AddressWidth( 8 ))
centroid_x_coords_prev_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(centroid_x_coords_prev_address0),
    .ce0(centroid_x_coords_prev_ce0),
    .we0(centroid_x_coords_prev_we0),
    .d0(grp_kmeans_Pipeline_1_fu_332_centroid_x_coords_prev_d0),
    .q0(centroid_x_coords_prev_q0)
);

kmeans_top_kmeans_Pipeline_1 grp_kmeans_Pipeline_1_fu_332(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(grp_kmeans_Pipeline_1_fu_332_ap_start),
    .ap_done(grp_kmeans_Pipeline_1_fu_332_ap_done),
    .ap_idle(grp_kmeans_Pipeline_1_fu_332_ap_idle),
    .ap_ready(grp_kmeans_Pipeline_1_fu_332_ap_ready),
    .centroid_x_coords_address0(grp_kmeans_Pipeline_1_fu_332_centroid_x_coords_address0),
    .centroid_x_coords_ce0(grp_kmeans_Pipeline_1_fu_332_centroid_x_coords_ce0),
    .centroid_x_coords_q0(centroid_x_coords_q0),
    .centroid_x_coords_prev_address0(grp_kmeans_Pipeline_1_fu_332_centroid_x_coords_prev_address0),
    .centroid_x_coords_prev_ce0(grp_kmeans_Pipeline_1_fu_332_centroid_x_coords_prev_ce0),
    .centroid_x_coords_prev_we0(grp_kmeans_Pipeline_1_fu_332_centroid_x_coords_prev_we0),
    .centroid_x_coords_prev_d0(grp_kmeans_Pipeline_1_fu_332_centroid_x_coords_prev_d0),
    .p_cast12(k)
);

kmeans_top_kmeans_Pipeline_2 grp_kmeans_Pipeline_2_fu_340(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(grp_kmeans_Pipeline_2_fu_340_ap_start),
    .ap_done(grp_kmeans_Pipeline_2_fu_340_ap_done),
    .ap_idle(grp_kmeans_Pipeline_2_fu_340_ap_idle),
    .ap_ready(grp_kmeans_Pipeline_2_fu_340_ap_ready),
    .cluster_cardinality_next_address0(grp_kmeans_Pipeline_2_fu_340_cluster_cardinality_next_address0),
    .cluster_cardinality_next_ce0(grp_kmeans_Pipeline_2_fu_340_cluster_cardinality_next_ce0),
    .cluster_cardinality_next_we0(grp_kmeans_Pipeline_2_fu_340_cluster_cardinality_next_we0),
    .cluster_cardinality_next_d0(grp_kmeans_Pipeline_2_fu_340_cluster_cardinality_next_d0),
    .p_cast3_cast(tmp_reg_623)
);

kmeans_top_kmeans_Pipeline_3 grp_kmeans_Pipeline_3_fu_346(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(grp_kmeans_Pipeline_3_fu_346_ap_start),
    .ap_done(grp_kmeans_Pipeline_3_fu_346_ap_done),
    .ap_idle(grp_kmeans_Pipeline_3_fu_346_ap_idle),
    .ap_ready(grp_kmeans_Pipeline_3_fu_346_ap_ready),
    .centroid_x_coords_next_address0(grp_kmeans_Pipeline_3_fu_346_centroid_x_coords_next_address0),
    .centroid_x_coords_next_ce0(grp_kmeans_Pipeline_3_fu_346_centroid_x_coords_next_ce0),
    .centroid_x_coords_next_we0(grp_kmeans_Pipeline_3_fu_346_centroid_x_coords_next_we0),
    .centroid_x_coords_next_d0(grp_kmeans_Pipeline_3_fu_346_centroid_x_coords_next_d0),
    .k_cast2_cast_cast(k)
);

kmeans_top_kmeans_Pipeline_4 grp_kmeans_Pipeline_4_fu_352(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(grp_kmeans_Pipeline_4_fu_352_ap_start),
    .ap_done(grp_kmeans_Pipeline_4_fu_352_ap_done),
    .ap_idle(grp_kmeans_Pipeline_4_fu_352_ap_idle),
    .ap_ready(grp_kmeans_Pipeline_4_fu_352_ap_ready),
    .centroid_y_coords_next_address0(grp_kmeans_Pipeline_4_fu_352_centroid_y_coords_next_address0),
    .centroid_y_coords_next_ce0(grp_kmeans_Pipeline_4_fu_352_centroid_y_coords_next_ce0),
    .centroid_y_coords_next_we0(grp_kmeans_Pipeline_4_fu_352_centroid_y_coords_next_we0),
    .centroid_y_coords_next_d0(grp_kmeans_Pipeline_4_fu_352_centroid_y_coords_next_d0),
    .k_cast2_cast_cast(k)
);

kmeans_top_kmeans_Pipeline_VITIS_LOOP_73_3 grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_ap_start),
    .ap_done(grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_ap_done),
    .ap_idle(grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_ap_idle),
    .ap_ready(grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_ap_ready),
    .node_x_coords_address0(grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_node_x_coords_address0),
    .node_x_coords_ce0(grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_node_x_coords_ce0),
    .node_x_coords_q0(node_x_coords_q0),
    .node_x_coords_address1(grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_node_x_coords_address1),
    .node_x_coords_ce1(grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_node_x_coords_ce1),
    .node_x_coords_q1(node_x_coords_q1),
    .zext_ln69(trunc_ln37_reg_648),
    .node_y_coords_address0(grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_node_y_coords_address0),
    .node_y_coords_ce0(grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_node_y_coords_ce0),
    .node_y_coords_q0(node_y_coords_q0),
    .node_y_coords_address1(grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_node_y_coords_address1),
    .node_y_coords_ce1(grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_node_y_coords_ce1),
    .node_y_coords_q1(node_y_coords_q1),
    .k(k),
    .centroid_y_coords_address0(grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_centroid_y_coords_address0),
    .centroid_y_coords_ce0(grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_centroid_y_coords_ce0),
    .centroid_y_coords_q0(centroid_y_coords_q0),
    .centroid_y_coords_address1(grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_centroid_y_coords_address1),
    .centroid_y_coords_ce1(grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_centroid_y_coords_ce1),
    .centroid_y_coords_q1(centroid_y_coords_q1),
    .centroid_x_coords_address0(grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_centroid_x_coords_address0),
    .centroid_x_coords_ce0(grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_centroid_x_coords_ce0),
    .centroid_x_coords_q0(centroid_x_coords_q0),
    .centroid_x_coords_address1(grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_centroid_x_coords_address1),
    .centroid_x_coords_ce1(grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_centroid_x_coords_ce1),
    .centroid_x_coords_q1(centroid_x_coords_q1),
    .min_dist_index_out(grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_min_dist_index_out),
    .min_dist_index_out_ap_vld(grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_min_dist_index_out_ap_vld)
);

kmeans_top_kmeans_Pipeline_VITIS_LOOP_116_6 grp_kmeans_Pipeline_VITIS_LOOP_116_6_fu_373(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(grp_kmeans_Pipeline_VITIS_LOOP_116_6_fu_373_ap_start),
    .ap_done(grp_kmeans_Pipeline_VITIS_LOOP_116_6_fu_373_ap_done),
    .ap_idle(grp_kmeans_Pipeline_VITIS_LOOP_116_6_fu_373_ap_idle),
    .ap_ready(grp_kmeans_Pipeline_VITIS_LOOP_116_6_fu_373_ap_ready),
    .k(empty_reg_602),
    .centroid_y_coords_address0(grp_kmeans_Pipeline_VITIS_LOOP_116_6_fu_373_centroid_y_coords_address0),
    .centroid_y_coords_ce0(grp_kmeans_Pipeline_VITIS_LOOP_116_6_fu_373_centroid_y_coords_ce0),
    .centroid_y_coords_q0(centroid_y_coords_q0),
    .centroid_x_coords_prev_address0(grp_kmeans_Pipeline_VITIS_LOOP_116_6_fu_373_centroid_x_coords_prev_address0),
    .centroid_x_coords_prev_ce0(grp_kmeans_Pipeline_VITIS_LOOP_116_6_fu_373_centroid_x_coords_prev_ce0),
    .centroid_x_coords_prev_q0(centroid_x_coords_prev_q0),
    .centroid_x_coords_address0(grp_kmeans_Pipeline_VITIS_LOOP_116_6_fu_373_centroid_x_coords_address0),
    .centroid_x_coords_ce0(grp_kmeans_Pipeline_VITIS_LOOP_116_6_fu_373_centroid_x_coords_ce0),
    .centroid_x_coords_q0(centroid_x_coords_q0),
    .ap_return(grp_kmeans_Pipeline_VITIS_LOOP_116_6_fu_373_ap_return)
);

kmeans_top_udiv_64ns_16ns_64_68_seq_1 #(
    .ID( 1 ),
    .NUM_STAGE( 68 ),
    .din0_WIDTH( 64 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 64 ))
udiv_64ns_16ns_64_68_seq_1_U44(
    .clk(ap_clk),
    .reset(ap_rst),
    .start(grp_fu_532_ap_start),
    .done(grp_fu_532_ap_done),
    .din0(centroid_x_coords_next_q0),
    .din1(grp_fu_532_p1),
    .ce(1'b1),
    .dout(grp_fu_532_p2)
);

kmeans_top_udiv_64ns_16ns_64_68_seq_1 #(
    .ID( 1 ),
    .NUM_STAGE( 68 ),
    .din0_WIDTH( 64 ),
    .din1_WIDTH( 16 ),
    .dout_WIDTH( 64 ))
udiv_64ns_16ns_64_68_seq_1_U45(
    .clk(ap_clk),
    .reset(ap_rst),
    .start(grp_fu_563_ap_start),
    .done(grp_fu_563_ap_done),
    .din0(centroid_y_coords_next_q0),
    .din1(grp_fu_563_p1),
    .ce(1'b1),
    .dout(grp_fu_563_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_return_preg <= 1'd0;
    end else begin
        if ((1'b1 == ap_CS_fsm_state150)) begin
            ap_return_preg <= converged_0_lcssa_reg_319;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        grp_kmeans_Pipeline_1_fu_332_ap_start_reg <= 1'b0;
    end else begin
        if (((icmp_ln53_fu_443_p2 == 1'd1) & (ap_phi_mux_converged_phi_fu_263_p4 == 1'd0) & (empty_76_reg_619 == 1'd0) & (1'b1 == ap_CS_fsm_state2))) begin
            grp_kmeans_Pipeline_1_fu_332_ap_start_reg <= 1'b1;
        end else if ((grp_kmeans_Pipeline_1_fu_332_ap_ready == 1'b1)) begin
            grp_kmeans_Pipeline_1_fu_332_ap_start_reg <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        grp_kmeans_Pipeline_2_fu_340_ap_start_reg <= 1'b0;
    end else begin
        if (((icmp_ln53_fu_443_p2 == 1'd1) & (ap_phi_mux_converged_phi_fu_263_p4 == 1'd0) & (empty_76_reg_619 == 1'd0) & (1'b1 == ap_CS_fsm_state2))) begin
            grp_kmeans_Pipeline_2_fu_340_ap_start_reg <= 1'b1;
        end else if ((grp_kmeans_Pipeline_2_fu_340_ap_ready == 1'b1)) begin
            grp_kmeans_Pipeline_2_fu_340_ap_start_reg <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        grp_kmeans_Pipeline_3_fu_346_ap_start_reg <= 1'b0;
    end else begin
        if (((icmp_ln53_fu_443_p2 == 1'd1) & (ap_phi_mux_converged_phi_fu_263_p4 == 1'd0) & (empty_76_reg_619 == 1'd0) & (1'b1 == ap_CS_fsm_state2))) begin
            grp_kmeans_Pipeline_3_fu_346_ap_start_reg <= 1'b1;
        end else if ((grp_kmeans_Pipeline_3_fu_346_ap_ready == 1'b1)) begin
            grp_kmeans_Pipeline_3_fu_346_ap_start_reg <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        grp_kmeans_Pipeline_4_fu_352_ap_start_reg <= 1'b0;
    end else begin
        if (((icmp_ln53_fu_443_p2 == 1'd1) & (ap_phi_mux_converged_phi_fu_263_p4 == 1'd0) & (empty_76_reg_619 == 1'd0) & (1'b1 == ap_CS_fsm_state2))) begin
            grp_kmeans_Pipeline_4_fu_352_ap_start_reg <= 1'b1;
        end else if ((grp_kmeans_Pipeline_4_fu_352_ap_ready == 1'b1)) begin
            grp_kmeans_Pipeline_4_fu_352_ap_start_reg <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        grp_kmeans_Pipeline_VITIS_LOOP_116_6_fu_373_ap_start_reg <= 1'b0;
    end else begin
        if (((icmp_ln107_fu_554_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state78))) begin
            grp_kmeans_Pipeline_VITIS_LOOP_116_6_fu_373_ap_start_reg <= 1'b1;
        end else if ((grp_kmeans_Pipeline_VITIS_LOOP_116_6_fu_373_ap_ready == 1'b1)) begin
            grp_kmeans_Pipeline_VITIS_LOOP_116_6_fu_373_ap_start_reg <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_ap_start_reg <= 1'b0;
    end else begin
        if (((icmp_ln69_fu_459_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state4))) begin
            grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_ap_start_reg <= 1'b1;
        end else if ((grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_ap_ready == 1'b1)) begin
            grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_ap_start_reg <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        if (((icmp_ln53_fu_443_p2 == 1'd0) & (ap_phi_mux_converged_phi_fu_263_p4 == 1'd0))) begin
            converged_0_lcssa_reg_319 <= 1'd0;
        end else if ((ap_phi_mux_converged_phi_fu_263_p4 == 1'd1)) begin
            converged_0_lcssa_reg_319 <= 1'd1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_state148_on_subcall_done) & (1'b1 == ap_CS_fsm_state148))) begin
        if (((cond_fu_570_p2 == 1'd0) & (cmp165_reg_628 == 1'd1))) begin
            converged_1_reg_304 <= 1'd0;
        end else if (((cond_fu_570_p2 == 1'd1) | (cmp165_reg_628 == 1'd0))) begin
            converged_1_reg_304 <= 1'd1;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state149)) begin
        converged_reg_259 <= converged_1_reg_304;
    end else if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
        converged_reg_259 <= 1'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
        current_iteration_fu_80 <= 32'd0;
    end else if (((1'b0 == ap_block_state148_on_subcall_done) & (1'b1 == ap_CS_fsm_state148))) begin
        current_iteration_fu_80 <= current_iteration_3_reg_632;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln69_fu_459_p2 == 1'd0) & (cmp165_reg_628 == 1'd1) & (1'b1 == ap_CS_fsm_state4))) begin
        i_1_reg_282 <= 31'd0;
    end else if ((1'b1 == ap_CS_fsm_state77)) begin
        i_1_reg_282 <= add_ln101_reg_678;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln101_fu_523_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state8))) begin
        i_2_reg_293 <= 31'd0;
    end else if ((1'b1 == ap_CS_fsm_state147)) begin
        i_2_reg_293 <= add_ln107_reg_716;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_state3_on_subcall_done) & (1'b1 == ap_CS_fsm_state3))) begin
        i_reg_270 <= 14'd0;
    end else if ((1'b1 == ap_CS_fsm_state7)) begin
        i_reg_270 <= add_ln69_reg_640;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state8)) begin
        add_ln101_reg_678 <= add_ln101_fu_508_p2;
        zext_ln101_reg_683[30 : 0] <= zext_ln101_fu_514_p1[30 : 0];
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state78)) begin
        add_ln107_reg_716 <= add_ln107_fu_539_p2;
        zext_ln107_reg_721[30 : 0] <= zext_ln107_fu_545_p1[30 : 0];
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        add_ln69_reg_640 <= add_ln69_fu_449_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state6)) begin
        centroid_x_coords_next_addr_reg_663 <= sext_ln94_fu_479_p1;
        centroid_y_coords_next_addr_reg_668 <= sext_ln94_fu_479_p1;
        cluster_cardinality_next_addr_reg_673 <= sext_ln94_fu_479_p1;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        cmp165_reg_628 <= cmp165_fu_416_p2;
        empty_76_reg_619 <= empty_76_fu_402_p2;
        empty_reg_602 <= empty_fu_393_p1;
        tmp_reg_623[33 : 2] <= tmp_fu_408_p3[33 : 2];
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        current_iteration_3_reg_632 <= current_iteration_3_fu_430_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state9)) begin
        icmp_ln103_reg_697 <= grp_fu_383_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state79)) begin
        icmp_ln109_reg_735 <= grp_fu_383_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
        max_iterations_assign_fu_88 <= max_iterations;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_state79) | (1'b1 == ap_CS_fsm_state9))) begin
        reg_389 <= cluster_cardinality_next_q0;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln69_fu_459_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state4))) begin
        trunc_ln37_reg_648 <= trunc_ln37_fu_464_p1;
    end
end

assign ap_ST_fsm_state100_blk = 1'b0;

assign ap_ST_fsm_state101_blk = 1'b0;

assign ap_ST_fsm_state102_blk = 1'b0;

assign ap_ST_fsm_state103_blk = 1'b0;

assign ap_ST_fsm_state104_blk = 1'b0;

assign ap_ST_fsm_state105_blk = 1'b0;

assign ap_ST_fsm_state106_blk = 1'b0;

assign ap_ST_fsm_state107_blk = 1'b0;

assign ap_ST_fsm_state108_blk = 1'b0;

assign ap_ST_fsm_state109_blk = 1'b0;

assign ap_ST_fsm_state10_blk = 1'b0;

assign ap_ST_fsm_state110_blk = 1'b0;

assign ap_ST_fsm_state111_blk = 1'b0;

assign ap_ST_fsm_state112_blk = 1'b0;

assign ap_ST_fsm_state113_blk = 1'b0;

assign ap_ST_fsm_state114_blk = 1'b0;

assign ap_ST_fsm_state115_blk = 1'b0;

assign ap_ST_fsm_state116_blk = 1'b0;

assign ap_ST_fsm_state117_blk = 1'b0;

assign ap_ST_fsm_state118_blk = 1'b0;

assign ap_ST_fsm_state119_blk = 1'b0;

assign ap_ST_fsm_state11_blk = 1'b0;

assign ap_ST_fsm_state120_blk = 1'b0;

assign ap_ST_fsm_state121_blk = 1'b0;

assign ap_ST_fsm_state122_blk = 1'b0;

assign ap_ST_fsm_state123_blk = 1'b0;

assign ap_ST_fsm_state124_blk = 1'b0;

assign ap_ST_fsm_state125_blk = 1'b0;

assign ap_ST_fsm_state126_blk = 1'b0;

assign ap_ST_fsm_state127_blk = 1'b0;

assign ap_ST_fsm_state128_blk = 1'b0;

assign ap_ST_fsm_state129_blk = 1'b0;

assign ap_ST_fsm_state12_blk = 1'b0;

assign ap_ST_fsm_state130_blk = 1'b0;

assign ap_ST_fsm_state131_blk = 1'b0;

assign ap_ST_fsm_state132_blk = 1'b0;

assign ap_ST_fsm_state133_blk = 1'b0;

assign ap_ST_fsm_state134_blk = 1'b0;

assign ap_ST_fsm_state135_blk = 1'b0;

assign ap_ST_fsm_state136_blk = 1'b0;

assign ap_ST_fsm_state137_blk = 1'b0;

assign ap_ST_fsm_state138_blk = 1'b0;

assign ap_ST_fsm_state139_blk = 1'b0;

assign ap_ST_fsm_state13_blk = 1'b0;

assign ap_ST_fsm_state140_blk = 1'b0;

assign ap_ST_fsm_state141_blk = 1'b0;

assign ap_ST_fsm_state142_blk = 1'b0;

assign ap_ST_fsm_state143_blk = 1'b0;

assign ap_ST_fsm_state144_blk = 1'b0;

assign ap_ST_fsm_state145_blk = 1'b0;

assign ap_ST_fsm_state146_blk = 1'b0;

assign ap_ST_fsm_state147_blk = 1'b0;

always @ (*) begin
    if ((1'b1 == ap_block_state148_on_subcall_done)) begin
        ap_ST_fsm_state148_blk = 1'b1;
    end else begin
        ap_ST_fsm_state148_blk = 1'b0;
    end
end

assign ap_ST_fsm_state149_blk = 1'b0;

assign ap_ST_fsm_state14_blk = 1'b0;

assign ap_ST_fsm_state150_blk = 1'b0;

assign ap_ST_fsm_state15_blk = 1'b0;

assign ap_ST_fsm_state16_blk = 1'b0;

assign ap_ST_fsm_state17_blk = 1'b0;

assign ap_ST_fsm_state18_blk = 1'b0;

assign ap_ST_fsm_state19_blk = 1'b0;

always @ (*) begin
    if ((ap_start == 1'b0)) begin
        ap_ST_fsm_state1_blk = 1'b1;
    end else begin
        ap_ST_fsm_state1_blk = 1'b0;
    end
end

assign ap_ST_fsm_state20_blk = 1'b0;

assign ap_ST_fsm_state21_blk = 1'b0;

assign ap_ST_fsm_state22_blk = 1'b0;

assign ap_ST_fsm_state23_blk = 1'b0;

assign ap_ST_fsm_state24_blk = 1'b0;

assign ap_ST_fsm_state25_blk = 1'b0;

assign ap_ST_fsm_state26_blk = 1'b0;

assign ap_ST_fsm_state27_blk = 1'b0;

assign ap_ST_fsm_state28_blk = 1'b0;

assign ap_ST_fsm_state29_blk = 1'b0;

assign ap_ST_fsm_state2_blk = 1'b0;

assign ap_ST_fsm_state30_blk = 1'b0;

assign ap_ST_fsm_state31_blk = 1'b0;

assign ap_ST_fsm_state32_blk = 1'b0;

assign ap_ST_fsm_state33_blk = 1'b0;

assign ap_ST_fsm_state34_blk = 1'b0;

assign ap_ST_fsm_state35_blk = 1'b0;

assign ap_ST_fsm_state36_blk = 1'b0;

assign ap_ST_fsm_state37_blk = 1'b0;

assign ap_ST_fsm_state38_blk = 1'b0;

assign ap_ST_fsm_state39_blk = 1'b0;

always @ (*) begin
    if ((1'b1 == ap_block_state3_on_subcall_done)) begin
        ap_ST_fsm_state3_blk = 1'b1;
    end else begin
        ap_ST_fsm_state3_blk = 1'b0;
    end
end

assign ap_ST_fsm_state40_blk = 1'b0;

assign ap_ST_fsm_state41_blk = 1'b0;

assign ap_ST_fsm_state42_blk = 1'b0;

assign ap_ST_fsm_state43_blk = 1'b0;

assign ap_ST_fsm_state44_blk = 1'b0;

assign ap_ST_fsm_state45_blk = 1'b0;

assign ap_ST_fsm_state46_blk = 1'b0;

assign ap_ST_fsm_state47_blk = 1'b0;

assign ap_ST_fsm_state48_blk = 1'b0;

assign ap_ST_fsm_state49_blk = 1'b0;

assign ap_ST_fsm_state4_blk = 1'b0;

assign ap_ST_fsm_state50_blk = 1'b0;

assign ap_ST_fsm_state51_blk = 1'b0;

assign ap_ST_fsm_state52_blk = 1'b0;

assign ap_ST_fsm_state53_blk = 1'b0;

assign ap_ST_fsm_state54_blk = 1'b0;

assign ap_ST_fsm_state55_blk = 1'b0;

assign ap_ST_fsm_state56_blk = 1'b0;

assign ap_ST_fsm_state57_blk = 1'b0;

assign ap_ST_fsm_state58_blk = 1'b0;

assign ap_ST_fsm_state59_blk = 1'b0;

always @ (*) begin
    if ((grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_ap_done == 1'b0)) begin
        ap_ST_fsm_state5_blk = 1'b1;
    end else begin
        ap_ST_fsm_state5_blk = 1'b0;
    end
end

assign ap_ST_fsm_state60_blk = 1'b0;

assign ap_ST_fsm_state61_blk = 1'b0;

assign ap_ST_fsm_state62_blk = 1'b0;

assign ap_ST_fsm_state63_blk = 1'b0;

assign ap_ST_fsm_state64_blk = 1'b0;

assign ap_ST_fsm_state65_blk = 1'b0;

assign ap_ST_fsm_state66_blk = 1'b0;

assign ap_ST_fsm_state67_blk = 1'b0;

assign ap_ST_fsm_state68_blk = 1'b0;

assign ap_ST_fsm_state69_blk = 1'b0;

assign ap_ST_fsm_state6_blk = 1'b0;

assign ap_ST_fsm_state70_blk = 1'b0;

assign ap_ST_fsm_state71_blk = 1'b0;

assign ap_ST_fsm_state72_blk = 1'b0;

assign ap_ST_fsm_state73_blk = 1'b0;

assign ap_ST_fsm_state74_blk = 1'b0;

assign ap_ST_fsm_state75_blk = 1'b0;

assign ap_ST_fsm_state76_blk = 1'b0;

assign ap_ST_fsm_state77_blk = 1'b0;

assign ap_ST_fsm_state78_blk = 1'b0;

assign ap_ST_fsm_state79_blk = 1'b0;

assign ap_ST_fsm_state7_blk = 1'b0;

assign ap_ST_fsm_state80_blk = 1'b0;

assign ap_ST_fsm_state81_blk = 1'b0;

assign ap_ST_fsm_state82_blk = 1'b0;

assign ap_ST_fsm_state83_blk = 1'b0;

assign ap_ST_fsm_state84_blk = 1'b0;

assign ap_ST_fsm_state85_blk = 1'b0;

assign ap_ST_fsm_state86_blk = 1'b0;

assign ap_ST_fsm_state87_blk = 1'b0;

assign ap_ST_fsm_state88_blk = 1'b0;

assign ap_ST_fsm_state89_blk = 1'b0;

assign ap_ST_fsm_state8_blk = 1'b0;

assign ap_ST_fsm_state90_blk = 1'b0;

assign ap_ST_fsm_state91_blk = 1'b0;

assign ap_ST_fsm_state92_blk = 1'b0;

assign ap_ST_fsm_state93_blk = 1'b0;

assign ap_ST_fsm_state94_blk = 1'b0;

assign ap_ST_fsm_state95_blk = 1'b0;

assign ap_ST_fsm_state96_blk = 1'b0;

assign ap_ST_fsm_state97_blk = 1'b0;

assign ap_ST_fsm_state98_blk = 1'b0;

assign ap_ST_fsm_state99_blk = 1'b0;

assign ap_ST_fsm_state9_blk = 1'b0;

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state150) | ((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0)))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state150)) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state150)) begin
        ap_return = converged_0_lcssa_reg_319;
    end else begin
        ap_return = ap_return_preg;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state77)) begin
        centroid_x_coords_address0 = zext_ln101_reg_683;
    end else if (((cmp165_reg_628 == 1'd1) & (1'b1 == ap_CS_fsm_state148))) begin
        centroid_x_coords_address0 = grp_kmeans_Pipeline_VITIS_LOOP_116_6_fu_373_centroid_x_coords_address0;
    end else if ((1'b1 == ap_CS_fsm_state5)) begin
        centroid_x_coords_address0 = grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_centroid_x_coords_address0;
    end else if (((empty_76_reg_619 == 1'd0) & (1'b1 == ap_CS_fsm_state3))) begin
        centroid_x_coords_address0 = grp_kmeans_Pipeline_1_fu_332_centroid_x_coords_address0;
    end else begin
        centroid_x_coords_address0 = 'bx;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state77)) begin
        centroid_x_coords_ce0 = 1'b1;
    end else if (((cmp165_reg_628 == 1'd1) & (1'b1 == ap_CS_fsm_state148))) begin
        centroid_x_coords_ce0 = grp_kmeans_Pipeline_VITIS_LOOP_116_6_fu_373_centroid_x_coords_ce0;
    end else if ((1'b1 == ap_CS_fsm_state5)) begin
        centroid_x_coords_ce0 = grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_centroid_x_coords_ce0;
    end else if (((empty_76_reg_619 == 1'd0) & (1'b1 == ap_CS_fsm_state3))) begin
        centroid_x_coords_ce0 = grp_kmeans_Pipeline_1_fu_332_centroid_x_coords_ce0;
    end else begin
        centroid_x_coords_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state5)) begin
        centroid_x_coords_ce1 = grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_centroid_x_coords_ce1;
    end else begin
        centroid_x_coords_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state9)) begin
        centroid_x_coords_next_address0 = zext_ln101_reg_683;
    end else if ((1'b1 == ap_CS_fsm_state7)) begin
        centroid_x_coords_next_address0 = centroid_x_coords_next_addr_reg_663;
    end else if ((1'b1 == ap_CS_fsm_state6)) begin
        centroid_x_coords_next_address0 = sext_ln94_fu_479_p1;
    end else if (((empty_76_reg_619 == 1'd0) & (1'b1 == ap_CS_fsm_state3))) begin
        centroid_x_coords_next_address0 = grp_kmeans_Pipeline_3_fu_346_centroid_x_coords_next_address0;
    end else begin
        centroid_x_coords_next_address0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state6) | (1'b1 == ap_CS_fsm_state9))) begin
        centroid_x_coords_next_ce0 = 1'b1;
    end else if (((empty_76_reg_619 == 1'd0) & (1'b1 == ap_CS_fsm_state3))) begin
        centroid_x_coords_next_ce0 = grp_kmeans_Pipeline_3_fu_346_centroid_x_coords_next_ce0;
    end else begin
        centroid_x_coords_next_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state7)) begin
        centroid_x_coords_next_d0 = add_ln95_fu_487_p2;
    end else if (((empty_76_reg_619 == 1'd0) & (1'b1 == ap_CS_fsm_state3))) begin
        centroid_x_coords_next_d0 = grp_kmeans_Pipeline_3_fu_346_centroid_x_coords_next_d0;
    end else begin
        centroid_x_coords_next_d0 = 'bx;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state7)) begin
        centroid_x_coords_next_we0 = 1'b1;
    end else if (((empty_76_reg_619 == 1'd0) & (1'b1 == ap_CS_fsm_state3))) begin
        centroid_x_coords_next_we0 = grp_kmeans_Pipeline_3_fu_346_centroid_x_coords_next_we0;
    end else begin
        centroid_x_coords_next_we0 = 1'b0;
    end
end

always @ (*) begin
    if (((cmp165_reg_628 == 1'd1) & (1'b1 == ap_CS_fsm_state148))) begin
        centroid_x_coords_prev_address0 = grp_kmeans_Pipeline_VITIS_LOOP_116_6_fu_373_centroid_x_coords_prev_address0;
    end else if (((empty_76_reg_619 == 1'd0) & (1'b1 == ap_CS_fsm_state3))) begin
        centroid_x_coords_prev_address0 = grp_kmeans_Pipeline_1_fu_332_centroid_x_coords_prev_address0;
    end else begin
        centroid_x_coords_prev_address0 = 'bx;
    end
end

always @ (*) begin
    if (((cmp165_reg_628 == 1'd1) & (1'b1 == ap_CS_fsm_state148))) begin
        centroid_x_coords_prev_ce0 = grp_kmeans_Pipeline_VITIS_LOOP_116_6_fu_373_centroid_x_coords_prev_ce0;
    end else if (((empty_76_reg_619 == 1'd0) & (1'b1 == ap_CS_fsm_state3))) begin
        centroid_x_coords_prev_ce0 = grp_kmeans_Pipeline_1_fu_332_centroid_x_coords_prev_ce0;
    end else begin
        centroid_x_coords_prev_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((empty_76_reg_619 == 1'd0) & (1'b1 == ap_CS_fsm_state3))) begin
        centroid_x_coords_prev_we0 = grp_kmeans_Pipeline_1_fu_332_centroid_x_coords_prev_we0;
    end else begin
        centroid_x_coords_prev_we0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln103_reg_697 == 1'd0) & (1'b1 == ap_CS_fsm_state77))) begin
        centroid_x_coords_we0 = 1'b1;
    end else begin
        centroid_x_coords_we0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state147)) begin
        centroid_y_coords_address0 = zext_ln107_reg_721;
    end else if (((cmp165_reg_628 == 1'd1) & (1'b1 == ap_CS_fsm_state148))) begin
        centroid_y_coords_address0 = grp_kmeans_Pipeline_VITIS_LOOP_116_6_fu_373_centroid_y_coords_address0;
    end else if ((1'b1 == ap_CS_fsm_state5)) begin
        centroid_y_coords_address0 = grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_centroid_y_coords_address0;
    end else begin
        centroid_y_coords_address0 = 'bx;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state147)) begin
        centroid_y_coords_ce0 = 1'b1;
    end else if (((cmp165_reg_628 == 1'd1) & (1'b1 == ap_CS_fsm_state148))) begin
        centroid_y_coords_ce0 = grp_kmeans_Pipeline_VITIS_LOOP_116_6_fu_373_centroid_y_coords_ce0;
    end else if ((1'b1 == ap_CS_fsm_state5)) begin
        centroid_y_coords_ce0 = grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_centroid_y_coords_ce0;
    end else begin
        centroid_y_coords_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state5)) begin
        centroid_y_coords_ce1 = grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_centroid_y_coords_ce1;
    end else begin
        centroid_y_coords_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state79)) begin
        centroid_y_coords_next_address0 = zext_ln107_reg_721;
    end else if ((1'b1 == ap_CS_fsm_state7)) begin
        centroid_y_coords_next_address0 = centroid_y_coords_next_addr_reg_668;
    end else if ((1'b1 == ap_CS_fsm_state6)) begin
        centroid_y_coords_next_address0 = sext_ln94_fu_479_p1;
    end else if (((empty_76_reg_619 == 1'd0) & (1'b1 == ap_CS_fsm_state3))) begin
        centroid_y_coords_next_address0 = grp_kmeans_Pipeline_4_fu_352_centroid_y_coords_next_address0;
    end else begin
        centroid_y_coords_next_address0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state6) | (1'b1 == ap_CS_fsm_state79))) begin
        centroid_y_coords_next_ce0 = 1'b1;
    end else if (((empty_76_reg_619 == 1'd0) & (1'b1 == ap_CS_fsm_state3))) begin
        centroid_y_coords_next_ce0 = grp_kmeans_Pipeline_4_fu_352_centroid_y_coords_next_ce0;
    end else begin
        centroid_y_coords_next_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state7)) begin
        centroid_y_coords_next_d0 = add_ln96_fu_494_p2;
    end else if (((empty_76_reg_619 == 1'd0) & (1'b1 == ap_CS_fsm_state3))) begin
        centroid_y_coords_next_d0 = grp_kmeans_Pipeline_4_fu_352_centroid_y_coords_next_d0;
    end else begin
        centroid_y_coords_next_d0 = 'bx;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state7)) begin
        centroid_y_coords_next_we0 = 1'b1;
    end else if (((empty_76_reg_619 == 1'd0) & (1'b1 == ap_CS_fsm_state3))) begin
        centroid_y_coords_next_we0 = grp_kmeans_Pipeline_4_fu_352_centroid_y_coords_next_we0;
    end else begin
        centroid_y_coords_next_we0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln109_reg_735 == 1'd0) & (1'b1 == ap_CS_fsm_state147))) begin
        centroid_y_coords_we0 = 1'b1;
    end else begin
        centroid_y_coords_we0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state78)) begin
        cluster_cardinality_next_address0 = zext_ln107_fu_545_p1;
    end else if ((1'b1 == ap_CS_fsm_state8)) begin
        cluster_cardinality_next_address0 = zext_ln101_fu_514_p1;
    end else if ((1'b1 == ap_CS_fsm_state7)) begin
        cluster_cardinality_next_address0 = cluster_cardinality_next_addr_reg_673;
    end else if ((1'b1 == ap_CS_fsm_state6)) begin
        cluster_cardinality_next_address0 = sext_ln94_fu_479_p1;
    end else if (((empty_76_reg_619 == 1'd0) & (1'b1 == ap_CS_fsm_state3))) begin
        cluster_cardinality_next_address0 = grp_kmeans_Pipeline_2_fu_340_cluster_cardinality_next_address0;
    end else begin
        cluster_cardinality_next_address0 = 'bx;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state78) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state6))) begin
        cluster_cardinality_next_ce0 = 1'b1;
    end else if (((empty_76_reg_619 == 1'd0) & (1'b1 == ap_CS_fsm_state3))) begin
        cluster_cardinality_next_ce0 = grp_kmeans_Pipeline_2_fu_340_cluster_cardinality_next_ce0;
    end else begin
        cluster_cardinality_next_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state7)) begin
        cluster_cardinality_next_d0 = add_ln97_fu_501_p2;
    end else if (((empty_76_reg_619 == 1'd0) & (1'b1 == ap_CS_fsm_state3))) begin
        cluster_cardinality_next_d0 = grp_kmeans_Pipeline_2_fu_340_cluster_cardinality_next_d0;
    end else begin
        cluster_cardinality_next_d0 = 'bx;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state7)) begin
        cluster_cardinality_next_we0 = 1'b1;
    end else if (((empty_76_reg_619 == 1'd0) & (1'b1 == ap_CS_fsm_state3))) begin
        cluster_cardinality_next_we0 = grp_kmeans_Pipeline_2_fu_340_cluster_cardinality_next_we0;
    end else begin
        cluster_cardinality_next_we0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state10)) begin
        grp_fu_532_ap_start = 1'b1;
    end else begin
        grp_fu_532_ap_start = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state80)) begin
        grp_fu_563_ap_start = 1'b1;
    end else begin
        grp_fu_563_ap_start = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state6)) begin
        node_cluster_assignments_ce1 = 1'b1;
    end else begin
        node_cluster_assignments_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state6)) begin
        node_cluster_assignments_we1 = 1'b1;
    end else begin
        node_cluster_assignments_we1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state6)) begin
        node_x_coords_address0 = zext_ln69_fu_469_p1;
    end else if ((1'b1 == ap_CS_fsm_state5)) begin
        node_x_coords_address0 = grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_node_x_coords_address0;
    end else begin
        node_x_coords_address0 = 'bx;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state6)) begin
        node_x_coords_ce0 = 1'b1;
    end else if ((1'b1 == ap_CS_fsm_state5)) begin
        node_x_coords_ce0 = grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_node_x_coords_ce0;
    end else begin
        node_x_coords_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state5)) begin
        node_x_coords_ce1 = grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_node_x_coords_ce1;
    end else begin
        node_x_coords_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state6)) begin
        node_y_coords_address0 = zext_ln69_fu_469_p1;
    end else if ((1'b1 == ap_CS_fsm_state5)) begin
        node_y_coords_address0 = grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_node_y_coords_address0;
    end else begin
        node_y_coords_address0 = 'bx;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state6)) begin
        node_y_coords_ce0 = 1'b1;
    end else if ((1'b1 == ap_CS_fsm_state5)) begin
        node_y_coords_ce0 = grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_node_y_coords_ce0;
    end else begin
        node_y_coords_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state5)) begin
        node_y_coords_ce1 = grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_node_y_coords_ce1;
    end else begin
        node_y_coords_ce1 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            if (((icmp_ln53_fu_443_p2 == 1'd1) & (ap_phi_mux_converged_phi_fu_263_p4 == 1'd0) & (1'b1 == ap_CS_fsm_state2))) begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state150;
            end
        end
        ap_ST_fsm_state3 : begin
            if (((1'b0 == ap_block_state3_on_subcall_done) & (1'b1 == ap_CS_fsm_state3))) begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
        end
        ap_ST_fsm_state4 : begin
            if (((icmp_ln69_fu_459_p2 == 1'd0) & (cmp165_reg_628 == 1'd1) & (1'b1 == ap_CS_fsm_state4))) begin
                ap_NS_fsm = ap_ST_fsm_state8;
            end else if (((icmp_ln69_fu_459_p2 == 1'd0) & (cmp165_reg_628 == 1'd0) & (1'b1 == ap_CS_fsm_state4))) begin
                ap_NS_fsm = ap_ST_fsm_state148;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state5;
            end
        end
        ap_ST_fsm_state5 : begin
            if (((grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state5))) begin
                ap_NS_fsm = ap_ST_fsm_state6;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state5;
            end
        end
        ap_ST_fsm_state6 : begin
            ap_NS_fsm = ap_ST_fsm_state7;
        end
        ap_ST_fsm_state7 : begin
            ap_NS_fsm = ap_ST_fsm_state4;
        end
        ap_ST_fsm_state8 : begin
            if (((icmp_ln101_fu_523_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state8))) begin
                ap_NS_fsm = ap_ST_fsm_state78;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state9;
            end
        end
        ap_ST_fsm_state9 : begin
            if (((grp_fu_383_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state9))) begin
                ap_NS_fsm = ap_ST_fsm_state77;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state10;
            end
        end
        ap_ST_fsm_state10 : begin
            ap_NS_fsm = ap_ST_fsm_state11;
        end
        ap_ST_fsm_state11 : begin
            ap_NS_fsm = ap_ST_fsm_state12;
        end
        ap_ST_fsm_state12 : begin
            ap_NS_fsm = ap_ST_fsm_state13;
        end
        ap_ST_fsm_state13 : begin
            ap_NS_fsm = ap_ST_fsm_state14;
        end
        ap_ST_fsm_state14 : begin
            ap_NS_fsm = ap_ST_fsm_state15;
        end
        ap_ST_fsm_state15 : begin
            ap_NS_fsm = ap_ST_fsm_state16;
        end
        ap_ST_fsm_state16 : begin
            ap_NS_fsm = ap_ST_fsm_state17;
        end
        ap_ST_fsm_state17 : begin
            ap_NS_fsm = ap_ST_fsm_state18;
        end
        ap_ST_fsm_state18 : begin
            ap_NS_fsm = ap_ST_fsm_state19;
        end
        ap_ST_fsm_state19 : begin
            ap_NS_fsm = ap_ST_fsm_state20;
        end
        ap_ST_fsm_state20 : begin
            ap_NS_fsm = ap_ST_fsm_state21;
        end
        ap_ST_fsm_state21 : begin
            ap_NS_fsm = ap_ST_fsm_state22;
        end
        ap_ST_fsm_state22 : begin
            ap_NS_fsm = ap_ST_fsm_state23;
        end
        ap_ST_fsm_state23 : begin
            ap_NS_fsm = ap_ST_fsm_state24;
        end
        ap_ST_fsm_state24 : begin
            ap_NS_fsm = ap_ST_fsm_state25;
        end
        ap_ST_fsm_state25 : begin
            ap_NS_fsm = ap_ST_fsm_state26;
        end
        ap_ST_fsm_state26 : begin
            ap_NS_fsm = ap_ST_fsm_state27;
        end
        ap_ST_fsm_state27 : begin
            ap_NS_fsm = ap_ST_fsm_state28;
        end
        ap_ST_fsm_state28 : begin
            ap_NS_fsm = ap_ST_fsm_state29;
        end
        ap_ST_fsm_state29 : begin
            ap_NS_fsm = ap_ST_fsm_state30;
        end
        ap_ST_fsm_state30 : begin
            ap_NS_fsm = ap_ST_fsm_state31;
        end
        ap_ST_fsm_state31 : begin
            ap_NS_fsm = ap_ST_fsm_state32;
        end
        ap_ST_fsm_state32 : begin
            ap_NS_fsm = ap_ST_fsm_state33;
        end
        ap_ST_fsm_state33 : begin
            ap_NS_fsm = ap_ST_fsm_state34;
        end
        ap_ST_fsm_state34 : begin
            ap_NS_fsm = ap_ST_fsm_state35;
        end
        ap_ST_fsm_state35 : begin
            ap_NS_fsm = ap_ST_fsm_state36;
        end
        ap_ST_fsm_state36 : begin
            ap_NS_fsm = ap_ST_fsm_state37;
        end
        ap_ST_fsm_state37 : begin
            ap_NS_fsm = ap_ST_fsm_state38;
        end
        ap_ST_fsm_state38 : begin
            ap_NS_fsm = ap_ST_fsm_state39;
        end
        ap_ST_fsm_state39 : begin
            ap_NS_fsm = ap_ST_fsm_state40;
        end
        ap_ST_fsm_state40 : begin
            ap_NS_fsm = ap_ST_fsm_state41;
        end
        ap_ST_fsm_state41 : begin
            ap_NS_fsm = ap_ST_fsm_state42;
        end
        ap_ST_fsm_state42 : begin
            ap_NS_fsm = ap_ST_fsm_state43;
        end
        ap_ST_fsm_state43 : begin
            ap_NS_fsm = ap_ST_fsm_state44;
        end
        ap_ST_fsm_state44 : begin
            ap_NS_fsm = ap_ST_fsm_state45;
        end
        ap_ST_fsm_state45 : begin
            ap_NS_fsm = ap_ST_fsm_state46;
        end
        ap_ST_fsm_state46 : begin
            ap_NS_fsm = ap_ST_fsm_state47;
        end
        ap_ST_fsm_state47 : begin
            ap_NS_fsm = ap_ST_fsm_state48;
        end
        ap_ST_fsm_state48 : begin
            ap_NS_fsm = ap_ST_fsm_state49;
        end
        ap_ST_fsm_state49 : begin
            ap_NS_fsm = ap_ST_fsm_state50;
        end
        ap_ST_fsm_state50 : begin
            ap_NS_fsm = ap_ST_fsm_state51;
        end
        ap_ST_fsm_state51 : begin
            ap_NS_fsm = ap_ST_fsm_state52;
        end
        ap_ST_fsm_state52 : begin
            ap_NS_fsm = ap_ST_fsm_state53;
        end
        ap_ST_fsm_state53 : begin
            ap_NS_fsm = ap_ST_fsm_state54;
        end
        ap_ST_fsm_state54 : begin
            ap_NS_fsm = ap_ST_fsm_state55;
        end
        ap_ST_fsm_state55 : begin
            ap_NS_fsm = ap_ST_fsm_state56;
        end
        ap_ST_fsm_state56 : begin
            ap_NS_fsm = ap_ST_fsm_state57;
        end
        ap_ST_fsm_state57 : begin
            ap_NS_fsm = ap_ST_fsm_state58;
        end
        ap_ST_fsm_state58 : begin
            ap_NS_fsm = ap_ST_fsm_state59;
        end
        ap_ST_fsm_state59 : begin
            ap_NS_fsm = ap_ST_fsm_state60;
        end
        ap_ST_fsm_state60 : begin
            ap_NS_fsm = ap_ST_fsm_state61;
        end
        ap_ST_fsm_state61 : begin
            ap_NS_fsm = ap_ST_fsm_state62;
        end
        ap_ST_fsm_state62 : begin
            ap_NS_fsm = ap_ST_fsm_state63;
        end
        ap_ST_fsm_state63 : begin
            ap_NS_fsm = ap_ST_fsm_state64;
        end
        ap_ST_fsm_state64 : begin
            ap_NS_fsm = ap_ST_fsm_state65;
        end
        ap_ST_fsm_state65 : begin
            ap_NS_fsm = ap_ST_fsm_state66;
        end
        ap_ST_fsm_state66 : begin
            ap_NS_fsm = ap_ST_fsm_state67;
        end
        ap_ST_fsm_state67 : begin
            ap_NS_fsm = ap_ST_fsm_state68;
        end
        ap_ST_fsm_state68 : begin
            ap_NS_fsm = ap_ST_fsm_state69;
        end
        ap_ST_fsm_state69 : begin
            ap_NS_fsm = ap_ST_fsm_state70;
        end
        ap_ST_fsm_state70 : begin
            ap_NS_fsm = ap_ST_fsm_state71;
        end
        ap_ST_fsm_state71 : begin
            ap_NS_fsm = ap_ST_fsm_state72;
        end
        ap_ST_fsm_state72 : begin
            ap_NS_fsm = ap_ST_fsm_state73;
        end
        ap_ST_fsm_state73 : begin
            ap_NS_fsm = ap_ST_fsm_state74;
        end
        ap_ST_fsm_state74 : begin
            ap_NS_fsm = ap_ST_fsm_state75;
        end
        ap_ST_fsm_state75 : begin
            ap_NS_fsm = ap_ST_fsm_state76;
        end
        ap_ST_fsm_state76 : begin
            ap_NS_fsm = ap_ST_fsm_state77;
        end
        ap_ST_fsm_state77 : begin
            ap_NS_fsm = ap_ST_fsm_state8;
        end
        ap_ST_fsm_state78 : begin
            if (((icmp_ln107_fu_554_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state78))) begin
                ap_NS_fsm = ap_ST_fsm_state148;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state79;
            end
        end
        ap_ST_fsm_state79 : begin
            if (((grp_fu_383_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state79))) begin
                ap_NS_fsm = ap_ST_fsm_state147;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state80;
            end
        end
        ap_ST_fsm_state80 : begin
            ap_NS_fsm = ap_ST_fsm_state81;
        end
        ap_ST_fsm_state81 : begin
            ap_NS_fsm = ap_ST_fsm_state82;
        end
        ap_ST_fsm_state82 : begin
            ap_NS_fsm = ap_ST_fsm_state83;
        end
        ap_ST_fsm_state83 : begin
            ap_NS_fsm = ap_ST_fsm_state84;
        end
        ap_ST_fsm_state84 : begin
            ap_NS_fsm = ap_ST_fsm_state85;
        end
        ap_ST_fsm_state85 : begin
            ap_NS_fsm = ap_ST_fsm_state86;
        end
        ap_ST_fsm_state86 : begin
            ap_NS_fsm = ap_ST_fsm_state87;
        end
        ap_ST_fsm_state87 : begin
            ap_NS_fsm = ap_ST_fsm_state88;
        end
        ap_ST_fsm_state88 : begin
            ap_NS_fsm = ap_ST_fsm_state89;
        end
        ap_ST_fsm_state89 : begin
            ap_NS_fsm = ap_ST_fsm_state90;
        end
        ap_ST_fsm_state90 : begin
            ap_NS_fsm = ap_ST_fsm_state91;
        end
        ap_ST_fsm_state91 : begin
            ap_NS_fsm = ap_ST_fsm_state92;
        end
        ap_ST_fsm_state92 : begin
            ap_NS_fsm = ap_ST_fsm_state93;
        end
        ap_ST_fsm_state93 : begin
            ap_NS_fsm = ap_ST_fsm_state94;
        end
        ap_ST_fsm_state94 : begin
            ap_NS_fsm = ap_ST_fsm_state95;
        end
        ap_ST_fsm_state95 : begin
            ap_NS_fsm = ap_ST_fsm_state96;
        end
        ap_ST_fsm_state96 : begin
            ap_NS_fsm = ap_ST_fsm_state97;
        end
        ap_ST_fsm_state97 : begin
            ap_NS_fsm = ap_ST_fsm_state98;
        end
        ap_ST_fsm_state98 : begin
            ap_NS_fsm = ap_ST_fsm_state99;
        end
        ap_ST_fsm_state99 : begin
            ap_NS_fsm = ap_ST_fsm_state100;
        end
        ap_ST_fsm_state100 : begin
            ap_NS_fsm = ap_ST_fsm_state101;
        end
        ap_ST_fsm_state101 : begin
            ap_NS_fsm = ap_ST_fsm_state102;
        end
        ap_ST_fsm_state102 : begin
            ap_NS_fsm = ap_ST_fsm_state103;
        end
        ap_ST_fsm_state103 : begin
            ap_NS_fsm = ap_ST_fsm_state104;
        end
        ap_ST_fsm_state104 : begin
            ap_NS_fsm = ap_ST_fsm_state105;
        end
        ap_ST_fsm_state105 : begin
            ap_NS_fsm = ap_ST_fsm_state106;
        end
        ap_ST_fsm_state106 : begin
            ap_NS_fsm = ap_ST_fsm_state107;
        end
        ap_ST_fsm_state107 : begin
            ap_NS_fsm = ap_ST_fsm_state108;
        end
        ap_ST_fsm_state108 : begin
            ap_NS_fsm = ap_ST_fsm_state109;
        end
        ap_ST_fsm_state109 : begin
            ap_NS_fsm = ap_ST_fsm_state110;
        end
        ap_ST_fsm_state110 : begin
            ap_NS_fsm = ap_ST_fsm_state111;
        end
        ap_ST_fsm_state111 : begin
            ap_NS_fsm = ap_ST_fsm_state112;
        end
        ap_ST_fsm_state112 : begin
            ap_NS_fsm = ap_ST_fsm_state113;
        end
        ap_ST_fsm_state113 : begin
            ap_NS_fsm = ap_ST_fsm_state114;
        end
        ap_ST_fsm_state114 : begin
            ap_NS_fsm = ap_ST_fsm_state115;
        end
        ap_ST_fsm_state115 : begin
            ap_NS_fsm = ap_ST_fsm_state116;
        end
        ap_ST_fsm_state116 : begin
            ap_NS_fsm = ap_ST_fsm_state117;
        end
        ap_ST_fsm_state117 : begin
            ap_NS_fsm = ap_ST_fsm_state118;
        end
        ap_ST_fsm_state118 : begin
            ap_NS_fsm = ap_ST_fsm_state119;
        end
        ap_ST_fsm_state119 : begin
            ap_NS_fsm = ap_ST_fsm_state120;
        end
        ap_ST_fsm_state120 : begin
            ap_NS_fsm = ap_ST_fsm_state121;
        end
        ap_ST_fsm_state121 : begin
            ap_NS_fsm = ap_ST_fsm_state122;
        end
        ap_ST_fsm_state122 : begin
            ap_NS_fsm = ap_ST_fsm_state123;
        end
        ap_ST_fsm_state123 : begin
            ap_NS_fsm = ap_ST_fsm_state124;
        end
        ap_ST_fsm_state124 : begin
            ap_NS_fsm = ap_ST_fsm_state125;
        end
        ap_ST_fsm_state125 : begin
            ap_NS_fsm = ap_ST_fsm_state126;
        end
        ap_ST_fsm_state126 : begin
            ap_NS_fsm = ap_ST_fsm_state127;
        end
        ap_ST_fsm_state127 : begin
            ap_NS_fsm = ap_ST_fsm_state128;
        end
        ap_ST_fsm_state128 : begin
            ap_NS_fsm = ap_ST_fsm_state129;
        end
        ap_ST_fsm_state129 : begin
            ap_NS_fsm = ap_ST_fsm_state130;
        end
        ap_ST_fsm_state130 : begin
            ap_NS_fsm = ap_ST_fsm_state131;
        end
        ap_ST_fsm_state131 : begin
            ap_NS_fsm = ap_ST_fsm_state132;
        end
        ap_ST_fsm_state132 : begin
            ap_NS_fsm = ap_ST_fsm_state133;
        end
        ap_ST_fsm_state133 : begin
            ap_NS_fsm = ap_ST_fsm_state134;
        end
        ap_ST_fsm_state134 : begin
            ap_NS_fsm = ap_ST_fsm_state135;
        end
        ap_ST_fsm_state135 : begin
            ap_NS_fsm = ap_ST_fsm_state136;
        end
        ap_ST_fsm_state136 : begin
            ap_NS_fsm = ap_ST_fsm_state137;
        end
        ap_ST_fsm_state137 : begin
            ap_NS_fsm = ap_ST_fsm_state138;
        end
        ap_ST_fsm_state138 : begin
            ap_NS_fsm = ap_ST_fsm_state139;
        end
        ap_ST_fsm_state139 : begin
            ap_NS_fsm = ap_ST_fsm_state140;
        end
        ap_ST_fsm_state140 : begin
            ap_NS_fsm = ap_ST_fsm_state141;
        end
        ap_ST_fsm_state141 : begin
            ap_NS_fsm = ap_ST_fsm_state142;
        end
        ap_ST_fsm_state142 : begin
            ap_NS_fsm = ap_ST_fsm_state143;
        end
        ap_ST_fsm_state143 : begin
            ap_NS_fsm = ap_ST_fsm_state144;
        end
        ap_ST_fsm_state144 : begin
            ap_NS_fsm = ap_ST_fsm_state145;
        end
        ap_ST_fsm_state145 : begin
            ap_NS_fsm = ap_ST_fsm_state146;
        end
        ap_ST_fsm_state146 : begin
            ap_NS_fsm = ap_ST_fsm_state147;
        end
        ap_ST_fsm_state147 : begin
            ap_NS_fsm = ap_ST_fsm_state78;
        end
        ap_ST_fsm_state148 : begin
            if (((1'b0 == ap_block_state148_on_subcall_done) & (1'b1 == ap_CS_fsm_state148))) begin
                ap_NS_fsm = ap_ST_fsm_state149;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state148;
            end
        end
        ap_ST_fsm_state149 : begin
            ap_NS_fsm = ap_ST_fsm_state2;
        end
        ap_ST_fsm_state150 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln101_fu_508_p2 = (i_1_reg_282 + 31'd1);

assign add_ln107_fu_539_p2 = (i_2_reg_293 + 31'd1);

assign add_ln69_fu_449_p2 = (i_reg_270 + 14'd1);

assign add_ln95_fu_487_p2 = (centroid_x_coords_next_q0 + node_x_coords_q0);

assign add_ln96_fu_494_p2 = (centroid_y_coords_next_q0 + node_y_coords_q0);

assign add_ln97_fu_501_p2 = (cluster_cardinality_next_q0 + 16'd1);

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state10 = ap_CS_fsm[32'd9];

assign ap_CS_fsm_state147 = ap_CS_fsm[32'd146];

assign ap_CS_fsm_state148 = ap_CS_fsm[32'd147];

assign ap_CS_fsm_state149 = ap_CS_fsm[32'd148];

assign ap_CS_fsm_state150 = ap_CS_fsm[32'd149];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

assign ap_CS_fsm_state5 = ap_CS_fsm[32'd4];

assign ap_CS_fsm_state6 = ap_CS_fsm[32'd5];

assign ap_CS_fsm_state7 = ap_CS_fsm[32'd6];

assign ap_CS_fsm_state77 = ap_CS_fsm[32'd76];

assign ap_CS_fsm_state78 = ap_CS_fsm[32'd77];

assign ap_CS_fsm_state79 = ap_CS_fsm[32'd78];

assign ap_CS_fsm_state8 = ap_CS_fsm[32'd7];

assign ap_CS_fsm_state80 = ap_CS_fsm[32'd79];

assign ap_CS_fsm_state9 = ap_CS_fsm[32'd8];

always @ (*) begin
    ap_block_state148_on_subcall_done = ((grp_kmeans_Pipeline_VITIS_LOOP_116_6_fu_373_ap_done == 1'b0) & (cmp165_reg_628 == 1'd1));
end

always @ (*) begin
    ap_block_state3_on_subcall_done = (((grp_kmeans_Pipeline_4_fu_352_ap_done == 1'b0) & (empty_76_reg_619 == 1'd0)) | ((grp_kmeans_Pipeline_3_fu_346_ap_done == 1'b0) & (empty_76_reg_619 == 1'd0)) | ((grp_kmeans_Pipeline_2_fu_340_ap_done == 1'b0) & (empty_76_reg_619 == 1'd0)) | ((grp_kmeans_Pipeline_1_fu_332_ap_done == 1'b0) & (empty_76_reg_619 == 1'd0)));
end

assign ap_phi_mux_converged_phi_fu_263_p4 = converged_reg_259;

assign centroid_x_coords_address1 = grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_centroid_x_coords_address1;

assign centroid_x_coords_d0 = grp_fu_532_p2;

assign centroid_y_coords_address1 = grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_centroid_y_coords_address1;

assign centroid_y_coords_d0 = grp_fu_563_p2;

assign cmp165_fu_416_p2 = (($signed(k) > $signed(32'd0)) ? 1'b1 : 1'b0);

assign cond_fu_570_p2 = ((grp_kmeans_Pipeline_VITIS_LOOP_116_6_fu_373_ap_return == 2'd0) ? 1'b1 : 1'b0);

assign current_iteration_3_fu_430_p2 = (current_iteration_fu_80 + 32'd1);

assign empty_76_fu_402_p2 = ((k == 32'd0) ? 1'b1 : 1'b0);

assign empty_fu_393_p1 = k[30:0];

assign grp_fu_383_p2 = ((cluster_cardinality_next_q0 == 16'd0) ? 1'b1 : 1'b0);

assign grp_fu_532_p1 = grp_fu_532_p10;

assign grp_fu_532_p10 = reg_389;

assign grp_fu_563_p1 = grp_fu_563_p10;

assign grp_fu_563_p10 = reg_389;

assign grp_kmeans_Pipeline_1_fu_332_ap_start = grp_kmeans_Pipeline_1_fu_332_ap_start_reg;

assign grp_kmeans_Pipeline_2_fu_340_ap_start = grp_kmeans_Pipeline_2_fu_340_ap_start_reg;

assign grp_kmeans_Pipeline_3_fu_346_ap_start = grp_kmeans_Pipeline_3_fu_346_ap_start_reg;

assign grp_kmeans_Pipeline_4_fu_352_ap_start = grp_kmeans_Pipeline_4_fu_352_ap_start_reg;

assign grp_kmeans_Pipeline_VITIS_LOOP_116_6_fu_373_ap_start = grp_kmeans_Pipeline_VITIS_LOOP_116_6_fu_373_ap_start_reg;

assign grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_ap_start = grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_ap_start_reg;

assign icmp_ln101_fu_523_p2 = ((zext_ln101_1_fu_519_p1 == k) ? 1'b1 : 1'b0);

assign icmp_ln107_fu_554_p2 = ((zext_ln107_1_fu_550_p1 == k) ? 1'b1 : 1'b0);

assign icmp_ln53_fu_443_p2 = ((max_iterations_assign_fu_88 > zext_ln53_fu_436_p1) ? 1'b1 : 1'b0);

assign icmp_ln69_fu_459_p2 = (($signed(zext_ln69_1_fu_455_p1) < $signed(n)) ? 1'b1 : 1'b0);

assign node_cluster_assignments_address1 = zext_ln69_fu_469_p1;

assign node_cluster_assignments_d1 = sext_ln94_fu_479_p1;

assign node_x_coords_address1 = grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_node_x_coords_address1;

assign node_y_coords_address1 = grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_node_y_coords_address1;

assign sext_ln94_fu_479_p1 = $signed(grp_kmeans_Pipeline_VITIS_LOOP_73_3_fu_358_min_dist_index_out);

assign tmp_fu_408_p3 = {{k}, {2'd0}};

assign trunc_ln37_fu_464_p1 = i_reg_270[12:0];

assign zext_ln101_1_fu_519_p1 = i_1_reg_282;

assign zext_ln101_fu_514_p1 = i_1_reg_282;

assign zext_ln107_1_fu_550_p1 = i_2_reg_293;

assign zext_ln107_fu_545_p1 = i_2_reg_293;

assign zext_ln53_fu_436_p1 = current_iteration_fu_80;

assign zext_ln69_1_fu_455_p1 = i_reg_270;

assign zext_ln69_fu_469_p1 = i_reg_270;

always @ (posedge ap_clk) begin
    tmp_reg_623[1:0] <= 2'b00;
    zext_ln101_reg_683[63:31] <= 33'b000000000000000000000000000000000;
    zext_ln107_reg_721[63:31] <= 33'b000000000000000000000000000000000;
end

endmodule //kmeans_top_kmeans


// Content from kmeans_top_kmeans_top_Pipeline_2.v
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2022.2 (64-bit)
// Version: 2022.2
// Copyright (C) Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module kmeans_top_kmeans_top_Pipeline_2 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        m_axi_mem_AWVALID,
        m_axi_mem_AWREADY,
        m_axi_mem_AWADDR,
        m_axi_mem_AWID,
        m_axi_mem_AWLEN,
        m_axi_mem_AWSIZE,
        m_axi_mem_AWBURST,
        m_axi_mem_AWLOCK,
        m_axi_mem_AWCACHE,
        m_axi_mem_AWPROT,
        m_axi_mem_AWQOS,
        m_axi_mem_AWREGION,
        m_axi_mem_AWUSER,
        m_axi_mem_WVALID,
        m_axi_mem_WREADY,
        m_axi_mem_WDATA,
        m_axi_mem_WSTRB,
        m_axi_mem_WLAST,
        m_axi_mem_WID,
        m_axi_mem_WUSER,
        m_axi_mem_ARVALID,
        m_axi_mem_ARREADY,
        m_axi_mem_ARADDR,
        m_axi_mem_ARID,
        m_axi_mem_ARLEN,
        m_axi_mem_ARSIZE,
        m_axi_mem_ARBURST,
        m_axi_mem_ARLOCK,
        m_axi_mem_ARCACHE,
        m_axi_mem_ARPROT,
        m_axi_mem_ARQOS,
        m_axi_mem_ARREGION,
        m_axi_mem_ARUSER,
        m_axi_mem_RVALID,
        m_axi_mem_RREADY,
        m_axi_mem_RDATA,
        m_axi_mem_RLAST,
        m_axi_mem_RID,
        m_axi_mem_RFIFONUM,
        m_axi_mem_RUSER,
        m_axi_mem_RRESP,
        m_axi_mem_BVALID,
        m_axi_mem_BREADY,
        m_axi_mem_BRESP,
        m_axi_mem_BID,
        m_axi_mem_BUSER,
        p_cast2_cast,
        node_y_coords_address1,
        node_y_coords_ce1,
        node_y_coords_we1,
        node_y_coords_d1,
        sext_ln182
);

parameter    ap_ST_fsm_pp0_stage0 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
output   m_axi_mem_AWVALID;
input   m_axi_mem_AWREADY;
output  [63:0] m_axi_mem_AWADDR;
output  [0:0] m_axi_mem_AWID;
output  [31:0] m_axi_mem_AWLEN;
output  [2:0] m_axi_mem_AWSIZE;
output  [1:0] m_axi_mem_AWBURST;
output  [1:0] m_axi_mem_AWLOCK;
output  [3:0] m_axi_mem_AWCACHE;
output  [2:0] m_axi_mem_AWPROT;
output  [3:0] m_axi_mem_AWQOS;
output  [3:0] m_axi_mem_AWREGION;
output  [0:0] m_axi_mem_AWUSER;
output   m_axi_mem_WVALID;
input   m_axi_mem_WREADY;
output  [63:0] m_axi_mem_WDATA;
output  [7:0] m_axi_mem_WSTRB;
output   m_axi_mem_WLAST;
output  [0:0] m_axi_mem_WID;
output  [0:0] m_axi_mem_WUSER;
output   m_axi_mem_ARVALID;
input   m_axi_mem_ARREADY;
output  [63:0] m_axi_mem_ARADDR;
output  [0:0] m_axi_mem_ARID;
output  [31:0] m_axi_mem_ARLEN;
output  [2:0] m_axi_mem_ARSIZE;
output  [1:0] m_axi_mem_ARBURST;
output  [1:0] m_axi_mem_ARLOCK;
output  [3:0] m_axi_mem_ARCACHE;
output  [2:0] m_axi_mem_ARPROT;
output  [3:0] m_axi_mem_ARQOS;
output  [3:0] m_axi_mem_ARREGION;
output  [0:0] m_axi_mem_ARUSER;
input   m_axi_mem_RVALID;
output   m_axi_mem_RREADY;
input  [63:0] m_axi_mem_RDATA;
input   m_axi_mem_RLAST;
input  [0:0] m_axi_mem_RID;
input  [8:0] m_axi_mem_RFIFONUM;
input  [0:0] m_axi_mem_RUSER;
input  [1:0] m_axi_mem_RRESP;
input   m_axi_mem_BVALID;
output   m_axi_mem_BREADY;
input  [1:0] m_axi_mem_BRESP;
input  [0:0] m_axi_mem_BID;
input  [0:0] m_axi_mem_BUSER;
input  [60:0] p_cast2_cast;
output  [12:0] node_y_coords_address1;
output   node_y_coords_ce1;
output   node_y_coords_we1;
output  [63:0] node_y_coords_d1;
input  [31:0] sext_ln182;

reg ap_idle;
reg m_axi_mem_RREADY;
reg node_y_coords_ce1;
reg node_y_coords_we1;

(* fsm_encoding = "none" *) reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_enable_reg_pp0_iter0;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter2;
reg    ap_idle_pp0;
wire    ap_block_state1_pp0_stage0_iter0;
reg    ap_block_state2_pp0_stage0_iter1;
wire    ap_block_state3_pp0_stage0_iter2;
reg    ap_block_pp0_stage0_subdone;
wire   [0:0] exitcond84_fu_126_p2;
reg    ap_condition_exit_pp0_iter1_stage0;
wire    ap_loop_exit_ready;
reg    ap_ready_int;
reg    mem_blk_n_R;
wire    ap_block_pp0_stage0;
wire  signed [60:0] sext_ln182_cast_fu_98_p1;
reg  signed [60:0] sext_ln182_cast_reg_147;
reg    ap_block_pp0_stage0_11001;
reg   [60:0] loop_index63_load_reg_157;
reg   [63:0] mem_addr_read_reg_162;
wire   [63:0] loop_index63_cast_fu_136_p1;
reg   [60:0] loop_index63_fu_60;
wire   [60:0] empty_fu_114_p2;
wire    ap_loop_init;
reg    ap_done_reg;
wire    ap_continue_int;
reg    ap_done_int;
reg    ap_loop_exit_ready_pp0_iter2_reg;
reg   [0:0] ap_NS_fsm;
wire    ap_enable_pp0;
wire    ap_start_int;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_CS_fsm = 1'd1;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_done_reg = 1'b0;
end

kmeans_top_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(ap_start),
    .ap_ready(ap_ready),
    .ap_done(ap_done),
    .ap_start_int(ap_start_int),
    .ap_loop_init(ap_loop_init),
    .ap_ready_int(ap_ready_int),
    .ap_loop_exit_ready(ap_condition_exit_pp0_iter1_stage0),
    .ap_loop_exit_done(ap_done_int),
    .ap_continue_int(ap_continue_int),
    .ap_done_int(ap_done_int)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue_int == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter2_reg == 1'b1))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b1 == ap_condition_exit_pp0_iter1_stage0)) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_enable_reg_pp0_iter1 <= ap_start_int;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready == 1'b0))) begin
        ap_loop_exit_ready_pp0_iter2_reg <= 1'b0;
    end else if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_loop_exit_ready_pp0_iter2_reg <= ap_loop_exit_ready;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        if ((ap_loop_init == 1'b1)) begin
            loop_index63_fu_60 <= 61'd0;
        end else if (((exitcond84_fu_126_p2 == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
            loop_index63_fu_60 <= empty_fu_114_p2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        loop_index63_load_reg_157 <= loop_index63_fu_60;
        mem_addr_read_reg_162 <= m_axi_mem_RDATA;
        sext_ln182_cast_reg_147 <= sext_ln182_cast_fu_98_p1;
    end
end

always @ (*) begin
    if (((exitcond84_fu_126_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_condition_exit_pp0_iter1_stage0 = 1'b1;
    end else begin
        ap_condition_exit_pp0_iter1_stage0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter2_reg == 1'b1))) begin
        ap_done_int = 1'b1;
    end else begin
        ap_done_int = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_idle_pp0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_start_int == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_ready_int = 1'b1;
    end else begin
        ap_ready_int = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        m_axi_mem_RREADY = 1'b1;
    end else begin
        m_axi_mem_RREADY = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        mem_blk_n_R = m_axi_mem_RVALID;
    end else begin
        mem_blk_n_R = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        node_y_coords_ce1 = 1'b1;
    end else begin
        node_y_coords_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        node_y_coords_we1 = 1'b1;
    end else begin
        node_y_coords_we1 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_pp0_stage0 : begin
            ap_NS_fsm = ap_ST_fsm_pp0_stage0;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_pp0_stage0_11001 = ((m_axi_mem_RVALID == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b1));
end

always @ (*) begin
    ap_block_pp0_stage0_subdone = ((m_axi_mem_RVALID == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b1));
end

assign ap_block_state1_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state2_pp0_stage0_iter1 = (m_axi_mem_RVALID == 1'b0);
end

assign ap_block_state3_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_enable_reg_pp0_iter0 = ap_start_int;

assign ap_loop_exit_ready = ap_condition_exit_pp0_iter1_stage0;

assign empty_fu_114_p2 = (loop_index63_fu_60 + 61'd1);

assign exitcond84_fu_126_p2 = ((empty_fu_114_p2 == sext_ln182_cast_reg_147) ? 1'b1 : 1'b0);

assign loop_index63_cast_fu_136_p1 = loop_index63_load_reg_157;

assign m_axi_mem_ARADDR = 64'd0;

assign m_axi_mem_ARBURST = 2'd0;

assign m_axi_mem_ARCACHE = 4'd0;

assign m_axi_mem_ARID = 1'd0;

assign m_axi_mem_ARLEN = 32'd0;

assign m_axi_mem_ARLOCK = 2'd0;

assign m_axi_mem_ARPROT = 3'd0;

assign m_axi_mem_ARQOS = 4'd0;

assign m_axi_mem_ARREGION = 4'd0;

assign m_axi_mem_ARSIZE = 3'd0;

assign m_axi_mem_ARUSER = 1'd0;

assign m_axi_mem_ARVALID = 1'b0;

assign m_axi_mem_AWADDR = 64'd0;

assign m_axi_mem_AWBURST = 2'd0;

assign m_axi_mem_AWCACHE = 4'd0;

assign m_axi_mem_AWID = 1'd0;

assign m_axi_mem_AWLEN = 32'd0;

assign m_axi_mem_AWLOCK = 2'd0;

assign m_axi_mem_AWPROT = 3'd0;

assign m_axi_mem_AWQOS = 4'd0;

assign m_axi_mem_AWREGION = 4'd0;

assign m_axi_mem_AWSIZE = 3'd0;

assign m_axi_mem_AWUSER = 1'd0;

assign m_axi_mem_AWVALID = 1'b0;

assign m_axi_mem_BREADY = 1'b0;

assign m_axi_mem_WDATA = 64'd0;

assign m_axi_mem_WID = 1'd0;

assign m_axi_mem_WLAST = 1'b0;

assign m_axi_mem_WSTRB = 8'd0;

assign m_axi_mem_WUSER = 1'd0;

assign m_axi_mem_WVALID = 1'b0;

assign node_y_coords_address1 = loop_index63_cast_fu_136_p1;

assign node_y_coords_d1 = mem_addr_read_reg_162;

assign sext_ln182_cast_fu_98_p1 = $signed(sext_ln182);

endmodule //kmeans_top_kmeans_top_Pipeline_2


// Content from kmeans_top_cfg_s_axi.v
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2022.2 (64-bit)
// Tool Version Limit: 2019.12
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1ns/1ps
module kmeans_top_cfg_s_axi
#(parameter
    C_S_AXI_ADDR_WIDTH = 8,
    C_S_AXI_DATA_WIDTH = 32
)(
    input  wire                          ACLK,
    input  wire                          ARESET,
    input  wire                          ACLK_EN,
    input  wire [C_S_AXI_ADDR_WIDTH-1:0] AWADDR,
    input  wire                          AWVALID,
    output wire                          AWREADY,
    input  wire [C_S_AXI_DATA_WIDTH-1:0] WDATA,
    input  wire [C_S_AXI_DATA_WIDTH/8-1:0] WSTRB,
    input  wire                          WVALID,
    output wire                          WREADY,
    output wire [1:0]                    BRESP,
    output wire                          BVALID,
    input  wire                          BREADY,
    input  wire [C_S_AXI_ADDR_WIDTH-1:0] ARADDR,
    input  wire                          ARVALID,
    output wire                          ARREADY,
    output wire [C_S_AXI_DATA_WIDTH-1:0] RDATA,
    output wire [1:0]                    RRESP,
    output wire                          RVALID,
    input  wire                          RREADY,
    output wire                          interrupt,
    output wire [31:0]                   n,
    output wire [31:0]                   k,
    output wire [31:0]                   control,
    output wire [63:0]                   buf_ptr_node_x_coords,
    output wire [63:0]                   buf_ptr_node_y_coords,
    output wire [63:0]                   buf_ptr_node_cluster_assignments,
    output wire [63:0]                   buf_ptr_centroid_x_coords,
    output wire [63:0]                   buf_ptr_centroid_y_coords,
    output wire [63:0]                   buf_ptr_intermediate_cluster_assignments,
    output wire [63:0]                   buf_ptr_intermediate_centroid_x_coords,
    output wire [63:0]                   buf_ptr_intermediate_centroid_y_coords,
    output wire [63:0]                   max_iterations,
    output wire [63:0]                   sub_iterations,
    output wire                          ap_start,
    input  wire                          ap_done,
    input  wire                          ap_ready,
    input  wire                          ap_idle
);
//------------------------Address Info-------------------
// 0x00 : Control signals
//        bit 0  - ap_start (Read/Write/COH)
//        bit 1  - ap_done (Read/COR)
//        bit 2  - ap_idle (Read)
//        bit 3  - ap_ready (Read/COR)
//        bit 7  - auto_restart (Read/Write)
//        bit 9  - interrupt (Read)
//        others - reserved
// 0x04 : Global Interrupt Enable Register
//        bit 0  - Global Interrupt Enable (Read/Write)
//        others - reserved
// 0x08 : IP Interrupt Enable Register (Read/Write)
//        bit 0 - enable ap_done interrupt (Read/Write)
//        bit 1 - enable ap_ready interrupt (Read/Write)
//        others - reserved
// 0x0c : IP Interrupt Status Register (Read/TOW)
//        bit 0 - ap_done (Read/TOW)
//        bit 1 - ap_ready (Read/TOW)
//        others - reserved
// 0x10 : Data signal of n
//        bit 31~0 - n[31:0] (Read/Write)
// 0x14 : reserved
// 0x18 : Data signal of k
//        bit 31~0 - k[31:0] (Read/Write)
// 0x1c : reserved
// 0x20 : Data signal of control
//        bit 31~0 - control[31:0] (Read/Write)
// 0x24 : reserved
// 0x28 : Data signal of buf_ptr_node_x_coords
//        bit 31~0 - buf_ptr_node_x_coords[31:0] (Read/Write)
// 0x2c : Data signal of buf_ptr_node_x_coords
//        bit 31~0 - buf_ptr_node_x_coords[63:32] (Read/Write)
// 0x30 : reserved
// 0x34 : Data signal of buf_ptr_node_y_coords
//        bit 31~0 - buf_ptr_node_y_coords[31:0] (Read/Write)
// 0x38 : Data signal of buf_ptr_node_y_coords
//        bit 31~0 - buf_ptr_node_y_coords[63:32] (Read/Write)
// 0x3c : reserved
// 0x40 : Data signal of buf_ptr_node_cluster_assignments
//        bit 31~0 - buf_ptr_node_cluster_assignments[31:0] (Read/Write)
// 0x44 : Data signal of buf_ptr_node_cluster_assignments
//        bit 31~0 - buf_ptr_node_cluster_assignments[63:32] (Read/Write)
// 0x48 : reserved
// 0x4c : Data signal of buf_ptr_centroid_x_coords
//        bit 31~0 - buf_ptr_centroid_x_coords[31:0] (Read/Write)
// 0x50 : Data signal of buf_ptr_centroid_x_coords
//        bit 31~0 - buf_ptr_centroid_x_coords[63:32] (Read/Write)
// 0x54 : reserved
// 0x58 : Data signal of buf_ptr_centroid_y_coords
//        bit 31~0 - buf_ptr_centroid_y_coords[31:0] (Read/Write)
// 0x5c : Data signal of buf_ptr_centroid_y_coords
//        bit 31~0 - buf_ptr_centroid_y_coords[63:32] (Read/Write)
// 0x60 : reserved
// 0x64 : Data signal of buf_ptr_intermediate_cluster_assignments
//        bit 31~0 - buf_ptr_intermediate_cluster_assignments[31:0] (Read/Write)
// 0x68 : Data signal of buf_ptr_intermediate_cluster_assignments
//        bit 31~0 - buf_ptr_intermediate_cluster_assignments[63:32] (Read/Write)
// 0x6c : reserved
// 0x70 : Data signal of buf_ptr_intermediate_centroid_x_coords
//        bit 31~0 - buf_ptr_intermediate_centroid_x_coords[31:0] (Read/Write)
// 0x74 : Data signal of buf_ptr_intermediate_centroid_x_coords
//        bit 31~0 - buf_ptr_intermediate_centroid_x_coords[63:32] (Read/Write)
// 0x78 : reserved
// 0x7c : Data signal of buf_ptr_intermediate_centroid_y_coords
//        bit 31~0 - buf_ptr_intermediate_centroid_y_coords[31:0] (Read/Write)
// 0x80 : Data signal of buf_ptr_intermediate_centroid_y_coords
//        bit 31~0 - buf_ptr_intermediate_centroid_y_coords[63:32] (Read/Write)
// 0x84 : reserved
// 0x88 : Data signal of max_iterations
//        bit 31~0 - max_iterations[31:0] (Read/Write)
// 0x8c : Data signal of max_iterations
//        bit 31~0 - max_iterations[63:32] (Read/Write)
// 0x90 : reserved
// 0x94 : Data signal of sub_iterations
//        bit 31~0 - sub_iterations[31:0] (Read/Write)
// 0x98 : Data signal of sub_iterations
//        bit 31~0 - sub_iterations[63:32] (Read/Write)
// 0x9c : reserved
// (SC = Self Clear, COR = Clear on Read, TOW = Toggle on Write, COH = Clear on Handshake)

//------------------------Parameter----------------------
localparam
    ADDR_AP_CTRL                                         = 8'h00,
    ADDR_GIE                                             = 8'h04,
    ADDR_IER                                             = 8'h08,
    ADDR_ISR                                             = 8'h0c,
    ADDR_N_DATA_0                                        = 8'h10,
    ADDR_N_CTRL                                          = 8'h14,
    ADDR_K_DATA_0                                        = 8'h18,
    ADDR_K_CTRL                                          = 8'h1c,
    ADDR_CONTROL_DATA_0                                  = 8'h20,
    ADDR_CONTROL_CTRL                                    = 8'h24,
    ADDR_BUF_PTR_NODE_X_COORDS_DATA_0                    = 8'h28,
    ADDR_BUF_PTR_NODE_X_COORDS_DATA_1                    = 8'h2c,
    ADDR_BUF_PTR_NODE_X_COORDS_CTRL                      = 8'h30,
    ADDR_BUF_PTR_NODE_Y_COORDS_DATA_0                    = 8'h34,
    ADDR_BUF_PTR_NODE_Y_COORDS_DATA_1                    = 8'h38,
    ADDR_BUF_PTR_NODE_Y_COORDS_CTRL                      = 8'h3c,
    ADDR_BUF_PTR_NODE_CLUSTER_ASSIGNMENTS_DATA_0         = 8'h40,
    ADDR_BUF_PTR_NODE_CLUSTER_ASSIGNMENTS_DATA_1         = 8'h44,
    ADDR_BUF_PTR_NODE_CLUSTER_ASSIGNMENTS_CTRL           = 8'h48,
    ADDR_BUF_PTR_CENTROID_X_COORDS_DATA_0                = 8'h4c,
    ADDR_BUF_PTR_CENTROID_X_COORDS_DATA_1                = 8'h50,
    ADDR_BUF_PTR_CENTROID_X_COORDS_CTRL                  = 8'h54,
    ADDR_BUF_PTR_CENTROID_Y_COORDS_DATA_0                = 8'h58,
    ADDR_BUF_PTR_CENTROID_Y_COORDS_DATA_1                = 8'h5c,
    ADDR_BUF_PTR_CENTROID_Y_COORDS_CTRL                  = 8'h60,
    ADDR_BUF_PTR_INTERMEDIATE_CLUSTER_ASSIGNMENTS_DATA_0 = 8'h64,
    ADDR_BUF_PTR_INTERMEDIATE_CLUSTER_ASSIGNMENTS_DATA_1 = 8'h68,
    ADDR_BUF_PTR_INTERMEDIATE_CLUSTER_ASSIGNMENTS_CTRL   = 8'h6c,
    ADDR_BUF_PTR_INTERMEDIATE_CENTROID_X_COORDS_DATA_0   = 8'h70,
    ADDR_BUF_PTR_INTERMEDIATE_CENTROID_X_COORDS_DATA_1   = 8'h74,
    ADDR_BUF_PTR_INTERMEDIATE_CENTROID_X_COORDS_CTRL     = 8'h78,
    ADDR_BUF_PTR_INTERMEDIATE_CENTROID_Y_COORDS_DATA_0   = 8'h7c,
    ADDR_BUF_PTR_INTERMEDIATE_CENTROID_Y_COORDS_DATA_1   = 8'h80,
    ADDR_BUF_PTR_INTERMEDIATE_CENTROID_Y_COORDS_CTRL     = 8'h84,
    ADDR_MAX_ITERATIONS_DATA_0                           = 8'h88,
    ADDR_MAX_ITERATIONS_DATA_1                           = 8'h8c,
    ADDR_MAX_ITERATIONS_CTRL                             = 8'h90,
    ADDR_SUB_ITERATIONS_DATA_0                           = 8'h94,
    ADDR_SUB_ITERATIONS_DATA_1                           = 8'h98,
    ADDR_SUB_ITERATIONS_CTRL                             = 8'h9c,
    WRIDLE                                               = 2'd0,
    WRDATA                                               = 2'd1,
    WRRESP                                               = 2'd2,
    WRRESET                                              = 2'd3,
    RDIDLE                                               = 2'd0,
    RDDATA                                               = 2'd1,
    RDRESET                                              = 2'd2,
    ADDR_BITS                = 8;

//------------------------Local signal-------------------
    reg  [1:0]                    wstate = WRRESET;
    reg  [1:0]                    wnext;
    reg  [ADDR_BITS-1:0]          waddr;
    wire [C_S_AXI_DATA_WIDTH-1:0] wmask;
    wire                          aw_hs;
    wire                          w_hs;
    reg  [1:0]                    rstate = RDRESET;
    reg  [1:0]                    rnext;
    reg  [C_S_AXI_DATA_WIDTH-1:0] rdata;
    wire                          ar_hs;
    wire [ADDR_BITS-1:0]          raddr;
    // internal registers
    reg                           int_ap_idle;
    reg                           int_ap_ready = 1'b0;
    wire                          task_ap_ready;
    reg                           int_ap_done = 1'b0;
    wire                          task_ap_done;
    reg                           int_task_ap_done = 1'b0;
    reg                           int_ap_start = 1'b0;
    reg                           int_interrupt = 1'b0;
    reg                           int_auto_restart = 1'b0;
    reg                           auto_restart_status = 1'b0;
    wire                          auto_restart_done;
    reg                           int_gie = 1'b0;
    reg  [1:0]                    int_ier = 2'b0;
    reg  [1:0]                    int_isr = 2'b0;
    reg  [31:0]                   int_n = 'b0;
    reg  [31:0]                   int_k = 'b0;
    reg  [31:0]                   int_control = 'b0;
    reg  [63:0]                   int_buf_ptr_node_x_coords = 'b0;
    reg  [63:0]                   int_buf_ptr_node_y_coords = 'b0;
    reg  [63:0]                   int_buf_ptr_node_cluster_assignments = 'b0;
    reg  [63:0]                   int_buf_ptr_centroid_x_coords = 'b0;
    reg  [63:0]                   int_buf_ptr_centroid_y_coords = 'b0;
    reg  [63:0]                   int_buf_ptr_intermediate_cluster_assignments = 'b0;
    reg  [63:0]                   int_buf_ptr_intermediate_centroid_x_coords = 'b0;
    reg  [63:0]                   int_buf_ptr_intermediate_centroid_y_coords = 'b0;
    reg  [63:0]                   int_max_iterations = 'b0;
    reg  [63:0]                   int_sub_iterations = 'b0;

//------------------------Instantiation------------------


//------------------------AXI write fsm------------------
assign AWREADY = (wstate == WRIDLE);
assign WREADY  = (wstate == WRDATA);
assign BRESP   = 2'b00;  // OKAY
assign BVALID  = (wstate == WRRESP);
assign wmask   = { {8{WSTRB[3]}}, {8{WSTRB[2]}}, {8{WSTRB[1]}}, {8{WSTRB[0]}} };
assign aw_hs   = AWVALID & AWREADY;
assign w_hs    = WVALID & WREADY;

// wstate
always @(posedge ACLK) begin
    if (ARESET)
        wstate <= WRRESET;
    else if (ACLK_EN)
        wstate <= wnext;
end

// wnext
always @(*) begin
    case (wstate)
        WRIDLE:
            if (AWVALID)
                wnext = WRDATA;
            else
                wnext = WRIDLE;
        WRDATA:
            if (WVALID)
                wnext = WRRESP;
            else
                wnext = WRDATA;
        WRRESP:
            if (BREADY)
                wnext = WRIDLE;
            else
                wnext = WRRESP;
        default:
            wnext = WRIDLE;
    endcase
end

// waddr
always @(posedge ACLK) begin
    if (ACLK_EN) begin
        if (aw_hs)
            waddr <= AWADDR[ADDR_BITS-1:0];
    end
end

//------------------------AXI read fsm-------------------
assign ARREADY = (rstate == RDIDLE);
assign RDATA   = rdata;
assign RRESP   = 2'b00;  // OKAY
assign RVALID  = (rstate == RDDATA);
assign ar_hs   = ARVALID & ARREADY;
assign raddr   = ARADDR[ADDR_BITS-1:0];

// rstate
always @(posedge ACLK) begin
    if (ARESET)
        rstate <= RDRESET;
    else if (ACLK_EN)
        rstate <= rnext;
end

// rnext
always @(*) begin
    case (rstate)
        RDIDLE:
            if (ARVALID)
                rnext = RDDATA;
            else
                rnext = RDIDLE;
        RDDATA:
            if (RREADY & RVALID)
                rnext = RDIDLE;
            else
                rnext = RDDATA;
        default:
            rnext = RDIDLE;
    endcase
end

// rdata
always @(posedge ACLK) begin
    if (ACLK_EN) begin
        if (ar_hs) begin
            rdata <= 'b0;
            case (raddr)
                ADDR_AP_CTRL: begin
                    rdata[0] <= int_ap_start;
                    rdata[1] <= int_task_ap_done;
                    rdata[2] <= int_ap_idle;
                    rdata[3] <= int_ap_ready;
                    rdata[7] <= int_auto_restart;
                    rdata[9] <= int_interrupt;
                end
                ADDR_GIE: begin
                    rdata <= int_gie;
                end
                ADDR_IER: begin
                    rdata <= int_ier;
                end
                ADDR_ISR: begin
                    rdata <= int_isr;
                end
                ADDR_N_DATA_0: begin
                    rdata <= int_n[31:0];
                end
                ADDR_K_DATA_0: begin
                    rdata <= int_k[31:0];
                end
                ADDR_CONTROL_DATA_0: begin
                    rdata <= int_control[31:0];
                end
                ADDR_BUF_PTR_NODE_X_COORDS_DATA_0: begin
                    rdata <= int_buf_ptr_node_x_coords[31:0];
                end
                ADDR_BUF_PTR_NODE_X_COORDS_DATA_1: begin
                    rdata <= int_buf_ptr_node_x_coords[63:32];
                end
                ADDR_BUF_PTR_NODE_Y_COORDS_DATA_0: begin
                    rdata <= int_buf_ptr_node_y_coords[31:0];
                end
                ADDR_BUF_PTR_NODE_Y_COORDS_DATA_1: begin
                    rdata <= int_buf_ptr_node_y_coords[63:32];
                end
                ADDR_BUF_PTR_NODE_CLUSTER_ASSIGNMENTS_DATA_0: begin
                    rdata <= int_buf_ptr_node_cluster_assignments[31:0];
                end
                ADDR_BUF_PTR_NODE_CLUSTER_ASSIGNMENTS_DATA_1: begin
                    rdata <= int_buf_ptr_node_cluster_assignments[63:32];
                end
                ADDR_BUF_PTR_CENTROID_X_COORDS_DATA_0: begin
                    rdata <= int_buf_ptr_centroid_x_coords[31:0];
                end
                ADDR_BUF_PTR_CENTROID_X_COORDS_DATA_1: begin
                    rdata <= int_buf_ptr_centroid_x_coords[63:32];
                end
                ADDR_BUF_PTR_CENTROID_Y_COORDS_DATA_0: begin
                    rdata <= int_buf_ptr_centroid_y_coords[31:0];
                end
                ADDR_BUF_PTR_CENTROID_Y_COORDS_DATA_1: begin
                    rdata <= int_buf_ptr_centroid_y_coords[63:32];
                end
                ADDR_BUF_PTR_INTERMEDIATE_CLUSTER_ASSIGNMENTS_DATA_0: begin
                    rdata <= int_buf_ptr_intermediate_cluster_assignments[31:0];
                end
                ADDR_BUF_PTR_INTERMEDIATE_CLUSTER_ASSIGNMENTS_DATA_1: begin
                    rdata <= int_buf_ptr_intermediate_cluster_assignments[63:32];
                end
                ADDR_BUF_PTR_INTERMEDIATE_CENTROID_X_COORDS_DATA_0: begin
                    rdata <= int_buf_ptr_intermediate_centroid_x_coords[31:0];
                end
                ADDR_BUF_PTR_INTERMEDIATE_CENTROID_X_COORDS_DATA_1: begin
                    rdata <= int_buf_ptr_intermediate_centroid_x_coords[63:32];
                end
                ADDR_BUF_PTR_INTERMEDIATE_CENTROID_Y_COORDS_DATA_0: begin
                    rdata <= int_buf_ptr_intermediate_centroid_y_coords[31:0];
                end
                ADDR_BUF_PTR_INTERMEDIATE_CENTROID_Y_COORDS_DATA_1: begin
                    rdata <= int_buf_ptr_intermediate_centroid_y_coords[63:32];
                end
                ADDR_MAX_ITERATIONS_DATA_0: begin
                    rdata <= int_max_iterations[31:0];
                end
                ADDR_MAX_ITERATIONS_DATA_1: begin
                    rdata <= int_max_iterations[63:32];
                end
                ADDR_SUB_ITERATIONS_DATA_0: begin
                    rdata <= int_sub_iterations[31:0];
                end
                ADDR_SUB_ITERATIONS_DATA_1: begin
                    rdata <= int_sub_iterations[63:32];
                end
            endcase
        end
    end
end


//------------------------Register logic-----------------
assign interrupt                                = int_interrupt;
assign ap_start                                 = int_ap_start;
assign task_ap_done                             = (ap_done && !auto_restart_status) || auto_restart_done;
assign task_ap_ready                            = ap_ready && !int_auto_restart;
assign auto_restart_done                        = auto_restart_status && (ap_idle && !int_ap_idle);
assign n                                        = int_n;
assign k                                        = int_k;
assign control                                  = int_control;
assign buf_ptr_node_x_coords                    = int_buf_ptr_node_x_coords;
assign buf_ptr_node_y_coords                    = int_buf_ptr_node_y_coords;
assign buf_ptr_node_cluster_assignments         = int_buf_ptr_node_cluster_assignments;
assign buf_ptr_centroid_x_coords                = int_buf_ptr_centroid_x_coords;
assign buf_ptr_centroid_y_coords                = int_buf_ptr_centroid_y_coords;
assign buf_ptr_intermediate_cluster_assignments = int_buf_ptr_intermediate_cluster_assignments;
assign buf_ptr_intermediate_centroid_x_coords   = int_buf_ptr_intermediate_centroid_x_coords;
assign buf_ptr_intermediate_centroid_y_coords   = int_buf_ptr_intermediate_centroid_y_coords;
assign max_iterations                           = int_max_iterations;
assign sub_iterations                           = int_sub_iterations;
// int_interrupt
always @(posedge ACLK) begin
    if (ARESET)
        int_interrupt <= 1'b0;
    else if (ACLK_EN) begin
        if (int_gie && (|int_isr))
            int_interrupt <= 1'b1;
        else
            int_interrupt <= 1'b0;
    end
end

// int_ap_start
always @(posedge ACLK) begin
    if (ARESET)
        int_ap_start <= 1'b0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_AP_CTRL && WSTRB[0] && WDATA[0])
            int_ap_start <= 1'b1;
        else if (ap_ready)
            int_ap_start <= int_auto_restart; // clear on handshake/auto restart
    end
end

// int_ap_done
always @(posedge ACLK) begin
    if (ARESET)
        int_ap_done <= 1'b0;
    else if (ACLK_EN) begin
            int_ap_done <= ap_done;
    end
end

// int_task_ap_done
always @(posedge ACLK) begin
    if (ARESET)
        int_task_ap_done <= 1'b0;
    else if (ACLK_EN) begin
        if (task_ap_done)
            int_task_ap_done <= 1'b1;
        else if (ar_hs && raddr == ADDR_AP_CTRL)
            int_task_ap_done <= 1'b0; // clear on read
    end
end

// int_ap_idle
always @(posedge ACLK) begin
    if (ARESET)
        int_ap_idle <= 1'b0;
    else if (ACLK_EN) begin
            int_ap_idle <= ap_idle;
    end
end

// int_ap_ready
always @(posedge ACLK) begin
    if (ARESET)
        int_ap_ready <= 1'b0;
    else if (ACLK_EN) begin
        if (task_ap_ready)
            int_ap_ready <= 1'b1;
        else if (ar_hs && raddr == ADDR_AP_CTRL)
            int_ap_ready <= 1'b0;
    end
end

// int_auto_restart
always @(posedge ACLK) begin
    if (ARESET)
        int_auto_restart <= 1'b0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_AP_CTRL && WSTRB[0])
            int_auto_restart <=  WDATA[7];
    end
end

// auto_restart_status
always @(posedge ACLK) begin
    if (ARESET)
        auto_restart_status <= 1'b0;
    else if (ACLK_EN) begin
        if (int_auto_restart)
            auto_restart_status <= 1'b1;
        else if (ap_idle)
            auto_restart_status <= 1'b0;
    end
end

// int_gie
always @(posedge ACLK) begin
    if (ARESET)
        int_gie <= 1'b0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_GIE && WSTRB[0])
            int_gie <= WDATA[0];
    end
end

// int_ier
always @(posedge ACLK) begin
    if (ARESET)
        int_ier <= 1'b0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_IER && WSTRB[0])
            int_ier <= WDATA[1:0];
    end
end

// int_isr[0]
always @(posedge ACLK) begin
    if (ARESET)
        int_isr[0] <= 1'b0;
    else if (ACLK_EN) begin
        if (int_ier[0] & ap_done)
            int_isr[0] <= 1'b1;
        else if (w_hs && waddr == ADDR_ISR && WSTRB[0])
            int_isr[0] <= int_isr[0] ^ WDATA[0]; // toggle on write
    end
end

// int_isr[1]
always @(posedge ACLK) begin
    if (ARESET)
        int_isr[1] <= 1'b0;
    else if (ACLK_EN) begin
        if (int_ier[1] & ap_ready)
            int_isr[1] <= 1'b1;
        else if (w_hs && waddr == ADDR_ISR && WSTRB[0])
            int_isr[1] <= int_isr[1] ^ WDATA[1]; // toggle on write
    end
end

// int_n[31:0]
always @(posedge ACLK) begin
    if (ARESET)
        int_n[31:0] <= 0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_N_DATA_0)
            int_n[31:0] <= (WDATA[31:0] & wmask) | (int_n[31:0] & ~wmask);
    end
end

// int_k[31:0]
always @(posedge ACLK) begin
    if (ARESET)
        int_k[31:0] <= 0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_K_DATA_0)
            int_k[31:0] <= (WDATA[31:0] & wmask) | (int_k[31:0] & ~wmask);
    end
end

// int_control[31:0]
always @(posedge ACLK) begin
    if (ARESET)
        int_control[31:0] <= 0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_CONTROL_DATA_0)
            int_control[31:0] <= (WDATA[31:0] & wmask) | (int_control[31:0] & ~wmask);
    end
end

// int_buf_ptr_node_x_coords[31:0]
always @(posedge ACLK) begin
    if (ARESET)
        int_buf_ptr_node_x_coords[31:0] <= 0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_BUF_PTR_NODE_X_COORDS_DATA_0)
            int_buf_ptr_node_x_coords[31:0] <= (WDATA[31:0] & wmask) | (int_buf_ptr_node_x_coords[31:0] & ~wmask);
    end
end

// int_buf_ptr_node_x_coords[63:32]
always @(posedge ACLK) begin
    if (ARESET)
        int_buf_ptr_node_x_coords[63:32] <= 0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_BUF_PTR_NODE_X_COORDS_DATA_1)
            int_buf_ptr_node_x_coords[63:32] <= (WDATA[31:0] & wmask) | (int_buf_ptr_node_x_coords[63:32] & ~wmask);
    end
end

// int_buf_ptr_node_y_coords[31:0]
always @(posedge ACLK) begin
    if (ARESET)
        int_buf_ptr_node_y_coords[31:0] <= 0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_BUF_PTR_NODE_Y_COORDS_DATA_0)
            int_buf_ptr_node_y_coords[31:0] <= (WDATA[31:0] & wmask) | (int_buf_ptr_node_y_coords[31:0] & ~wmask);
    end
end

// int_buf_ptr_node_y_coords[63:32]
always @(posedge ACLK) begin
    if (ARESET)
        int_buf_ptr_node_y_coords[63:32] <= 0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_BUF_PTR_NODE_Y_COORDS_DATA_1)
            int_buf_ptr_node_y_coords[63:32] <= (WDATA[31:0] & wmask) | (int_buf_ptr_node_y_coords[63:32] & ~wmask);
    end
end

// int_buf_ptr_node_cluster_assignments[31:0]
always @(posedge ACLK) begin
    if (ARESET)
        int_buf_ptr_node_cluster_assignments[31:0] <= 0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_BUF_PTR_NODE_CLUSTER_ASSIGNMENTS_DATA_0)
            int_buf_ptr_node_cluster_assignments[31:0] <= (WDATA[31:0] & wmask) | (int_buf_ptr_node_cluster_assignments[31:0] & ~wmask);
    end
end

// int_buf_ptr_node_cluster_assignments[63:32]
always @(posedge ACLK) begin
    if (ARESET)
        int_buf_ptr_node_cluster_assignments[63:32] <= 0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_BUF_PTR_NODE_CLUSTER_ASSIGNMENTS_DATA_1)
            int_buf_ptr_node_cluster_assignments[63:32] <= (WDATA[31:0] & wmask) | (int_buf_ptr_node_cluster_assignments[63:32] & ~wmask);
    end
end

// int_buf_ptr_centroid_x_coords[31:0]
always @(posedge ACLK) begin
    if (ARESET)
        int_buf_ptr_centroid_x_coords[31:0] <= 0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_BUF_PTR_CENTROID_X_COORDS_DATA_0)
            int_buf_ptr_centroid_x_coords[31:0] <= (WDATA[31:0] & wmask) | (int_buf_ptr_centroid_x_coords[31:0] & ~wmask);
    end
end

// int_buf_ptr_centroid_x_coords[63:32]
always @(posedge ACLK) begin
    if (ARESET)
        int_buf_ptr_centroid_x_coords[63:32] <= 0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_BUF_PTR_CENTROID_X_COORDS_DATA_1)
            int_buf_ptr_centroid_x_coords[63:32] <= (WDATA[31:0] & wmask) | (int_buf_ptr_centroid_x_coords[63:32] & ~wmask);
    end
end

// int_buf_ptr_centroid_y_coords[31:0]
always @(posedge ACLK) begin
    if (ARESET)
        int_buf_ptr_centroid_y_coords[31:0] <= 0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_BUF_PTR_CENTROID_Y_COORDS_DATA_0)
            int_buf_ptr_centroid_y_coords[31:0] <= (WDATA[31:0] & wmask) | (int_buf_ptr_centroid_y_coords[31:0] & ~wmask);
    end
end

// int_buf_ptr_centroid_y_coords[63:32]
always @(posedge ACLK) begin
    if (ARESET)
        int_buf_ptr_centroid_y_coords[63:32] <= 0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_BUF_PTR_CENTROID_Y_COORDS_DATA_1)
            int_buf_ptr_centroid_y_coords[63:32] <= (WDATA[31:0] & wmask) | (int_buf_ptr_centroid_y_coords[63:32] & ~wmask);
    end
end

// int_buf_ptr_intermediate_cluster_assignments[31:0]
always @(posedge ACLK) begin
    if (ARESET)
        int_buf_ptr_intermediate_cluster_assignments[31:0] <= 0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_BUF_PTR_INTERMEDIATE_CLUSTER_ASSIGNMENTS_DATA_0)
            int_buf_ptr_intermediate_cluster_assignments[31:0] <= (WDATA[31:0] & wmask) | (int_buf_ptr_intermediate_cluster_assignments[31:0] & ~wmask);
    end
end

// int_buf_ptr_intermediate_cluster_assignments[63:32]
always @(posedge ACLK) begin
    if (ARESET)
        int_buf_ptr_intermediate_cluster_assignments[63:32] <= 0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_BUF_PTR_INTERMEDIATE_CLUSTER_ASSIGNMENTS_DATA_1)
            int_buf_ptr_intermediate_cluster_assignments[63:32] <= (WDATA[31:0] & wmask) | (int_buf_ptr_intermediate_cluster_assignments[63:32] & ~wmask);
    end
end

// int_buf_ptr_intermediate_centroid_x_coords[31:0]
always @(posedge ACLK) begin
    if (ARESET)
        int_buf_ptr_intermediate_centroid_x_coords[31:0] <= 0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_BUF_PTR_INTERMEDIATE_CENTROID_X_COORDS_DATA_0)
            int_buf_ptr_intermediate_centroid_x_coords[31:0] <= (WDATA[31:0] & wmask) | (int_buf_ptr_intermediate_centroid_x_coords[31:0] & ~wmask);
    end
end

// int_buf_ptr_intermediate_centroid_x_coords[63:32]
always @(posedge ACLK) begin
    if (ARESET)
        int_buf_ptr_intermediate_centroid_x_coords[63:32] <= 0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_BUF_PTR_INTERMEDIATE_CENTROID_X_COORDS_DATA_1)
            int_buf_ptr_intermediate_centroid_x_coords[63:32] <= (WDATA[31:0] & wmask) | (int_buf_ptr_intermediate_centroid_x_coords[63:32] & ~wmask);
    end
end

// int_buf_ptr_intermediate_centroid_y_coords[31:0]
always @(posedge ACLK) begin
    if (ARESET)
        int_buf_ptr_intermediate_centroid_y_coords[31:0] <= 0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_BUF_PTR_INTERMEDIATE_CENTROID_Y_COORDS_DATA_0)
            int_buf_ptr_intermediate_centroid_y_coords[31:0] <= (WDATA[31:0] & wmask) | (int_buf_ptr_intermediate_centroid_y_coords[31:0] & ~wmask);
    end
end

// int_buf_ptr_intermediate_centroid_y_coords[63:32]
always @(posedge ACLK) begin
    if (ARESET)
        int_buf_ptr_intermediate_centroid_y_coords[63:32] <= 0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_BUF_PTR_INTERMEDIATE_CENTROID_Y_COORDS_DATA_1)
            int_buf_ptr_intermediate_centroid_y_coords[63:32] <= (WDATA[31:0] & wmask) | (int_buf_ptr_intermediate_centroid_y_coords[63:32] & ~wmask);
    end
end

// int_max_iterations[31:0]
always @(posedge ACLK) begin
    if (ARESET)
        int_max_iterations[31:0] <= 0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_MAX_ITERATIONS_DATA_0)
            int_max_iterations[31:0] <= (WDATA[31:0] & wmask) | (int_max_iterations[31:0] & ~wmask);
    end
end

// int_max_iterations[63:32]
always @(posedge ACLK) begin
    if (ARESET)
        int_max_iterations[63:32] <= 0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_MAX_ITERATIONS_DATA_1)
            int_max_iterations[63:32] <= (WDATA[31:0] & wmask) | (int_max_iterations[63:32] & ~wmask);
    end
end

// int_sub_iterations[31:0]
always @(posedge ACLK) begin
    if (ARESET)
        int_sub_iterations[31:0] <= 0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_SUB_ITERATIONS_DATA_0)
            int_sub_iterations[31:0] <= (WDATA[31:0] & wmask) | (int_sub_iterations[31:0] & ~wmask);
    end
end

// int_sub_iterations[63:32]
always @(posedge ACLK) begin
    if (ARESET)
        int_sub_iterations[63:32] <= 0;
    else if (ACLK_EN) begin
        if (w_hs && waddr == ADDR_SUB_ITERATIONS_DATA_1)
            int_sub_iterations[63:32] <= (WDATA[31:0] & wmask) | (int_sub_iterations[63:32] & ~wmask);
    end
end

//synthesis translate_off
always @(posedge ACLK) begin
    if (ACLK_EN) begin
        if (int_gie & ~int_isr[0] & int_ier[0] & ap_done)
            $display ("// Interrupt Monitor : interrupt for ap_done detected @ \"%0t\"", $time);
        if (int_gie & ~int_isr[1] & int_ier[1] & ap_ready)
            $display ("// Interrupt Monitor : interrupt for ap_ready detected @ \"%0t\"", $time);
    end
end
//synthesis translate_on

//------------------------Memory logic-------------------

endmodule


// Content from kmeans_top_node_cluster_assignments_RAM_2P_URAM_1R1W.v
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2022.2 (64-bit)
// Version: 2022.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module kmeans_top_node_cluster_assignments_RAM_2P_URAM_1R1W (
     
    address0, ce0,
    
    q0, 
      
    address1, ce1,
    d1, we1, 
    
     
    reset, clk);

parameter DataWidth = 64;
parameter AddressWidth = 13;
parameter AddressRange = 8192;
 
input[AddressWidth-1:0] address0;
input ce0;

output reg[DataWidth-1:0] q0; 
 
input[AddressWidth-1:0] address1;
input ce1;
input[DataWidth-1:0] d1;
input we1; 


input reset;
input clk;

(* ram_style = "hls_ultra" , cascade_height = 1 *)reg [DataWidth-1:0] ram[0:AddressRange-1];


 



always @(posedge clk) 
begin 
    if (ce0) begin
        q0 <= ram[address0];
    end
end 

 
  

always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[address1] <= d1; 
    end
end 



 
 

endmodule



// Content from kmeans_top_kmeans_Pipeline_VITIS_LOOP_116_6.v
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2022.2 (64-bit)
// Version: 2022.2
// Copyright (C) Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module kmeans_top_kmeans_Pipeline_VITIS_LOOP_116_6 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        k,
        centroid_y_coords_address0,
        centroid_y_coords_ce0,
        centroid_y_coords_q0,
        centroid_x_coords_prev_address0,
        centroid_x_coords_prev_ce0,
        centroid_x_coords_prev_q0,
        centroid_x_coords_address0,
        centroid_x_coords_ce0,
        centroid_x_coords_q0,
        ap_return
);

parameter    ap_ST_fsm_state1 = 3'd1;
parameter    ap_ST_fsm_state2 = 3'd2;
parameter    ap_ST_fsm_state3 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
input  [30:0] k;
output  [7:0] centroid_y_coords_address0;
output   centroid_y_coords_ce0;
input  [63:0] centroid_y_coords_q0;
output  [7:0] centroid_x_coords_prev_address0;
output   centroid_x_coords_prev_ce0;
input  [63:0] centroid_x_coords_prev_q0;
output  [7:0] centroid_x_coords_address0;
output   centroid_x_coords_ce0;
input  [63:0] centroid_x_coords_q0;
output  [1:0] ap_return;

reg ap_idle;
reg centroid_y_coords_ce0;
reg[7:0] centroid_x_coords_prev_address0;
reg centroid_x_coords_prev_ce0;
reg centroid_x_coords_ce0;
reg[1:0] ap_return;

(* fsm_encoding = "none" *) reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
wire    ap_CS_fsm_state3;
wire    ap_block_state3_pp0_stage2_iter0;
wire   [0:0] icmp_ln117_1_fu_133_p2;
reg   [0:0] icmp_ln117_reg_174;
reg   [0:0] icmp_ln116_reg_150;
reg    ap_condition_exit_pp0_iter0_stage2;
wire    ap_loop_exit_ready;
reg    ap_ready_int;
reg   [1:0] merge_reg_85;
wire   [0:0] icmp_ln116_fu_109_p2;
reg    ap_block_state1_pp0_stage0_iter0;
wire   [30:0] add_ln116_fu_115_p2;
reg   [30:0] add_ln116_reg_154;
wire   [63:0] i_3_cast7_fu_121_p1;
reg   [63:0] i_3_cast7_reg_159;
reg   [7:0] centroid_x_coords_prev_addr_reg_164;
wire   [0:0] icmp_ln117_fu_127_p2;
wire    ap_CS_fsm_state2;
wire    ap_block_state2_pp0_stage1_iter0;
reg   [1:0] ap_phi_mux_merge_phi_fu_90_p6;
reg   [30:0] i_fu_36;
wire    ap_loop_init;
reg   [30:0] ap_sig_allocacmp_i_1;
reg   [1:0] ap_return_preg;
reg    ap_done_reg;
wire    ap_continue_int;
reg    ap_done_int;
reg   [2:0] ap_NS_fsm;
reg    ap_ST_fsm_state1_blk;
wire    ap_ST_fsm_state2_blk;
wire    ap_ST_fsm_state3_blk;
wire    ap_start_int;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_CS_fsm = 3'd1;
#0 ap_return_preg = 2'd0;
#0 ap_done_reg = 1'b0;
end

kmeans_top_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(ap_start),
    .ap_ready(ap_ready),
    .ap_done(ap_done),
    .ap_start_int(ap_start_int),
    .ap_loop_init(ap_loop_init),
    .ap_ready_int(ap_ready_int),
    .ap_loop_exit_ready(ap_condition_exit_pp0_iter0_stage2),
    .ap_loop_exit_done(ap_done_int),
    .ap_continue_int(ap_continue_int),
    .ap_done_int(ap_done_int)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue_int == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((ap_loop_exit_ready == 1'b1) & (1'b1 == ap_CS_fsm_state3))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_return_preg <= 2'd0;
    end else begin
        if (((1'b1 == ap_CS_fsm_state3) & ((icmp_ln116_reg_150 == 1'd0) | ((icmp_ln117_reg_174 == 1'd0) | (icmp_ln117_1_fu_133_p2 == 1'd0))))) begin
            ap_return_preg <= ap_phi_mux_merge_phi_fu_90_p6;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start_int == 1'b1) & (ap_loop_init == 1'b1))) begin
        i_fu_36 <= 31'd0;
    end else if (((icmp_ln116_reg_150 == 1'd1) & (icmp_ln117_reg_174 == 1'd1) & (icmp_ln117_1_fu_133_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state3))) begin
        i_fu_36 <= add_ln116_reg_154;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln116_reg_150 == 1'd1) & (1'b1 == ap_CS_fsm_state2) & (icmp_ln117_fu_127_p2 == 1'd0))) begin
        merge_reg_85 <= 2'd2;
    end else if (((icmp_ln116_reg_150 == 1'd1) & (icmp_ln117_reg_174 == 1'd1) & (icmp_ln117_1_fu_133_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state3))) begin
        merge_reg_85 <= 2'd1;
    end else if (((icmp_ln116_fu_109_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state1) & (ap_start_int == 1'b1))) begin
        merge_reg_85 <= 2'd0;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start_int == 1'b1))) begin
        add_ln116_reg_154 <= add_ln116_fu_115_p2;
        icmp_ln116_reg_150 <= icmp_ln116_fu_109_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln116_fu_109_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1) & (ap_start_int == 1'b1))) begin
        centroid_x_coords_prev_addr_reg_164 <= i_3_cast7_fu_121_p1;
        i_3_cast7_reg_159[30 : 0] <= i_3_cast7_fu_121_p1[30 : 0];
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln116_reg_150 == 1'd1) & (1'b1 == ap_CS_fsm_state2))) begin
        icmp_ln117_reg_174 <= icmp_ln117_fu_127_p2;
    end
end

always @ (*) begin
    if ((ap_start_int == 1'b0)) begin
        ap_ST_fsm_state1_blk = 1'b1;
    end else begin
        ap_ST_fsm_state1_blk = 1'b0;
    end
end

assign ap_ST_fsm_state2_blk = 1'b0;

assign ap_ST_fsm_state3_blk = 1'b0;

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state3) & ((icmp_ln116_reg_150 == 1'd0) | ((icmp_ln117_reg_174 == 1'd0) | (icmp_ln117_1_fu_133_p2 == 1'd0))))) begin
        ap_condition_exit_pp0_iter0_stage2 = 1'b1;
    end else begin
        ap_condition_exit_pp0_iter0_stage2 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_loop_exit_ready == 1'b1) & (1'b1 == ap_CS_fsm_state3))) begin
        ap_done_int = 1'b1;
    end else begin
        ap_done_int = ap_done_reg;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start_int == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln116_reg_150 == 1'd1) & (icmp_ln117_reg_174 == 1'd1) & (icmp_ln117_1_fu_133_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state3))) begin
        ap_phi_mux_merge_phi_fu_90_p6 = 2'd1;
    end else begin
        ap_phi_mux_merge_phi_fu_90_p6 = merge_reg_85;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        ap_ready_int = 1'b1;
    end else begin
        ap_ready_int = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state3) & ((icmp_ln116_reg_150 == 1'd0) | ((icmp_ln117_reg_174 == 1'd0) | (icmp_ln117_1_fu_133_p2 == 1'd0))))) begin
        ap_return = ap_phi_mux_merge_phi_fu_90_p6;
    end else begin
        ap_return = ap_return_preg;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_loop_init == 1'b1))) begin
        ap_sig_allocacmp_i_1 = 31'd0;
    end else begin
        ap_sig_allocacmp_i_1 = i_fu_36;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start_int == 1'b1))) begin
        centroid_x_coords_ce0 = 1'b1;
    end else begin
        centroid_x_coords_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln116_reg_150 == 1'd1) & (1'b1 == ap_CS_fsm_state2) & (icmp_ln117_fu_127_p2 == 1'd1))) begin
        centroid_x_coords_prev_address0 = centroid_x_coords_prev_addr_reg_164;
    end else if (((icmp_ln116_fu_109_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1))) begin
        centroid_x_coords_prev_address0 = i_3_cast7_fu_121_p1;
    end else begin
        centroid_x_coords_prev_address0 = 'bx;
    end
end

always @ (*) begin
    if ((((icmp_ln116_reg_150 == 1'd1) & (1'b1 == ap_CS_fsm_state2) & (icmp_ln117_fu_127_p2 == 1'd1)) | ((icmp_ln116_fu_109_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state1) & (ap_start_int == 1'b1)))) begin
        centroid_x_coords_prev_ce0 = 1'b1;
    end else begin
        centroid_x_coords_prev_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        centroid_y_coords_ce0 = 1'b1;
    end else begin
        centroid_y_coords_ce0 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if (((1'b1 == ap_CS_fsm_state1) & (ap_start_int == 1'b1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            ap_NS_fsm = ap_ST_fsm_state3;
        end
        ap_ST_fsm_state3 : begin
            ap_NS_fsm = ap_ST_fsm_state1;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln116_fu_115_p2 = (ap_sig_allocacmp_i_1 + 31'd1);

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

always @ (*) begin
    ap_block_state1_pp0_stage0_iter0 = (ap_start_int == 1'b0);
end

assign ap_block_state2_pp0_stage1_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage2_iter0 = ~(1'b1 == 1'b1);

assign ap_loop_exit_ready = ap_condition_exit_pp0_iter0_stage2;

assign centroid_x_coords_address0 = i_3_cast7_fu_121_p1;

assign centroid_y_coords_address0 = i_3_cast7_reg_159;

assign i_3_cast7_fu_121_p1 = ap_sig_allocacmp_i_1;

assign icmp_ln116_fu_109_p2 = ((ap_sig_allocacmp_i_1 < k) ? 1'b1 : 1'b0);

assign icmp_ln117_1_fu_133_p2 = ((centroid_x_coords_prev_q0 == centroid_y_coords_q0) ? 1'b1 : 1'b0);

assign icmp_ln117_fu_127_p2 = ((centroid_x_coords_prev_q0 == centroid_x_coords_q0) ? 1'b1 : 1'b0);

always @ (posedge ap_clk) begin
    i_3_cast7_reg_159[63:31] <= 33'b000000000000000000000000000000000;
end

endmodule //kmeans_top_kmeans_Pipeline_VITIS_LOOP_116_6


// Content from kmeans_top_kmeans_top_Pipeline_10.v
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2022.2 (64-bit)
// Version: 2022.2
// Copyright (C) Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module kmeans_top_kmeans_top_Pipeline_10 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        m_axi_mem_AWVALID,
        m_axi_mem_AWREADY,
        m_axi_mem_AWADDR,
        m_axi_mem_AWID,
        m_axi_mem_AWLEN,
        m_axi_mem_AWSIZE,
        m_axi_mem_AWBURST,
        m_axi_mem_AWLOCK,
        m_axi_mem_AWCACHE,
        m_axi_mem_AWPROT,
        m_axi_mem_AWQOS,
        m_axi_mem_AWREGION,
        m_axi_mem_AWUSER,
        m_axi_mem_WVALID,
        m_axi_mem_WREADY,
        m_axi_mem_WDATA,
        m_axi_mem_WSTRB,
        m_axi_mem_WLAST,
        m_axi_mem_WID,
        m_axi_mem_WUSER,
        m_axi_mem_ARVALID,
        m_axi_mem_ARREADY,
        m_axi_mem_ARADDR,
        m_axi_mem_ARID,
        m_axi_mem_ARLEN,
        m_axi_mem_ARSIZE,
        m_axi_mem_ARBURST,
        m_axi_mem_ARLOCK,
        m_axi_mem_ARCACHE,
        m_axi_mem_ARPROT,
        m_axi_mem_ARQOS,
        m_axi_mem_ARREGION,
        m_axi_mem_ARUSER,
        m_axi_mem_RVALID,
        m_axi_mem_RREADY,
        m_axi_mem_RDATA,
        m_axi_mem_RLAST,
        m_axi_mem_RID,
        m_axi_mem_RFIFONUM,
        m_axi_mem_RUSER,
        m_axi_mem_RRESP,
        m_axi_mem_BVALID,
        m_axi_mem_BREADY,
        m_axi_mem_BRESP,
        m_axi_mem_BID,
        m_axi_mem_BUSER,
        p_cast8_cast,
        node_y_coords_address0,
        node_y_coords_ce0,
        node_y_coords_q0,
        sext_ln182
);

parameter    ap_ST_fsm_pp0_stage0 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
output   m_axi_mem_AWVALID;
input   m_axi_mem_AWREADY;
output  [63:0] m_axi_mem_AWADDR;
output  [0:0] m_axi_mem_AWID;
output  [31:0] m_axi_mem_AWLEN;
output  [2:0] m_axi_mem_AWSIZE;
output  [1:0] m_axi_mem_AWBURST;
output  [1:0] m_axi_mem_AWLOCK;
output  [3:0] m_axi_mem_AWCACHE;
output  [2:0] m_axi_mem_AWPROT;
output  [3:0] m_axi_mem_AWQOS;
output  [3:0] m_axi_mem_AWREGION;
output  [0:0] m_axi_mem_AWUSER;
output   m_axi_mem_WVALID;
input   m_axi_mem_WREADY;
output  [63:0] m_axi_mem_WDATA;
output  [7:0] m_axi_mem_WSTRB;
output   m_axi_mem_WLAST;
output  [0:0] m_axi_mem_WID;
output  [0:0] m_axi_mem_WUSER;
output   m_axi_mem_ARVALID;
input   m_axi_mem_ARREADY;
output  [63:0] m_axi_mem_ARADDR;
output  [0:0] m_axi_mem_ARID;
output  [31:0] m_axi_mem_ARLEN;
output  [2:0] m_axi_mem_ARSIZE;
output  [1:0] m_axi_mem_ARBURST;
output  [1:0] m_axi_mem_ARLOCK;
output  [3:0] m_axi_mem_ARCACHE;
output  [2:0] m_axi_mem_ARPROT;
output  [3:0] m_axi_mem_ARQOS;
output  [3:0] m_axi_mem_ARREGION;
output  [0:0] m_axi_mem_ARUSER;
input   m_axi_mem_RVALID;
output   m_axi_mem_RREADY;
input  [63:0] m_axi_mem_RDATA;
input   m_axi_mem_RLAST;
input  [0:0] m_axi_mem_RID;
input  [8:0] m_axi_mem_RFIFONUM;
input  [0:0] m_axi_mem_RUSER;
input  [1:0] m_axi_mem_RRESP;
input   m_axi_mem_BVALID;
output   m_axi_mem_BREADY;
input  [1:0] m_axi_mem_BRESP;
input  [0:0] m_axi_mem_BID;
input  [0:0] m_axi_mem_BUSER;
input  [60:0] p_cast8_cast;
output  [12:0] node_y_coords_address0;
output   node_y_coords_ce0;
input  [63:0] node_y_coords_q0;
input  [31:0] sext_ln182;

reg ap_idle;
reg m_axi_mem_WVALID;
reg node_y_coords_ce0;

(* fsm_encoding = "none" *) reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_enable_reg_pp0_iter0;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter2;
reg    ap_enable_reg_pp0_iter3;
reg    ap_idle_pp0;
wire    ap_block_state1_pp0_stage0_iter0;
wire    ap_block_state2_pp0_stage0_iter1;
wire    ap_block_state3_pp0_stage0_iter2;
wire    ap_block_state4_pp0_stage0_iter3;
reg    ap_block_pp0_stage0_subdone;
wire   [0:0] exitcond76_fu_126_p2;
reg    ap_condition_exit_pp0_iter1_stage0;
wire    ap_loop_exit_ready;
reg    ap_ready_int;
reg    mem_blk_n_W;
wire    ap_block_pp0_stage0;
wire  signed [60:0] sext_ln182_cast_fu_99_p1;
reg  signed [60:0] sext_ln182_cast_reg_149;
reg    ap_block_pp0_stage0_11001;
reg   [63:0] node_y_coords_load_reg_168;
wire   [63:0] loop_index15_cast_fu_121_p1;
wire    ap_block_pp0_stage0_01001;
reg   [60:0] loop_index15_fu_62;
wire   [60:0] empty_fu_115_p2;
wire    ap_loop_init;
reg    ap_done_reg;
wire    ap_continue_int;
reg    ap_done_int;
reg    ap_loop_exit_ready_pp0_iter2_reg;
reg    ap_loop_exit_ready_pp0_iter3_reg;
reg   [0:0] ap_NS_fsm;
wire    ap_enable_pp0;
wire    ap_start_int;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_CS_fsm = 1'd1;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_done_reg = 1'b0;
end

kmeans_top_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(ap_start),
    .ap_ready(ap_ready),
    .ap_done(ap_done),
    .ap_start_int(ap_start_int),
    .ap_loop_init(ap_loop_init),
    .ap_ready_int(ap_ready_int),
    .ap_loop_exit_ready(ap_condition_exit_pp0_iter1_stage0),
    .ap_loop_exit_done(ap_done_int),
    .ap_continue_int(ap_continue_int),
    .ap_done_int(ap_done_int)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue_int == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter3_reg == 1'b1))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b1 == ap_condition_exit_pp0_iter1_stage0)) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_enable_reg_pp0_iter1 <= ap_start_int;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter2_reg == 1'b0))) begin
        ap_loop_exit_ready_pp0_iter3_reg <= 1'b0;
    end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        ap_loop_exit_ready_pp0_iter3_reg <= ap_loop_exit_ready_pp0_iter2_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        if ((ap_loop_init == 1'b1)) begin
            loop_index15_fu_62 <= 61'd0;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (exitcond76_fu_126_p2 == 1'd0))) begin
            loop_index15_fu_62 <= empty_fu_115_p2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_loop_exit_ready_pp0_iter2_reg <= ap_loop_exit_ready;
        sext_ln182_cast_reg_149 <= sext_ln182_cast_fu_99_p1;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        node_y_coords_load_reg_168 <= node_y_coords_q0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (exitcond76_fu_126_p2 == 1'd1))) begin
        ap_condition_exit_pp0_iter1_stage0 = 1'b1;
    end else begin
        ap_condition_exit_pp0_iter1_stage0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter3_reg == 1'b1))) begin
        ap_done_int = 1'b1;
    end else begin
        ap_done_int = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_idle_pp0 == 1'b1) & (ap_start_int == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_ready_int = 1'b1;
    end else begin
        ap_ready_int = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1))) begin
        m_axi_mem_WVALID = 1'b1;
    end else begin
        m_axi_mem_WVALID = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter3 == 1'b1))) begin
        mem_blk_n_W = m_axi_mem_WREADY;
    end else begin
        mem_blk_n_W = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        node_y_coords_ce0 = 1'b1;
    end else begin
        node_y_coords_ce0 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_pp0_stage0 : begin
            ap_NS_fsm = ap_ST_fsm_pp0_stage0;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_01001 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_pp0_stage0_11001 = ((m_axi_mem_WREADY == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b1));
end

always @ (*) begin
    ap_block_pp0_stage0_subdone = ((m_axi_mem_WREADY == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b1));
end

assign ap_block_state1_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_enable_reg_pp0_iter0 = ap_start_int;

assign ap_loop_exit_ready = ap_condition_exit_pp0_iter1_stage0;

assign empty_fu_115_p2 = (loop_index15_fu_62 + 61'd1);

assign exitcond76_fu_126_p2 = ((empty_fu_115_p2 == sext_ln182_cast_reg_149) ? 1'b1 : 1'b0);

assign loop_index15_cast_fu_121_p1 = loop_index15_fu_62;

assign m_axi_mem_ARADDR = 64'd0;

assign m_axi_mem_ARBURST = 2'd0;

assign m_axi_mem_ARCACHE = 4'd0;

assign m_axi_mem_ARID = 1'd0;

assign m_axi_mem_ARLEN = 32'd0;

assign m_axi_mem_ARLOCK = 2'd0;

assign m_axi_mem_ARPROT = 3'd0;

assign m_axi_mem_ARQOS = 4'd0;

assign m_axi_mem_ARREGION = 4'd0;

assign m_axi_mem_ARSIZE = 3'd0;

assign m_axi_mem_ARUSER = 1'd0;

assign m_axi_mem_ARVALID = 1'b0;

assign m_axi_mem_AWADDR = 64'd0;

assign m_axi_mem_AWBURST = 2'd0;

assign m_axi_mem_AWCACHE = 4'd0;

assign m_axi_mem_AWID = 1'd0;

assign m_axi_mem_AWLEN = 32'd0;

assign m_axi_mem_AWLOCK = 2'd0;

assign m_axi_mem_AWPROT = 3'd0;

assign m_axi_mem_AWQOS = 4'd0;

assign m_axi_mem_AWREGION = 4'd0;

assign m_axi_mem_AWSIZE = 3'd0;

assign m_axi_mem_AWUSER = 1'd0;

assign m_axi_mem_AWVALID = 1'b0;

assign m_axi_mem_BREADY = 1'b0;

assign m_axi_mem_RREADY = 1'b0;

assign m_axi_mem_WDATA = node_y_coords_load_reg_168;

assign m_axi_mem_WID = 1'd0;

assign m_axi_mem_WLAST = 1'b0;

assign m_axi_mem_WSTRB = 8'd255;

assign m_axi_mem_WUSER = 1'd0;

assign node_y_coords_address0 = loop_index15_cast_fu_121_p1;

assign sext_ln182_cast_fu_99_p1 = $signed(sext_ln182);

endmodule //kmeans_top_kmeans_top_Pipeline_10


// Content from kmeans_top_kmeans_top_Pipeline_11.v
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2022.2 (64-bit)
// Version: 2022.2
// Copyright (C) Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module kmeans_top_kmeans_top_Pipeline_11 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        m_axi_mem_AWVALID,
        m_axi_mem_AWREADY,
        m_axi_mem_AWADDR,
        m_axi_mem_AWID,
        m_axi_mem_AWLEN,
        m_axi_mem_AWSIZE,
        m_axi_mem_AWBURST,
        m_axi_mem_AWLOCK,
        m_axi_mem_AWCACHE,
        m_axi_mem_AWPROT,
        m_axi_mem_AWQOS,
        m_axi_mem_AWREGION,
        m_axi_mem_AWUSER,
        m_axi_mem_WVALID,
        m_axi_mem_WREADY,
        m_axi_mem_WDATA,
        m_axi_mem_WSTRB,
        m_axi_mem_WLAST,
        m_axi_mem_WID,
        m_axi_mem_WUSER,
        m_axi_mem_ARVALID,
        m_axi_mem_ARREADY,
        m_axi_mem_ARADDR,
        m_axi_mem_ARID,
        m_axi_mem_ARLEN,
        m_axi_mem_ARSIZE,
        m_axi_mem_ARBURST,
        m_axi_mem_ARLOCK,
        m_axi_mem_ARCACHE,
        m_axi_mem_ARPROT,
        m_axi_mem_ARQOS,
        m_axi_mem_ARREGION,
        m_axi_mem_ARUSER,
        m_axi_mem_RVALID,
        m_axi_mem_RREADY,
        m_axi_mem_RDATA,
        m_axi_mem_RLAST,
        m_axi_mem_RID,
        m_axi_mem_RFIFONUM,
        m_axi_mem_RUSER,
        m_axi_mem_RRESP,
        m_axi_mem_BVALID,
        m_axi_mem_BREADY,
        m_axi_mem_BRESP,
        m_axi_mem_BID,
        m_axi_mem_BUSER,
        p_cast6_cast,
        node_cluster_assignments_address0,
        node_cluster_assignments_ce0,
        node_cluster_assignments_q0,
        sext_ln182
);

parameter    ap_ST_fsm_pp0_stage0 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
output   m_axi_mem_AWVALID;
input   m_axi_mem_AWREADY;
output  [63:0] m_axi_mem_AWADDR;
output  [0:0] m_axi_mem_AWID;
output  [31:0] m_axi_mem_AWLEN;
output  [2:0] m_axi_mem_AWSIZE;
output  [1:0] m_axi_mem_AWBURST;
output  [1:0] m_axi_mem_AWLOCK;
output  [3:0] m_axi_mem_AWCACHE;
output  [2:0] m_axi_mem_AWPROT;
output  [3:0] m_axi_mem_AWQOS;
output  [3:0] m_axi_mem_AWREGION;
output  [0:0] m_axi_mem_AWUSER;
output   m_axi_mem_WVALID;
input   m_axi_mem_WREADY;
output  [63:0] m_axi_mem_WDATA;
output  [7:0] m_axi_mem_WSTRB;
output   m_axi_mem_WLAST;
output  [0:0] m_axi_mem_WID;
output  [0:0] m_axi_mem_WUSER;
output   m_axi_mem_ARVALID;
input   m_axi_mem_ARREADY;
output  [63:0] m_axi_mem_ARADDR;
output  [0:0] m_axi_mem_ARID;
output  [31:0] m_axi_mem_ARLEN;
output  [2:0] m_axi_mem_ARSIZE;
output  [1:0] m_axi_mem_ARBURST;
output  [1:0] m_axi_mem_ARLOCK;
output  [3:0] m_axi_mem_ARCACHE;
output  [2:0] m_axi_mem_ARPROT;
output  [3:0] m_axi_mem_ARQOS;
output  [3:0] m_axi_mem_ARREGION;
output  [0:0] m_axi_mem_ARUSER;
input   m_axi_mem_RVALID;
output   m_axi_mem_RREADY;
input  [63:0] m_axi_mem_RDATA;
input   m_axi_mem_RLAST;
input  [0:0] m_axi_mem_RID;
input  [8:0] m_axi_mem_RFIFONUM;
input  [0:0] m_axi_mem_RUSER;
input  [1:0] m_axi_mem_RRESP;
input   m_axi_mem_BVALID;
output   m_axi_mem_BREADY;
input  [1:0] m_axi_mem_BRESP;
input  [0:0] m_axi_mem_BID;
input  [0:0] m_axi_mem_BUSER;
input  [60:0] p_cast6_cast;
output  [12:0] node_cluster_assignments_address0;
output   node_cluster_assignments_ce0;
input  [63:0] node_cluster_assignments_q0;
input  [31:0] sext_ln182;

reg ap_idle;
reg m_axi_mem_WVALID;
reg node_cluster_assignments_ce0;

(* fsm_encoding = "none" *) reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_enable_reg_pp0_iter0;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter2;
reg    ap_enable_reg_pp0_iter3;
reg    ap_idle_pp0;
wire    ap_block_state1_pp0_stage0_iter0;
wire    ap_block_state2_pp0_stage0_iter1;
wire    ap_block_state3_pp0_stage0_iter2;
wire    ap_block_state4_pp0_stage0_iter3;
reg    ap_block_pp0_stage0_subdone;
wire   [0:0] exitcond75_fu_126_p2;
reg    ap_condition_exit_pp0_iter1_stage0;
wire    ap_loop_exit_ready;
reg    ap_ready_int;
reg    mem_blk_n_W;
wire    ap_block_pp0_stage0;
wire  signed [60:0] sext_ln182_cast_fu_99_p1;
reg  signed [60:0] sext_ln182_cast_reg_149;
reg    ap_block_pp0_stage0_11001;
reg   [63:0] node_cluster_assignments_load_reg_168;
wire   [63:0] loop_index9_cast_fu_121_p1;
wire    ap_block_pp0_stage0_01001;
reg   [60:0] loop_index9_fu_62;
wire   [60:0] empty_fu_115_p2;
wire    ap_loop_init;
reg    ap_done_reg;
wire    ap_continue_int;
reg    ap_done_int;
reg    ap_loop_exit_ready_pp0_iter2_reg;
reg    ap_loop_exit_ready_pp0_iter3_reg;
reg   [0:0] ap_NS_fsm;
wire    ap_enable_pp0;
wire    ap_start_int;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_CS_fsm = 1'd1;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_done_reg = 1'b0;
end

kmeans_top_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(ap_start),
    .ap_ready(ap_ready),
    .ap_done(ap_done),
    .ap_start_int(ap_start_int),
    .ap_loop_init(ap_loop_init),
    .ap_ready_int(ap_ready_int),
    .ap_loop_exit_ready(ap_condition_exit_pp0_iter1_stage0),
    .ap_loop_exit_done(ap_done_int),
    .ap_continue_int(ap_continue_int),
    .ap_done_int(ap_done_int)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue_int == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter3_reg == 1'b1))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b1 == ap_condition_exit_pp0_iter1_stage0)) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_enable_reg_pp0_iter1 <= ap_start_int;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter2_reg == 1'b0))) begin
        ap_loop_exit_ready_pp0_iter3_reg <= 1'b0;
    end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        ap_loop_exit_ready_pp0_iter3_reg <= ap_loop_exit_ready_pp0_iter2_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        if ((ap_loop_init == 1'b1)) begin
            loop_index9_fu_62 <= 61'd0;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (exitcond75_fu_126_p2 == 1'd0))) begin
            loop_index9_fu_62 <= empty_fu_115_p2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_loop_exit_ready_pp0_iter2_reg <= ap_loop_exit_ready;
        sext_ln182_cast_reg_149 <= sext_ln182_cast_fu_99_p1;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        node_cluster_assignments_load_reg_168 <= node_cluster_assignments_q0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (exitcond75_fu_126_p2 == 1'd1))) begin
        ap_condition_exit_pp0_iter1_stage0 = 1'b1;
    end else begin
        ap_condition_exit_pp0_iter1_stage0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter3_reg == 1'b1))) begin
        ap_done_int = 1'b1;
    end else begin
        ap_done_int = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_idle_pp0 == 1'b1) & (ap_start_int == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_ready_int = 1'b1;
    end else begin
        ap_ready_int = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1))) begin
        m_axi_mem_WVALID = 1'b1;
    end else begin
        m_axi_mem_WVALID = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter3 == 1'b1))) begin
        mem_blk_n_W = m_axi_mem_WREADY;
    end else begin
        mem_blk_n_W = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        node_cluster_assignments_ce0 = 1'b1;
    end else begin
        node_cluster_assignments_ce0 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_pp0_stage0 : begin
            ap_NS_fsm = ap_ST_fsm_pp0_stage0;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_01001 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_pp0_stage0_11001 = ((m_axi_mem_WREADY == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b1));
end

always @ (*) begin
    ap_block_pp0_stage0_subdone = ((m_axi_mem_WREADY == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b1));
end

assign ap_block_state1_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_enable_reg_pp0_iter0 = ap_start_int;

assign ap_loop_exit_ready = ap_condition_exit_pp0_iter1_stage0;

assign empty_fu_115_p2 = (loop_index9_fu_62 + 61'd1);

assign exitcond75_fu_126_p2 = ((empty_fu_115_p2 == sext_ln182_cast_reg_149) ? 1'b1 : 1'b0);

assign loop_index9_cast_fu_121_p1 = loop_index9_fu_62;

assign m_axi_mem_ARADDR = 64'd0;

assign m_axi_mem_ARBURST = 2'd0;

assign m_axi_mem_ARCACHE = 4'd0;

assign m_axi_mem_ARID = 1'd0;

assign m_axi_mem_ARLEN = 32'd0;

assign m_axi_mem_ARLOCK = 2'd0;

assign m_axi_mem_ARPROT = 3'd0;

assign m_axi_mem_ARQOS = 4'd0;

assign m_axi_mem_ARREGION = 4'd0;

assign m_axi_mem_ARSIZE = 3'd0;

assign m_axi_mem_ARUSER = 1'd0;

assign m_axi_mem_ARVALID = 1'b0;

assign m_axi_mem_AWADDR = 64'd0;

assign m_axi_mem_AWBURST = 2'd0;

assign m_axi_mem_AWCACHE = 4'd0;

assign m_axi_mem_AWID = 1'd0;

assign m_axi_mem_AWLEN = 32'd0;

assign m_axi_mem_AWLOCK = 2'd0;

assign m_axi_mem_AWPROT = 3'd0;

assign m_axi_mem_AWQOS = 4'd0;

assign m_axi_mem_AWREGION = 4'd0;

assign m_axi_mem_AWSIZE = 3'd0;

assign m_axi_mem_AWUSER = 1'd0;

assign m_axi_mem_AWVALID = 1'b0;

assign m_axi_mem_BREADY = 1'b0;

assign m_axi_mem_RREADY = 1'b0;

assign m_axi_mem_WDATA = node_cluster_assignments_load_reg_168;

assign m_axi_mem_WID = 1'd0;

assign m_axi_mem_WLAST = 1'b0;

assign m_axi_mem_WSTRB = 8'd255;

assign m_axi_mem_WUSER = 1'd0;

assign node_cluster_assignments_address0 = loop_index9_cast_fu_121_p1;

assign sext_ln182_cast_fu_99_p1 = $signed(sext_ln182);

endmodule //kmeans_top_kmeans_top_Pipeline_11


// Content from kmeans_top_kmeans_cluster_cardinality_next_RAM_AUTO_1R1W.v
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2022.2 (64-bit)
// Version: 2022.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module kmeans_top_kmeans_cluster_cardinality_next_RAM_AUTO_1R1W (
     
    address0, ce0,
    d0, we0, 
    q0, 
     
    reset, clk);

parameter DataWidth = 16;
parameter AddressWidth = 8;
parameter AddressRange = 256;
 
input[AddressWidth-1:0] address0;
input ce0;
input[DataWidth-1:0] d0;
input we0; 
output reg[DataWidth-1:0] q0; 

input reset;
input clk;

(* ram_style = "auto"  *)reg [DataWidth-1:0] ram[0:AddressRange-1];


 





//read first
always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[address0] <= d0; 
        q0 <= ram[address0];

    end
end 
 
 

endmodule



// Content from kmeans_top_flow_control_loop_pipe_sequential_init.v
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2022.2 (64-bit)
// Tool Version Limit: 2019.12
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module kmeans_top_flow_control_loop_pipe_sequential_init(
        ap_clk,
        ap_rst,
        ap_start,
        ap_ready,
        ap_done,
        ap_start_int,
        ap_ready_int,
        ap_done_int,
        ap_continue_int,
        ap_loop_init,
        ap_loop_exit_ready,
        ap_loop_exit_done
);

input   ap_clk;
input   ap_rst;

//Block level handshake with outside loop
input   ap_start;
output  ap_ready;
output  ap_done;

//Block level handshake with loop body
output  ap_start_int;
input   ap_ready_int;
input   ap_done_int;
output  ap_continue_int;

//Init live in variables
output   ap_loop_init;
wire     ap_loop_init;
reg ap_loop_init_int;
reg ap_done;
reg ap_done_cache;

//Exit signal from loop body
input   ap_loop_exit_ready;
input   ap_loop_exit_done;

// power-on initialization
initial begin
#0 ap_loop_init_int = 1'b1;
#0 ap_done_cache = 1'b0;
end

assign ap_start_int = ap_start;

assign ap_continue_int = 1'b1;

assign ap_ready = ap_loop_exit_ready;

//ap_loop_init is valid for the first II
//of the first loop run so as to enable
//the init block ops which are pushed into
//the first state of the pipeline region
always @ (posedge ap_clk)
begin
    if (ap_rst == 1'b1) begin
        ap_loop_init_int <= 1'b1;
    end else if(ap_loop_exit_done == 1'b1) begin
        ap_loop_init_int <= 1'b1;
    end else if(ap_ready_int == 1'b1) begin
        ap_loop_init_int <= 1'b0;
    end
end

assign ap_loop_init = ap_loop_init_int & ap_start;

// if no ap_continue port and current module is not top module, 
// ap_done handshakes with ap_start. Internally, flow control sends out 
// ap_conintue_int = 1'b1 so the ap_done_int is asserted high for 1 clock cycle.
// ap_done_cache is used to record ap_done_int, and de-assert if ap_start_int
// is asserted, so DUT can start the next run
always @(posedge ap_clk)
begin
    if (ap_rst == 1'b1) begin
        ap_done_cache <= 1'b0;
    end else if (ap_done_int == 1'b1) begin
        ap_done_cache <= 1'b1;
    end else if (ap_start_int == 1'b1) begin
        ap_done_cache <= 1'b0;
    end
end

// if no ap_continue port and current module is not top module, ap_done handshakes with ap_start
always @(*)
begin
    if ((ap_done_int == 1'b1) || ((ap_done_cache == 1'b1) && (ap_start_int == 1'b0))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

endmodule
        


// Content from kmeans_top_node_x_coords_RAM_2P_URAM_1R1W.v
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2022.2 (64-bit)
// Version: 2022.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module kmeans_top_node_x_coords_RAM_2P_URAM_1R1W (
     
    address0, ce0,
    
    q0, 
      
    address1, ce1,
    d1, we1, 
    q1, 
     
    reset, clk);

parameter DataWidth = 64;
parameter AddressWidth = 13;
parameter AddressRange = 8192;
 
input[AddressWidth-1:0] address0;
input ce0;

output reg[DataWidth-1:0] q0; 
  
input[AddressWidth-1:0] address1;
input ce1;
input[DataWidth-1:0] d1;
input we1; 
output reg[DataWidth-1:0] q1; 
 
input reset;
input clk;

(* ram_style = "hls_ultra" , cascade_height = 1 *)reg [DataWidth-1:0] ram[0:AddressRange-1];


 



always @(posedge clk) 
begin 
    if (ce0) begin
        q0 <= ram[address0];
    end
end 

 
  






always @(posedge clk)  
begin 
    if (ce1) begin
        if (we1) 
            ram[address1] <= d1; 
        else 
            q1 <= ram[address1];
    end
end 
 
 

endmodule



// Content from kmeans_top_udiv_64ns_16ns_64_68_seq_1.v
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2022.2 (64-bit)
// Version: 2022.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps

module kmeans_top_udiv_64ns_16ns_64_68_seq_1_divseq
#(parameter
    in0_WIDTH = 32,
    in1_WIDTH = 32,
    out_WIDTH = 32
)
(
    input                       clk,
    input                       reset,
    input                       ce,
    input                       start,
    input       [in0_WIDTH-1:0] dividend,
    input       [in1_WIDTH-1:0] divisor,
    output wire                 done,
    output wire [out_WIDTH-1:0] quot,
    output wire [out_WIDTH-1:0] remd
);

localparam cal_WIDTH = (in0_WIDTH > in1_WIDTH)? in0_WIDTH : in1_WIDTH;

//------------------------Local signal-------------------
reg     [in0_WIDTH-1:0] dividend0;
reg     [in1_WIDTH-1:0] divisor0;
reg     [in0_WIDTH-1:0] dividend_tmp;
reg     [in0_WIDTH-1:0] remd_tmp;
wire    [in0_WIDTH-1:0] dividend_tmp_mux;
wire    [in0_WIDTH-1:0] remd_tmp_mux;
wire    [in0_WIDTH-1:0] comb_tmp;
wire    [cal_WIDTH:0]   cal_tmp;

//------------------------Body---------------------------
assign  quot   = dividend_tmp;
assign  remd   = remd_tmp;

// dividend0, divisor0
always @(posedge clk)
begin
    if (start) begin
        dividend0 <= dividend;
        divisor0  <= divisor;
    end
end

// One-Hot Register
// r_stage[0]=1:accept input; r_stage[in0_WIDTH]=1:done
reg     [in0_WIDTH:0]     r_stage;
assign done = r_stage[in0_WIDTH];
always @(posedge clk)
begin
    if (reset == 1'b1)
        r_stage[in0_WIDTH:0] <= {in0_WIDTH{1'b0}};
    else if (ce)
        r_stage[in0_WIDTH:0] <= {r_stage[in0_WIDTH-1:0], start};
end

// MUXs
assign  dividend_tmp_mux = r_stage[0]? dividend0 : dividend_tmp;
assign  remd_tmp_mux     = r_stage[0]? {in0_WIDTH{1'b0}} : remd_tmp;

if (in0_WIDTH == 1) assign comb_tmp = dividend_tmp_mux[0];
else                assign comb_tmp = {remd_tmp_mux[in0_WIDTH-2:0], dividend_tmp_mux[in0_WIDTH-1]};

assign  cal_tmp  = {1'b0, comb_tmp} - {1'b0, divisor0};

always @(posedge clk)
begin
    if (ce) begin
        if (in0_WIDTH == 1) dividend_tmp <= ~cal_tmp[cal_WIDTH];
        else           dividend_tmp <= {dividend_tmp_mux[in0_WIDTH-2:0], ~cal_tmp[cal_WIDTH]};
        remd_tmp     <= cal_tmp[cal_WIDTH]? comb_tmp : cal_tmp[in0_WIDTH-1:0];
    end
end

endmodule

module kmeans_top_udiv_64ns_16ns_64_68_seq_1
#(parameter
        ID   = 1,
        NUM_STAGE   = 2,
        din0_WIDTH   = 32,
        din1_WIDTH   = 32,
        dout_WIDTH   = 32
)
(
        input                           clk,
        input                           reset,
        input                           ce,
        input                           start,
        output  reg                     done,
        input           [din0_WIDTH-1:0] din0,
        input           [din1_WIDTH-1:0] din1,
        output          [dout_WIDTH-1:0] dout
);
//------------------------Local signal-------------------
reg                       start0 = 'b0;
wire                      done0;
reg     [din0_WIDTH-1:0] dividend0;
reg     [din1_WIDTH-1:0] divisor0;
wire    [din0_WIDTH-1:0] dividend_u;
wire    [din1_WIDTH-1:0] divisor_u;
wire    [dout_WIDTH-1:0] quot_u;
wire    [dout_WIDTH-1:0] remd_u;
reg     [dout_WIDTH-1:0] quot;
reg     [dout_WIDTH-1:0] remd;
//------------------------Instantiation------------------
kmeans_top_udiv_64ns_16ns_64_68_seq_1_divseq #(
    .in0_WIDTH      ( din0_WIDTH ),
    .in1_WIDTH      ( din1_WIDTH ),
    .out_WIDTH      ( dout_WIDTH )
) kmeans_top_udiv_64ns_16ns_64_68_seq_1_divseq_u (
    .clk      ( clk ),
    .reset    ( reset ),
    .ce       ( ce ),
    .start    ( start0 ),
    .done     ( done0 ),
    .dividend ( dividend_u ),
    .divisor  ( divisor_u ),
    .quot     ( quot_u ),
    .remd     ( remd_u )
);
//------------------------Body---------------------------
assign dividend_u = dividend0;
assign divisor_u = divisor0;

always @(posedge clk)
begin
    if (ce) begin
        dividend0 <= din0;
        divisor0  <= din1;
        start0    <= start;
    end
end

always @(posedge clk)
begin
    done <= done0;
end

always @(posedge clk)
begin
    if (done0) begin
        quot <= quot_u;
        remd <= remd_u;
    end
end

assign dout = quot;

endmodule




// Content from kmeans_top_kmeans_Pipeline_4.v
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2022.2 (64-bit)
// Version: 2022.2
// Copyright (C) Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module kmeans_top_kmeans_Pipeline_4 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        centroid_y_coords_next_address0,
        centroid_y_coords_next_ce0,
        centroid_y_coords_next_we0,
        centroid_y_coords_next_d0,
        k_cast2_cast_cast
);

parameter    ap_ST_fsm_pp0_stage0 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
output  [7:0] centroid_y_coords_next_address0;
output   centroid_y_coords_next_ce0;
output   centroid_y_coords_next_we0;
output  [63:0] centroid_y_coords_next_d0;
input  [31:0] k_cast2_cast_cast;

reg ap_idle;
reg centroid_y_coords_next_ce0;
reg centroid_y_coords_next_we0;

(* fsm_encoding = "none" *) reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_enable_reg_pp0_iter0;
reg    ap_enable_reg_pp0_iter1;
reg    ap_idle_pp0;
wire    ap_block_state1_pp0_stage0_iter0;
wire    ap_block_state2_pp0_stage0_iter1;
wire    ap_block_pp0_stage0_subdone;
wire   [0:0] exitcond1_fu_71_p2;
reg    ap_condition_exit_pp0_iter1_stage0;
wire    ap_loop_exit_ready;
reg    ap_ready_int;
wire   [63:0] k_cast2_cast_cast_cast_cast_fu_52_p1;
reg   [63:0] k_cast2_cast_cast_cast_cast_reg_88;
wire    ap_block_pp0_stage0_11001;
wire    ap_block_pp0_stage0;
reg   [63:0] empty_fu_24;
wire   [63:0] empty_69_fu_65_p2;
wire    ap_loop_init;
wire  signed [60:0] k_cast2_cast_cast_cast_fu_48_p1;
reg    ap_done_reg;
wire    ap_continue_int;
reg    ap_done_int;
reg   [0:0] ap_NS_fsm;
wire    ap_enable_pp0;
wire    ap_start_int;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_CS_fsm = 1'd1;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_done_reg = 1'b0;
end

kmeans_top_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(ap_start),
    .ap_ready(ap_ready),
    .ap_done(ap_done),
    .ap_start_int(ap_start_int),
    .ap_loop_init(ap_loop_init),
    .ap_ready_int(ap_ready_int),
    .ap_loop_exit_ready(ap_condition_exit_pp0_iter1_stage0),
    .ap_loop_exit_done(ap_done_int),
    .ap_continue_int(ap_continue_int),
    .ap_done_int(ap_done_int)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue_int == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((ap_loop_exit_ready == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b1 == ap_condition_exit_pp0_iter1_stage0)) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_enable_reg_pp0_iter1 <= ap_start_int;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        if ((ap_loop_init == 1'b1)) begin
            empty_fu_24 <= 64'd0;
        end else if (((exitcond1_fu_71_p2 == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
            empty_fu_24 <= empty_69_fu_65_p2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        k_cast2_cast_cast_cast_cast_reg_88[60 : 0] <= k_cast2_cast_cast_cast_cast_fu_52_p1[60 : 0];
    end
end

always @ (*) begin
    if (((exitcond1_fu_71_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_condition_exit_pp0_iter1_stage0 = 1'b1;
    end else begin
        ap_condition_exit_pp0_iter1_stage0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_loop_exit_ready == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_done_int = 1'b1;
    end else begin
        ap_done_int = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_idle_pp0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_start_int == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_ready_int = 1'b1;
    end else begin
        ap_ready_int = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        centroid_y_coords_next_ce0 = 1'b1;
    end else begin
        centroid_y_coords_next_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        centroid_y_coords_next_we0 = 1'b1;
    end else begin
        centroid_y_coords_next_we0 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_pp0_stage0 : begin
            ap_NS_fsm = ap_ST_fsm_pp0_stage0;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

assign ap_block_state1_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_enable_reg_pp0_iter0 = ap_start_int;

assign ap_loop_exit_ready = ap_condition_exit_pp0_iter1_stage0;

assign centroid_y_coords_next_address0 = empty_fu_24;

assign centroid_y_coords_next_d0 = 64'd0;

assign empty_69_fu_65_p2 = (empty_fu_24 + 64'd1);

assign exitcond1_fu_71_p2 = ((empty_69_fu_65_p2 == k_cast2_cast_cast_cast_cast_reg_88) ? 1'b1 : 1'b0);

assign k_cast2_cast_cast_cast_cast_fu_52_p1 = $unsigned(k_cast2_cast_cast_cast_fu_48_p1);

assign k_cast2_cast_cast_cast_fu_48_p1 = $signed(k_cast2_cast_cast);

always @ (posedge ap_clk) begin
    k_cast2_cast_cast_cast_cast_reg_88[63:61] <= 3'b000;
end

endmodule //kmeans_top_kmeans_Pipeline_4


// Content from kmeans_top_mul_29s_29s_29_1_1.v
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2022.2 (64-bit)
// Version: 2022.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module kmeans_top_mul_29s_29s_29_1_1(din0, din1, dout);
parameter ID = 1;
parameter NUM_STAGE = 0;
parameter din0_WIDTH = 14;
parameter din1_WIDTH = 12;
parameter dout_WIDTH = 26;
input [din0_WIDTH - 1 : 0] din0; 
input [din1_WIDTH - 1 : 0] din1; 
output [dout_WIDTH - 1 : 0] dout;

assign dout = $signed(din0) * $signed(din1);
endmodule


// Content from kmeans_top_kmeans_top_Pipeline_13.v
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2022.2 (64-bit)
// Version: 2022.2
// Copyright (C) Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module kmeans_top_kmeans_top_Pipeline_13 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        m_axi_mem_AWVALID,
        m_axi_mem_AWREADY,
        m_axi_mem_AWADDR,
        m_axi_mem_AWID,
        m_axi_mem_AWLEN,
        m_axi_mem_AWSIZE,
        m_axi_mem_AWBURST,
        m_axi_mem_AWLOCK,
        m_axi_mem_AWCACHE,
        m_axi_mem_AWPROT,
        m_axi_mem_AWQOS,
        m_axi_mem_AWREGION,
        m_axi_mem_AWUSER,
        m_axi_mem_WVALID,
        m_axi_mem_WREADY,
        m_axi_mem_WDATA,
        m_axi_mem_WSTRB,
        m_axi_mem_WLAST,
        m_axi_mem_WID,
        m_axi_mem_WUSER,
        m_axi_mem_ARVALID,
        m_axi_mem_ARREADY,
        m_axi_mem_ARADDR,
        m_axi_mem_ARID,
        m_axi_mem_ARLEN,
        m_axi_mem_ARSIZE,
        m_axi_mem_ARBURST,
        m_axi_mem_ARLOCK,
        m_axi_mem_ARCACHE,
        m_axi_mem_ARPROT,
        m_axi_mem_ARQOS,
        m_axi_mem_ARREGION,
        m_axi_mem_ARUSER,
        m_axi_mem_RVALID,
        m_axi_mem_RREADY,
        m_axi_mem_RDATA,
        m_axi_mem_RLAST,
        m_axi_mem_RID,
        m_axi_mem_RFIFONUM,
        m_axi_mem_RUSER,
        m_axi_mem_RRESP,
        m_axi_mem_BVALID,
        m_axi_mem_BREADY,
        m_axi_mem_BRESP,
        m_axi_mem_BID,
        m_axi_mem_BUSER,
        p_cast12_cast,
        centroid_y_coords_address0,
        centroid_y_coords_ce0,
        centroid_y_coords_q0,
        sext_ln185
);

parameter    ap_ST_fsm_pp0_stage0 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
output   m_axi_mem_AWVALID;
input   m_axi_mem_AWREADY;
output  [63:0] m_axi_mem_AWADDR;
output  [0:0] m_axi_mem_AWID;
output  [31:0] m_axi_mem_AWLEN;
output  [2:0] m_axi_mem_AWSIZE;
output  [1:0] m_axi_mem_AWBURST;
output  [1:0] m_axi_mem_AWLOCK;
output  [3:0] m_axi_mem_AWCACHE;
output  [2:0] m_axi_mem_AWPROT;
output  [3:0] m_axi_mem_AWQOS;
output  [3:0] m_axi_mem_AWREGION;
output  [0:0] m_axi_mem_AWUSER;
output   m_axi_mem_WVALID;
input   m_axi_mem_WREADY;
output  [63:0] m_axi_mem_WDATA;
output  [7:0] m_axi_mem_WSTRB;
output   m_axi_mem_WLAST;
output  [0:0] m_axi_mem_WID;
output  [0:0] m_axi_mem_WUSER;
output   m_axi_mem_ARVALID;
input   m_axi_mem_ARREADY;
output  [63:0] m_axi_mem_ARADDR;
output  [0:0] m_axi_mem_ARID;
output  [31:0] m_axi_mem_ARLEN;
output  [2:0] m_axi_mem_ARSIZE;
output  [1:0] m_axi_mem_ARBURST;
output  [1:0] m_axi_mem_ARLOCK;
output  [3:0] m_axi_mem_ARCACHE;
output  [2:0] m_axi_mem_ARPROT;
output  [3:0] m_axi_mem_ARQOS;
output  [3:0] m_axi_mem_ARREGION;
output  [0:0] m_axi_mem_ARUSER;
input   m_axi_mem_RVALID;
output   m_axi_mem_RREADY;
input  [63:0] m_axi_mem_RDATA;
input   m_axi_mem_RLAST;
input  [0:0] m_axi_mem_RID;
input  [8:0] m_axi_mem_RFIFONUM;
input  [0:0] m_axi_mem_RUSER;
input  [1:0] m_axi_mem_RRESP;
input   m_axi_mem_BVALID;
output   m_axi_mem_BREADY;
input  [1:0] m_axi_mem_BRESP;
input  [0:0] m_axi_mem_BID;
input  [0:0] m_axi_mem_BUSER;
input  [60:0] p_cast12_cast;
output  [7:0] centroid_y_coords_address0;
output   centroid_y_coords_ce0;
input  [63:0] centroid_y_coords_q0;
input  [31:0] sext_ln185;

reg ap_idle;
reg m_axi_mem_WVALID;
reg centroid_y_coords_ce0;

(* fsm_encoding = "none" *) reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_enable_reg_pp0_iter0;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter2;
reg    ap_enable_reg_pp0_iter3;
reg    ap_idle_pp0;
wire    ap_block_state1_pp0_stage0_iter0;
wire    ap_block_state2_pp0_stage0_iter1;
wire    ap_block_state3_pp0_stage0_iter2;
wire    ap_block_state4_pp0_stage0_iter3;
reg    ap_block_pp0_stage0_subdone;
wire   [0:0] exitcond_fu_118_p2;
reg    ap_condition_exit_pp0_iter1_stage0;
wire    ap_loop_exit_ready;
reg    ap_ready_int;
reg    mem_blk_n_W;
wire    ap_block_pp0_stage0;
wire  signed [60:0] sext_ln185_cast_fu_91_p1;
reg  signed [60:0] sext_ln185_cast_reg_141;
reg    ap_block_pp0_stage0_11001;
reg   [63:0] centroid_y_coords_load_reg_160;
wire   [63:0] loop_index_cast_fu_113_p1;
wire    ap_block_pp0_stage0_01001;
reg   [60:0] loop_index_fu_54;
wire   [60:0] empty_fu_107_p2;
wire    ap_loop_init;
reg    ap_done_reg;
wire    ap_continue_int;
reg    ap_done_int;
reg    ap_loop_exit_ready_pp0_iter2_reg;
reg    ap_loop_exit_ready_pp0_iter3_reg;
reg   [0:0] ap_NS_fsm;
wire    ap_enable_pp0;
wire    ap_start_int;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_CS_fsm = 1'd1;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_done_reg = 1'b0;
end

kmeans_top_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(ap_start),
    .ap_ready(ap_ready),
    .ap_done(ap_done),
    .ap_start_int(ap_start_int),
    .ap_loop_init(ap_loop_init),
    .ap_ready_int(ap_ready_int),
    .ap_loop_exit_ready(ap_condition_exit_pp0_iter1_stage0),
    .ap_loop_exit_done(ap_done_int),
    .ap_continue_int(ap_continue_int),
    .ap_done_int(ap_done_int)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue_int == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter3_reg == 1'b1))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b1 == ap_condition_exit_pp0_iter1_stage0)) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_enable_reg_pp0_iter1 <= ap_start_int;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter2_reg == 1'b0))) begin
        ap_loop_exit_ready_pp0_iter3_reg <= 1'b0;
    end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        ap_loop_exit_ready_pp0_iter3_reg <= ap_loop_exit_ready_pp0_iter2_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        if ((ap_loop_init == 1'b1)) begin
            loop_index_fu_54 <= 61'd0;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (exitcond_fu_118_p2 == 1'd0))) begin
            loop_index_fu_54 <= empty_fu_107_p2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_loop_exit_ready_pp0_iter2_reg <= ap_loop_exit_ready;
        sext_ln185_cast_reg_141 <= sext_ln185_cast_fu_91_p1;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        centroid_y_coords_load_reg_160 <= centroid_y_coords_q0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (exitcond_fu_118_p2 == 1'd1))) begin
        ap_condition_exit_pp0_iter1_stage0 = 1'b1;
    end else begin
        ap_condition_exit_pp0_iter1_stage0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter3_reg == 1'b1))) begin
        ap_done_int = 1'b1;
    end else begin
        ap_done_int = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_idle_pp0 == 1'b1) & (ap_start_int == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_ready_int = 1'b1;
    end else begin
        ap_ready_int = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        centroid_y_coords_ce0 = 1'b1;
    end else begin
        centroid_y_coords_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1))) begin
        m_axi_mem_WVALID = 1'b1;
    end else begin
        m_axi_mem_WVALID = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter3 == 1'b1))) begin
        mem_blk_n_W = m_axi_mem_WREADY;
    end else begin
        mem_blk_n_W = 1'b1;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_pp0_stage0 : begin
            ap_NS_fsm = ap_ST_fsm_pp0_stage0;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_01001 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_pp0_stage0_11001 = ((m_axi_mem_WREADY == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b1));
end

always @ (*) begin
    ap_block_pp0_stage0_subdone = ((m_axi_mem_WREADY == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b1));
end

assign ap_block_state1_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_enable_reg_pp0_iter0 = ap_start_int;

assign ap_loop_exit_ready = ap_condition_exit_pp0_iter1_stage0;

assign centroid_y_coords_address0 = loop_index_cast_fu_113_p1;

assign empty_fu_107_p2 = (loop_index_fu_54 + 61'd1);

assign exitcond_fu_118_p2 = ((empty_fu_107_p2 == sext_ln185_cast_reg_141) ? 1'b1 : 1'b0);

assign loop_index_cast_fu_113_p1 = loop_index_fu_54;

assign m_axi_mem_ARADDR = 64'd0;

assign m_axi_mem_ARBURST = 2'd0;

assign m_axi_mem_ARCACHE = 4'd0;

assign m_axi_mem_ARID = 1'd0;

assign m_axi_mem_ARLEN = 32'd0;

assign m_axi_mem_ARLOCK = 2'd0;

assign m_axi_mem_ARPROT = 3'd0;

assign m_axi_mem_ARQOS = 4'd0;

assign m_axi_mem_ARREGION = 4'd0;

assign m_axi_mem_ARSIZE = 3'd0;

assign m_axi_mem_ARUSER = 1'd0;

assign m_axi_mem_ARVALID = 1'b0;

assign m_axi_mem_AWADDR = 64'd0;

assign m_axi_mem_AWBURST = 2'd0;

assign m_axi_mem_AWCACHE = 4'd0;

assign m_axi_mem_AWID = 1'd0;

assign m_axi_mem_AWLEN = 32'd0;

assign m_axi_mem_AWLOCK = 2'd0;

assign m_axi_mem_AWPROT = 3'd0;

assign m_axi_mem_AWQOS = 4'd0;

assign m_axi_mem_AWREGION = 4'd0;

assign m_axi_mem_AWSIZE = 3'd0;

assign m_axi_mem_AWUSER = 1'd0;

assign m_axi_mem_AWVALID = 1'b0;

assign m_axi_mem_BREADY = 1'b0;

assign m_axi_mem_RREADY = 1'b0;

assign m_axi_mem_WDATA = centroid_y_coords_load_reg_160;

assign m_axi_mem_WID = 1'd0;

assign m_axi_mem_WLAST = 1'b0;

assign m_axi_mem_WSTRB = 8'd255;

assign m_axi_mem_WUSER = 1'd0;

assign sext_ln185_cast_fu_91_p1 = $signed(sext_ln185);

endmodule //kmeans_top_kmeans_top_Pipeline_13


// Content from kmeans_top_kmeans_top_Pipeline_5.v
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2022.2 (64-bit)
// Version: 2022.2
// Copyright (C) Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module kmeans_top_kmeans_top_Pipeline_5 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        m_axi_mem_AWVALID,
        m_axi_mem_AWREADY,
        m_axi_mem_AWADDR,
        m_axi_mem_AWID,
        m_axi_mem_AWLEN,
        m_axi_mem_AWSIZE,
        m_axi_mem_AWBURST,
        m_axi_mem_AWLOCK,
        m_axi_mem_AWCACHE,
        m_axi_mem_AWPROT,
        m_axi_mem_AWQOS,
        m_axi_mem_AWREGION,
        m_axi_mem_AWUSER,
        m_axi_mem_WVALID,
        m_axi_mem_WREADY,
        m_axi_mem_WDATA,
        m_axi_mem_WSTRB,
        m_axi_mem_WLAST,
        m_axi_mem_WID,
        m_axi_mem_WUSER,
        m_axi_mem_ARVALID,
        m_axi_mem_ARREADY,
        m_axi_mem_ARADDR,
        m_axi_mem_ARID,
        m_axi_mem_ARLEN,
        m_axi_mem_ARSIZE,
        m_axi_mem_ARBURST,
        m_axi_mem_ARLOCK,
        m_axi_mem_ARCACHE,
        m_axi_mem_ARPROT,
        m_axi_mem_ARQOS,
        m_axi_mem_ARREGION,
        m_axi_mem_ARUSER,
        m_axi_mem_RVALID,
        m_axi_mem_RREADY,
        m_axi_mem_RDATA,
        m_axi_mem_RLAST,
        m_axi_mem_RID,
        m_axi_mem_RFIFONUM,
        m_axi_mem_RUSER,
        m_axi_mem_RRESP,
        m_axi_mem_BVALID,
        m_axi_mem_BREADY,
        m_axi_mem_BRESP,
        m_axi_mem_BID,
        m_axi_mem_BUSER,
        p_cast3_cast,
        centroid_y_coords_address0,
        centroid_y_coords_ce0,
        centroid_y_coords_we0,
        centroid_y_coords_d0,
        sext_ln185
);

parameter    ap_ST_fsm_pp0_stage0 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
output   m_axi_mem_AWVALID;
input   m_axi_mem_AWREADY;
output  [63:0] m_axi_mem_AWADDR;
output  [0:0] m_axi_mem_AWID;
output  [31:0] m_axi_mem_AWLEN;
output  [2:0] m_axi_mem_AWSIZE;
output  [1:0] m_axi_mem_AWBURST;
output  [1:0] m_axi_mem_AWLOCK;
output  [3:0] m_axi_mem_AWCACHE;
output  [2:0] m_axi_mem_AWPROT;
output  [3:0] m_axi_mem_AWQOS;
output  [3:0] m_axi_mem_AWREGION;
output  [0:0] m_axi_mem_AWUSER;
output   m_axi_mem_WVALID;
input   m_axi_mem_WREADY;
output  [63:0] m_axi_mem_WDATA;
output  [7:0] m_axi_mem_WSTRB;
output   m_axi_mem_WLAST;
output  [0:0] m_axi_mem_WID;
output  [0:0] m_axi_mem_WUSER;
output   m_axi_mem_ARVALID;
input   m_axi_mem_ARREADY;
output  [63:0] m_axi_mem_ARADDR;
output  [0:0] m_axi_mem_ARID;
output  [31:0] m_axi_mem_ARLEN;
output  [2:0] m_axi_mem_ARSIZE;
output  [1:0] m_axi_mem_ARBURST;
output  [1:0] m_axi_mem_ARLOCK;
output  [3:0] m_axi_mem_ARCACHE;
output  [2:0] m_axi_mem_ARPROT;
output  [3:0] m_axi_mem_ARQOS;
output  [3:0] m_axi_mem_ARREGION;
output  [0:0] m_axi_mem_ARUSER;
input   m_axi_mem_RVALID;
output   m_axi_mem_RREADY;
input  [63:0] m_axi_mem_RDATA;
input   m_axi_mem_RLAST;
input  [0:0] m_axi_mem_RID;
input  [8:0] m_axi_mem_RFIFONUM;
input  [0:0] m_axi_mem_RUSER;
input  [1:0] m_axi_mem_RRESP;
input   m_axi_mem_BVALID;
output   m_axi_mem_BREADY;
input  [1:0] m_axi_mem_BRESP;
input  [0:0] m_axi_mem_BID;
input  [0:0] m_axi_mem_BUSER;
input  [60:0] p_cast3_cast;
output  [7:0] centroid_y_coords_address0;
output   centroid_y_coords_ce0;
output   centroid_y_coords_we0;
output  [63:0] centroid_y_coords_d0;
input  [31:0] sext_ln185;

reg ap_idle;
reg m_axi_mem_RREADY;
reg centroid_y_coords_ce0;
reg centroid_y_coords_we0;

(* fsm_encoding = "none" *) reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_enable_reg_pp0_iter0;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter2;
reg    ap_idle_pp0;
wire    ap_block_state1_pp0_stage0_iter0;
reg    ap_block_state2_pp0_stage0_iter1;
wire    ap_block_state3_pp0_stage0_iter2;
reg    ap_block_pp0_stage0_subdone;
wire   [0:0] exitcond81_fu_114_p2;
reg    ap_condition_exit_pp0_iter1_stage0;
wire    ap_loop_exit_ready;
reg    ap_ready_int;
reg    mem_blk_n_R;
wire    ap_block_pp0_stage0;
wire  signed [60:0] sext_ln185_cast_fu_86_p1;
reg  signed [60:0] sext_ln185_cast_reg_135;
reg    ap_block_pp0_stage0_11001;
reg   [60:0] loop_index45_load_reg_145;
reg   [63:0] mem_addr_read_reg_150;
wire   [63:0] loop_index45_cast_fu_124_p1;
reg   [60:0] loop_index45_fu_52;
wire   [60:0] empty_fu_102_p2;
wire    ap_loop_init;
reg    ap_done_reg;
wire    ap_continue_int;
reg    ap_done_int;
reg    ap_loop_exit_ready_pp0_iter2_reg;
reg   [0:0] ap_NS_fsm;
wire    ap_enable_pp0;
wire    ap_start_int;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_CS_fsm = 1'd1;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_done_reg = 1'b0;
end

kmeans_top_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(ap_start),
    .ap_ready(ap_ready),
    .ap_done(ap_done),
    .ap_start_int(ap_start_int),
    .ap_loop_init(ap_loop_init),
    .ap_ready_int(ap_ready_int),
    .ap_loop_exit_ready(ap_condition_exit_pp0_iter1_stage0),
    .ap_loop_exit_done(ap_done_int),
    .ap_continue_int(ap_continue_int),
    .ap_done_int(ap_done_int)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue_int == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter2_reg == 1'b1))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b1 == ap_condition_exit_pp0_iter1_stage0)) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_enable_reg_pp0_iter1 <= ap_start_int;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready == 1'b0))) begin
        ap_loop_exit_ready_pp0_iter2_reg <= 1'b0;
    end else if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_loop_exit_ready_pp0_iter2_reg <= ap_loop_exit_ready;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        if ((ap_loop_init == 1'b1)) begin
            loop_index45_fu_52 <= 61'd0;
        end else if (((exitcond81_fu_114_p2 == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
            loop_index45_fu_52 <= empty_fu_102_p2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        loop_index45_load_reg_145 <= loop_index45_fu_52;
        mem_addr_read_reg_150 <= m_axi_mem_RDATA;
        sext_ln185_cast_reg_135 <= sext_ln185_cast_fu_86_p1;
    end
end

always @ (*) begin
    if (((exitcond81_fu_114_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_condition_exit_pp0_iter1_stage0 = 1'b1;
    end else begin
        ap_condition_exit_pp0_iter1_stage0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter2_reg == 1'b1))) begin
        ap_done_int = 1'b1;
    end else begin
        ap_done_int = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_idle_pp0 == 1'b1) & (ap_start_int == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_ready_int = 1'b1;
    end else begin
        ap_ready_int = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        centroid_y_coords_ce0 = 1'b1;
    end else begin
        centroid_y_coords_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        centroid_y_coords_we0 = 1'b1;
    end else begin
        centroid_y_coords_we0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        m_axi_mem_RREADY = 1'b1;
    end else begin
        m_axi_mem_RREADY = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        mem_blk_n_R = m_axi_mem_RVALID;
    end else begin
        mem_blk_n_R = 1'b1;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_pp0_stage0 : begin
            ap_NS_fsm = ap_ST_fsm_pp0_stage0;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_pp0_stage0_11001 = ((m_axi_mem_RVALID == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b1));
end

always @ (*) begin
    ap_block_pp0_stage0_subdone = ((m_axi_mem_RVALID == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b1));
end

assign ap_block_state1_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state2_pp0_stage0_iter1 = (m_axi_mem_RVALID == 1'b0);
end

assign ap_block_state3_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_enable_reg_pp0_iter0 = ap_start_int;

assign ap_loop_exit_ready = ap_condition_exit_pp0_iter1_stage0;

assign centroid_y_coords_address0 = loop_index45_cast_fu_124_p1;

assign centroid_y_coords_d0 = mem_addr_read_reg_150;

assign empty_fu_102_p2 = (loop_index45_fu_52 + 61'd1);

assign exitcond81_fu_114_p2 = ((empty_fu_102_p2 == sext_ln185_cast_reg_135) ? 1'b1 : 1'b0);

assign loop_index45_cast_fu_124_p1 = loop_index45_load_reg_145;

assign m_axi_mem_ARADDR = 64'd0;

assign m_axi_mem_ARBURST = 2'd0;

assign m_axi_mem_ARCACHE = 4'd0;

assign m_axi_mem_ARID = 1'd0;

assign m_axi_mem_ARLEN = 32'd0;

assign m_axi_mem_ARLOCK = 2'd0;

assign m_axi_mem_ARPROT = 3'd0;

assign m_axi_mem_ARQOS = 4'd0;

assign m_axi_mem_ARREGION = 4'd0;

assign m_axi_mem_ARSIZE = 3'd0;

assign m_axi_mem_ARUSER = 1'd0;

assign m_axi_mem_ARVALID = 1'b0;

assign m_axi_mem_AWADDR = 64'd0;

assign m_axi_mem_AWBURST = 2'd0;

assign m_axi_mem_AWCACHE = 4'd0;

assign m_axi_mem_AWID = 1'd0;

assign m_axi_mem_AWLEN = 32'd0;

assign m_axi_mem_AWLOCK = 2'd0;

assign m_axi_mem_AWPROT = 3'd0;

assign m_axi_mem_AWQOS = 4'd0;

assign m_axi_mem_AWREGION = 4'd0;

assign m_axi_mem_AWSIZE = 3'd0;

assign m_axi_mem_AWUSER = 1'd0;

assign m_axi_mem_AWVALID = 1'b0;

assign m_axi_mem_BREADY = 1'b0;

assign m_axi_mem_WDATA = 64'd0;

assign m_axi_mem_WID = 1'd0;

assign m_axi_mem_WLAST = 1'b0;

assign m_axi_mem_WSTRB = 8'd0;

assign m_axi_mem_WUSER = 1'd0;

assign m_axi_mem_WVALID = 1'b0;

assign sext_ln185_cast_fu_86_p1 = $signed(sext_ln185);

endmodule //kmeans_top_kmeans_top_Pipeline_5


// Content from kmeans_top_kmeans_top_Pipeline_9.v
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2022.2 (64-bit)
// Version: 2022.2
// Copyright (C) Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module kmeans_top_kmeans_top_Pipeline_9 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        m_axi_mem_AWVALID,
        m_axi_mem_AWREADY,
        m_axi_mem_AWADDR,
        m_axi_mem_AWID,
        m_axi_mem_AWLEN,
        m_axi_mem_AWSIZE,
        m_axi_mem_AWBURST,
        m_axi_mem_AWLOCK,
        m_axi_mem_AWCACHE,
        m_axi_mem_AWPROT,
        m_axi_mem_AWQOS,
        m_axi_mem_AWREGION,
        m_axi_mem_AWUSER,
        m_axi_mem_WVALID,
        m_axi_mem_WREADY,
        m_axi_mem_WDATA,
        m_axi_mem_WSTRB,
        m_axi_mem_WLAST,
        m_axi_mem_WID,
        m_axi_mem_WUSER,
        m_axi_mem_ARVALID,
        m_axi_mem_ARREADY,
        m_axi_mem_ARADDR,
        m_axi_mem_ARID,
        m_axi_mem_ARLEN,
        m_axi_mem_ARSIZE,
        m_axi_mem_ARBURST,
        m_axi_mem_ARLOCK,
        m_axi_mem_ARCACHE,
        m_axi_mem_ARPROT,
        m_axi_mem_ARQOS,
        m_axi_mem_ARREGION,
        m_axi_mem_ARUSER,
        m_axi_mem_RVALID,
        m_axi_mem_RREADY,
        m_axi_mem_RDATA,
        m_axi_mem_RLAST,
        m_axi_mem_RID,
        m_axi_mem_RFIFONUM,
        m_axi_mem_RUSER,
        m_axi_mem_RRESP,
        m_axi_mem_BVALID,
        m_axi_mem_BREADY,
        m_axi_mem_BRESP,
        m_axi_mem_BID,
        m_axi_mem_BUSER,
        p_cast5_cast,
        node_x_coords_address0,
        node_x_coords_ce0,
        node_x_coords_q0,
        sext_ln182
);

parameter    ap_ST_fsm_pp0_stage0 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
output   m_axi_mem_AWVALID;
input   m_axi_mem_AWREADY;
output  [63:0] m_axi_mem_AWADDR;
output  [0:0] m_axi_mem_AWID;
output  [31:0] m_axi_mem_AWLEN;
output  [2:0] m_axi_mem_AWSIZE;
output  [1:0] m_axi_mem_AWBURST;
output  [1:0] m_axi_mem_AWLOCK;
output  [3:0] m_axi_mem_AWCACHE;
output  [2:0] m_axi_mem_AWPROT;
output  [3:0] m_axi_mem_AWQOS;
output  [3:0] m_axi_mem_AWREGION;
output  [0:0] m_axi_mem_AWUSER;
output   m_axi_mem_WVALID;
input   m_axi_mem_WREADY;
output  [63:0] m_axi_mem_WDATA;
output  [7:0] m_axi_mem_WSTRB;
output   m_axi_mem_WLAST;
output  [0:0] m_axi_mem_WID;
output  [0:0] m_axi_mem_WUSER;
output   m_axi_mem_ARVALID;
input   m_axi_mem_ARREADY;
output  [63:0] m_axi_mem_ARADDR;
output  [0:0] m_axi_mem_ARID;
output  [31:0] m_axi_mem_ARLEN;
output  [2:0] m_axi_mem_ARSIZE;
output  [1:0] m_axi_mem_ARBURST;
output  [1:0] m_axi_mem_ARLOCK;
output  [3:0] m_axi_mem_ARCACHE;
output  [2:0] m_axi_mem_ARPROT;
output  [3:0] m_axi_mem_ARQOS;
output  [3:0] m_axi_mem_ARREGION;
output  [0:0] m_axi_mem_ARUSER;
input   m_axi_mem_RVALID;
output   m_axi_mem_RREADY;
input  [63:0] m_axi_mem_RDATA;
input   m_axi_mem_RLAST;
input  [0:0] m_axi_mem_RID;
input  [8:0] m_axi_mem_RFIFONUM;
input  [0:0] m_axi_mem_RUSER;
input  [1:0] m_axi_mem_RRESP;
input   m_axi_mem_BVALID;
output   m_axi_mem_BREADY;
input  [1:0] m_axi_mem_BRESP;
input  [0:0] m_axi_mem_BID;
input  [0:0] m_axi_mem_BUSER;
input  [60:0] p_cast5_cast;
output  [12:0] node_x_coords_address0;
output   node_x_coords_ce0;
input  [63:0] node_x_coords_q0;
input  [31:0] sext_ln182;

reg ap_idle;
reg m_axi_mem_WVALID;
reg node_x_coords_ce0;

(* fsm_encoding = "none" *) reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_enable_reg_pp0_iter0;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter2;
reg    ap_enable_reg_pp0_iter3;
reg    ap_idle_pp0;
wire    ap_block_state1_pp0_stage0_iter0;
wire    ap_block_state2_pp0_stage0_iter1;
wire    ap_block_state3_pp0_stage0_iter2;
wire    ap_block_state4_pp0_stage0_iter3;
reg    ap_block_pp0_stage0_subdone;
wire   [0:0] exitcond77_fu_126_p2;
reg    ap_condition_exit_pp0_iter1_stage0;
wire    ap_loop_exit_ready;
reg    ap_ready_int;
reg    mem_blk_n_W;
wire    ap_block_pp0_stage0;
wire  signed [60:0] sext_ln182_cast_fu_99_p1;
reg  signed [60:0] sext_ln182_cast_reg_149;
reg    ap_block_pp0_stage0_11001;
reg   [63:0] node_x_coords_load_reg_168;
wire   [63:0] loop_index21_cast_fu_121_p1;
wire    ap_block_pp0_stage0_01001;
reg   [60:0] loop_index21_fu_62;
wire   [60:0] empty_fu_115_p2;
wire    ap_loop_init;
reg    ap_done_reg;
wire    ap_continue_int;
reg    ap_done_int;
reg    ap_loop_exit_ready_pp0_iter2_reg;
reg    ap_loop_exit_ready_pp0_iter3_reg;
reg   [0:0] ap_NS_fsm;
wire    ap_enable_pp0;
wire    ap_start_int;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_CS_fsm = 1'd1;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_done_reg = 1'b0;
end

kmeans_top_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(ap_start),
    .ap_ready(ap_ready),
    .ap_done(ap_done),
    .ap_start_int(ap_start_int),
    .ap_loop_init(ap_loop_init),
    .ap_ready_int(ap_ready_int),
    .ap_loop_exit_ready(ap_condition_exit_pp0_iter1_stage0),
    .ap_loop_exit_done(ap_done_int),
    .ap_continue_int(ap_continue_int),
    .ap_done_int(ap_done_int)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue_int == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter3_reg == 1'b1))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b1 == ap_condition_exit_pp0_iter1_stage0)) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_enable_reg_pp0_iter1 <= ap_start_int;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter2_reg == 1'b0))) begin
        ap_loop_exit_ready_pp0_iter3_reg <= 1'b0;
    end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        ap_loop_exit_ready_pp0_iter3_reg <= ap_loop_exit_ready_pp0_iter2_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        if ((ap_loop_init == 1'b1)) begin
            loop_index21_fu_62 <= 61'd0;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (exitcond77_fu_126_p2 == 1'd0))) begin
            loop_index21_fu_62 <= empty_fu_115_p2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_loop_exit_ready_pp0_iter2_reg <= ap_loop_exit_ready;
        sext_ln182_cast_reg_149 <= sext_ln182_cast_fu_99_p1;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        node_x_coords_load_reg_168 <= node_x_coords_q0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (exitcond77_fu_126_p2 == 1'd1))) begin
        ap_condition_exit_pp0_iter1_stage0 = 1'b1;
    end else begin
        ap_condition_exit_pp0_iter1_stage0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter3_reg == 1'b1))) begin
        ap_done_int = 1'b1;
    end else begin
        ap_done_int = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_idle_pp0 == 1'b1) & (ap_start_int == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_ready_int = 1'b1;
    end else begin
        ap_ready_int = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1))) begin
        m_axi_mem_WVALID = 1'b1;
    end else begin
        m_axi_mem_WVALID = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter3 == 1'b1))) begin
        mem_blk_n_W = m_axi_mem_WREADY;
    end else begin
        mem_blk_n_W = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        node_x_coords_ce0 = 1'b1;
    end else begin
        node_x_coords_ce0 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_pp0_stage0 : begin
            ap_NS_fsm = ap_ST_fsm_pp0_stage0;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_01001 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_pp0_stage0_11001 = ((m_axi_mem_WREADY == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b1));
end

always @ (*) begin
    ap_block_pp0_stage0_subdone = ((m_axi_mem_WREADY == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b1));
end

assign ap_block_state1_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_enable_reg_pp0_iter0 = ap_start_int;

assign ap_loop_exit_ready = ap_condition_exit_pp0_iter1_stage0;

assign empty_fu_115_p2 = (loop_index21_fu_62 + 61'd1);

assign exitcond77_fu_126_p2 = ((empty_fu_115_p2 == sext_ln182_cast_reg_149) ? 1'b1 : 1'b0);

assign loop_index21_cast_fu_121_p1 = loop_index21_fu_62;

assign m_axi_mem_ARADDR = 64'd0;

assign m_axi_mem_ARBURST = 2'd0;

assign m_axi_mem_ARCACHE = 4'd0;

assign m_axi_mem_ARID = 1'd0;

assign m_axi_mem_ARLEN = 32'd0;

assign m_axi_mem_ARLOCK = 2'd0;

assign m_axi_mem_ARPROT = 3'd0;

assign m_axi_mem_ARQOS = 4'd0;

assign m_axi_mem_ARREGION = 4'd0;

assign m_axi_mem_ARSIZE = 3'd0;

assign m_axi_mem_ARUSER = 1'd0;

assign m_axi_mem_ARVALID = 1'b0;

assign m_axi_mem_AWADDR = 64'd0;

assign m_axi_mem_AWBURST = 2'd0;

assign m_axi_mem_AWCACHE = 4'd0;

assign m_axi_mem_AWID = 1'd0;

assign m_axi_mem_AWLEN = 32'd0;

assign m_axi_mem_AWLOCK = 2'd0;

assign m_axi_mem_AWPROT = 3'd0;

assign m_axi_mem_AWQOS = 4'd0;

assign m_axi_mem_AWREGION = 4'd0;

assign m_axi_mem_AWSIZE = 3'd0;

assign m_axi_mem_AWUSER = 1'd0;

assign m_axi_mem_AWVALID = 1'b0;

assign m_axi_mem_BREADY = 1'b0;

assign m_axi_mem_RREADY = 1'b0;

assign m_axi_mem_WDATA = node_x_coords_load_reg_168;

assign m_axi_mem_WID = 1'd0;

assign m_axi_mem_WLAST = 1'b0;

assign m_axi_mem_WSTRB = 8'd255;

assign m_axi_mem_WUSER = 1'd0;

assign node_x_coords_address0 = loop_index21_cast_fu_121_p1;

assign sext_ln182_cast_fu_99_p1 = $signed(sext_ln182);

endmodule //kmeans_top_kmeans_top_Pipeline_9


// Content from kmeans_top_kmeans_top_Pipeline_7.v
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2022.2 (64-bit)
// Version: 2022.2
// Copyright (C) Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module kmeans_top_kmeans_top_Pipeline_7 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        m_axi_mem_AWVALID,
        m_axi_mem_AWREADY,
        m_axi_mem_AWADDR,
        m_axi_mem_AWID,
        m_axi_mem_AWLEN,
        m_axi_mem_AWSIZE,
        m_axi_mem_AWBURST,
        m_axi_mem_AWLOCK,
        m_axi_mem_AWCACHE,
        m_axi_mem_AWPROT,
        m_axi_mem_AWQOS,
        m_axi_mem_AWREGION,
        m_axi_mem_AWUSER,
        m_axi_mem_WVALID,
        m_axi_mem_WREADY,
        m_axi_mem_WDATA,
        m_axi_mem_WSTRB,
        m_axi_mem_WLAST,
        m_axi_mem_WID,
        m_axi_mem_WUSER,
        m_axi_mem_ARVALID,
        m_axi_mem_ARREADY,
        m_axi_mem_ARADDR,
        m_axi_mem_ARID,
        m_axi_mem_ARLEN,
        m_axi_mem_ARSIZE,
        m_axi_mem_ARBURST,
        m_axi_mem_ARLOCK,
        m_axi_mem_ARCACHE,
        m_axi_mem_ARPROT,
        m_axi_mem_ARQOS,
        m_axi_mem_ARREGION,
        m_axi_mem_ARUSER,
        m_axi_mem_RVALID,
        m_axi_mem_RREADY,
        m_axi_mem_RDATA,
        m_axi_mem_RLAST,
        m_axi_mem_RID,
        m_axi_mem_RFIFONUM,
        m_axi_mem_RUSER,
        m_axi_mem_RRESP,
        m_axi_mem_BVALID,
        m_axi_mem_BREADY,
        m_axi_mem_BRESP,
        m_axi_mem_BID,
        m_axi_mem_BUSER,
        p_cast11_cast,
        centroid_x_coords_address0,
        centroid_x_coords_ce0,
        centroid_x_coords_q0,
        sext_ln185
);

parameter    ap_ST_fsm_pp0_stage0 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
output   m_axi_mem_AWVALID;
input   m_axi_mem_AWREADY;
output  [63:0] m_axi_mem_AWADDR;
output  [0:0] m_axi_mem_AWID;
output  [31:0] m_axi_mem_AWLEN;
output  [2:0] m_axi_mem_AWSIZE;
output  [1:0] m_axi_mem_AWBURST;
output  [1:0] m_axi_mem_AWLOCK;
output  [3:0] m_axi_mem_AWCACHE;
output  [2:0] m_axi_mem_AWPROT;
output  [3:0] m_axi_mem_AWQOS;
output  [3:0] m_axi_mem_AWREGION;
output  [0:0] m_axi_mem_AWUSER;
output   m_axi_mem_WVALID;
input   m_axi_mem_WREADY;
output  [63:0] m_axi_mem_WDATA;
output  [7:0] m_axi_mem_WSTRB;
output   m_axi_mem_WLAST;
output  [0:0] m_axi_mem_WID;
output  [0:0] m_axi_mem_WUSER;
output   m_axi_mem_ARVALID;
input   m_axi_mem_ARREADY;
output  [63:0] m_axi_mem_ARADDR;
output  [0:0] m_axi_mem_ARID;
output  [31:0] m_axi_mem_ARLEN;
output  [2:0] m_axi_mem_ARSIZE;
output  [1:0] m_axi_mem_ARBURST;
output  [1:0] m_axi_mem_ARLOCK;
output  [3:0] m_axi_mem_ARCACHE;
output  [2:0] m_axi_mem_ARPROT;
output  [3:0] m_axi_mem_ARQOS;
output  [3:0] m_axi_mem_ARREGION;
output  [0:0] m_axi_mem_ARUSER;
input   m_axi_mem_RVALID;
output   m_axi_mem_RREADY;
input  [63:0] m_axi_mem_RDATA;
input   m_axi_mem_RLAST;
input  [0:0] m_axi_mem_RID;
input  [8:0] m_axi_mem_RFIFONUM;
input  [0:0] m_axi_mem_RUSER;
input  [1:0] m_axi_mem_RRESP;
input   m_axi_mem_BVALID;
output   m_axi_mem_BREADY;
input  [1:0] m_axi_mem_BRESP;
input  [0:0] m_axi_mem_BID;
input  [0:0] m_axi_mem_BUSER;
input  [60:0] p_cast11_cast;
output  [7:0] centroid_x_coords_address0;
output   centroid_x_coords_ce0;
input  [63:0] centroid_x_coords_q0;
input  [31:0] sext_ln185;

reg ap_idle;
reg m_axi_mem_WVALID;
reg centroid_x_coords_ce0;

(* fsm_encoding = "none" *) reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_enable_reg_pp0_iter0;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter2;
reg    ap_enable_reg_pp0_iter3;
reg    ap_idle_pp0;
wire    ap_block_state1_pp0_stage0_iter0;
wire    ap_block_state2_pp0_stage0_iter1;
wire    ap_block_state3_pp0_stage0_iter2;
wire    ap_block_state4_pp0_stage0_iter3;
reg    ap_block_pp0_stage0_subdone;
wire   [0:0] exitcond79_fu_118_p2;
reg    ap_condition_exit_pp0_iter1_stage0;
wire    ap_loop_exit_ready;
reg    ap_ready_int;
reg    mem_blk_n_W;
wire    ap_block_pp0_stage0;
wire  signed [60:0] sext_ln185_cast_fu_91_p1;
reg  signed [60:0] sext_ln185_cast_reg_141;
reg    ap_block_pp0_stage0_11001;
reg   [63:0] centroid_x_coords_load_reg_160;
wire   [63:0] loop_index33_cast_fu_113_p1;
wire    ap_block_pp0_stage0_01001;
reg   [60:0] loop_index33_fu_54;
wire   [60:0] empty_fu_107_p2;
wire    ap_loop_init;
reg    ap_done_reg;
wire    ap_continue_int;
reg    ap_done_int;
reg    ap_loop_exit_ready_pp0_iter2_reg;
reg    ap_loop_exit_ready_pp0_iter3_reg;
reg   [0:0] ap_NS_fsm;
wire    ap_enable_pp0;
wire    ap_start_int;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_CS_fsm = 1'd1;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_done_reg = 1'b0;
end

kmeans_top_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(ap_start),
    .ap_ready(ap_ready),
    .ap_done(ap_done),
    .ap_start_int(ap_start_int),
    .ap_loop_init(ap_loop_init),
    .ap_ready_int(ap_ready_int),
    .ap_loop_exit_ready(ap_condition_exit_pp0_iter1_stage0),
    .ap_loop_exit_done(ap_done_int),
    .ap_continue_int(ap_continue_int),
    .ap_done_int(ap_done_int)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue_int == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter3_reg == 1'b1))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b1 == ap_condition_exit_pp0_iter1_stage0)) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_enable_reg_pp0_iter1 <= ap_start_int;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter2_reg == 1'b0))) begin
        ap_loop_exit_ready_pp0_iter3_reg <= 1'b0;
    end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        ap_loop_exit_ready_pp0_iter3_reg <= ap_loop_exit_ready_pp0_iter2_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        if ((ap_loop_init == 1'b1)) begin
            loop_index33_fu_54 <= 61'd0;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (exitcond79_fu_118_p2 == 1'd0))) begin
            loop_index33_fu_54 <= empty_fu_107_p2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_loop_exit_ready_pp0_iter2_reg <= ap_loop_exit_ready;
        sext_ln185_cast_reg_141 <= sext_ln185_cast_fu_91_p1;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        centroid_x_coords_load_reg_160 <= centroid_x_coords_q0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (exitcond79_fu_118_p2 == 1'd1))) begin
        ap_condition_exit_pp0_iter1_stage0 = 1'b1;
    end else begin
        ap_condition_exit_pp0_iter1_stage0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter3_reg == 1'b1))) begin
        ap_done_int = 1'b1;
    end else begin
        ap_done_int = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_idle_pp0 == 1'b1) & (ap_start_int == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_ready_int = 1'b1;
    end else begin
        ap_ready_int = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        centroid_x_coords_ce0 = 1'b1;
    end else begin
        centroid_x_coords_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1))) begin
        m_axi_mem_WVALID = 1'b1;
    end else begin
        m_axi_mem_WVALID = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter3 == 1'b1))) begin
        mem_blk_n_W = m_axi_mem_WREADY;
    end else begin
        mem_blk_n_W = 1'b1;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_pp0_stage0 : begin
            ap_NS_fsm = ap_ST_fsm_pp0_stage0;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_01001 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_pp0_stage0_11001 = ((m_axi_mem_WREADY == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b1));
end

always @ (*) begin
    ap_block_pp0_stage0_subdone = ((m_axi_mem_WREADY == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b1));
end

assign ap_block_state1_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_enable_reg_pp0_iter0 = ap_start_int;

assign ap_loop_exit_ready = ap_condition_exit_pp0_iter1_stage0;

assign centroid_x_coords_address0 = loop_index33_cast_fu_113_p1;

assign empty_fu_107_p2 = (loop_index33_fu_54 + 61'd1);

assign exitcond79_fu_118_p2 = ((empty_fu_107_p2 == sext_ln185_cast_reg_141) ? 1'b1 : 1'b0);

assign loop_index33_cast_fu_113_p1 = loop_index33_fu_54;

assign m_axi_mem_ARADDR = 64'd0;

assign m_axi_mem_ARBURST = 2'd0;

assign m_axi_mem_ARCACHE = 4'd0;

assign m_axi_mem_ARID = 1'd0;

assign m_axi_mem_ARLEN = 32'd0;

assign m_axi_mem_ARLOCK = 2'd0;

assign m_axi_mem_ARPROT = 3'd0;

assign m_axi_mem_ARQOS = 4'd0;

assign m_axi_mem_ARREGION = 4'd0;

assign m_axi_mem_ARSIZE = 3'd0;

assign m_axi_mem_ARUSER = 1'd0;

assign m_axi_mem_ARVALID = 1'b0;

assign m_axi_mem_AWADDR = 64'd0;

assign m_axi_mem_AWBURST = 2'd0;

assign m_axi_mem_AWCACHE = 4'd0;

assign m_axi_mem_AWID = 1'd0;

assign m_axi_mem_AWLEN = 32'd0;

assign m_axi_mem_AWLOCK = 2'd0;

assign m_axi_mem_AWPROT = 3'd0;

assign m_axi_mem_AWQOS = 4'd0;

assign m_axi_mem_AWREGION = 4'd0;

assign m_axi_mem_AWSIZE = 3'd0;

assign m_axi_mem_AWUSER = 1'd0;

assign m_axi_mem_AWVALID = 1'b0;

assign m_axi_mem_BREADY = 1'b0;

assign m_axi_mem_RREADY = 1'b0;

assign m_axi_mem_WDATA = centroid_x_coords_load_reg_160;

assign m_axi_mem_WID = 1'd0;

assign m_axi_mem_WLAST = 1'b0;

assign m_axi_mem_WSTRB = 8'd255;

assign m_axi_mem_WUSER = 1'd0;

assign sext_ln185_cast_fu_91_p1 = $signed(sext_ln185);

endmodule //kmeans_top_kmeans_top_Pipeline_7


// Content from kmeans_top_kmeans_top_Pipeline_3.v
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2022.2 (64-bit)
// Version: 2022.2
// Copyright (C) Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module kmeans_top_kmeans_top_Pipeline_3 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        m_axi_mem_AWVALID,
        m_axi_mem_AWREADY,
        m_axi_mem_AWADDR,
        m_axi_mem_AWID,
        m_axi_mem_AWLEN,
        m_axi_mem_AWSIZE,
        m_axi_mem_AWBURST,
        m_axi_mem_AWLOCK,
        m_axi_mem_AWCACHE,
        m_axi_mem_AWPROT,
        m_axi_mem_AWQOS,
        m_axi_mem_AWREGION,
        m_axi_mem_AWUSER,
        m_axi_mem_WVALID,
        m_axi_mem_WREADY,
        m_axi_mem_WDATA,
        m_axi_mem_WSTRB,
        m_axi_mem_WLAST,
        m_axi_mem_WID,
        m_axi_mem_WUSER,
        m_axi_mem_ARVALID,
        m_axi_mem_ARREADY,
        m_axi_mem_ARADDR,
        m_axi_mem_ARID,
        m_axi_mem_ARLEN,
        m_axi_mem_ARSIZE,
        m_axi_mem_ARBURST,
        m_axi_mem_ARLOCK,
        m_axi_mem_ARCACHE,
        m_axi_mem_ARPROT,
        m_axi_mem_ARQOS,
        m_axi_mem_ARREGION,
        m_axi_mem_ARUSER,
        m_axi_mem_RVALID,
        m_axi_mem_RREADY,
        m_axi_mem_RDATA,
        m_axi_mem_RLAST,
        m_axi_mem_RID,
        m_axi_mem_RFIFONUM,
        m_axi_mem_RUSER,
        m_axi_mem_RRESP,
        m_axi_mem_BVALID,
        m_axi_mem_BREADY,
        m_axi_mem_BRESP,
        m_axi_mem_BID,
        m_axi_mem_BUSER,
        p_cast4_cast,
        node_cluster_assignments_address1,
        node_cluster_assignments_ce1,
        node_cluster_assignments_we1,
        node_cluster_assignments_d1,
        sext_ln182
);

parameter    ap_ST_fsm_pp0_stage0 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
output   m_axi_mem_AWVALID;
input   m_axi_mem_AWREADY;
output  [63:0] m_axi_mem_AWADDR;
output  [0:0] m_axi_mem_AWID;
output  [31:0] m_axi_mem_AWLEN;
output  [2:0] m_axi_mem_AWSIZE;
output  [1:0] m_axi_mem_AWBURST;
output  [1:0] m_axi_mem_AWLOCK;
output  [3:0] m_axi_mem_AWCACHE;
output  [2:0] m_axi_mem_AWPROT;
output  [3:0] m_axi_mem_AWQOS;
output  [3:0] m_axi_mem_AWREGION;
output  [0:0] m_axi_mem_AWUSER;
output   m_axi_mem_WVALID;
input   m_axi_mem_WREADY;
output  [63:0] m_axi_mem_WDATA;
output  [7:0] m_axi_mem_WSTRB;
output   m_axi_mem_WLAST;
output  [0:0] m_axi_mem_WID;
output  [0:0] m_axi_mem_WUSER;
output   m_axi_mem_ARVALID;
input   m_axi_mem_ARREADY;
output  [63:0] m_axi_mem_ARADDR;
output  [0:0] m_axi_mem_ARID;
output  [31:0] m_axi_mem_ARLEN;
output  [2:0] m_axi_mem_ARSIZE;
output  [1:0] m_axi_mem_ARBURST;
output  [1:0] m_axi_mem_ARLOCK;
output  [3:0] m_axi_mem_ARCACHE;
output  [2:0] m_axi_mem_ARPROT;
output  [3:0] m_axi_mem_ARQOS;
output  [3:0] m_axi_mem_ARREGION;
output  [0:0] m_axi_mem_ARUSER;
input   m_axi_mem_RVALID;
output   m_axi_mem_RREADY;
input  [63:0] m_axi_mem_RDATA;
input   m_axi_mem_RLAST;
input  [0:0] m_axi_mem_RID;
input  [8:0] m_axi_mem_RFIFONUM;
input  [0:0] m_axi_mem_RUSER;
input  [1:0] m_axi_mem_RRESP;
input   m_axi_mem_BVALID;
output   m_axi_mem_BREADY;
input  [1:0] m_axi_mem_BRESP;
input  [0:0] m_axi_mem_BID;
input  [0:0] m_axi_mem_BUSER;
input  [60:0] p_cast4_cast;
output  [12:0] node_cluster_assignments_address1;
output   node_cluster_assignments_ce1;
output   node_cluster_assignments_we1;
output  [63:0] node_cluster_assignments_d1;
input  [31:0] sext_ln182;

reg ap_idle;
reg m_axi_mem_RREADY;
reg node_cluster_assignments_ce1;
reg node_cluster_assignments_we1;

(* fsm_encoding = "none" *) reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_enable_reg_pp0_iter0;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter2;
reg    ap_idle_pp0;
wire    ap_block_state1_pp0_stage0_iter0;
reg    ap_block_state2_pp0_stage0_iter1;
wire    ap_block_state3_pp0_stage0_iter2;
reg    ap_block_pp0_stage0_subdone;
wire   [0:0] exitcond83_fu_126_p2;
reg    ap_condition_exit_pp0_iter1_stage0;
wire    ap_loop_exit_ready;
reg    ap_ready_int;
reg    mem_blk_n_R;
wire    ap_block_pp0_stage0;
wire  signed [60:0] sext_ln182_cast_fu_98_p1;
reg  signed [60:0] sext_ln182_cast_reg_147;
reg    ap_block_pp0_stage0_11001;
reg   [60:0] loop_index57_load_reg_157;
reg   [63:0] mem_addr_read_reg_162;
wire   [63:0] loop_index57_cast_fu_136_p1;
reg   [60:0] loop_index57_fu_60;
wire   [60:0] empty_fu_114_p2;
wire    ap_loop_init;
reg    ap_done_reg;
wire    ap_continue_int;
reg    ap_done_int;
reg    ap_loop_exit_ready_pp0_iter2_reg;
reg   [0:0] ap_NS_fsm;
wire    ap_enable_pp0;
wire    ap_start_int;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_CS_fsm = 1'd1;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_done_reg = 1'b0;
end

kmeans_top_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(ap_start),
    .ap_ready(ap_ready),
    .ap_done(ap_done),
    .ap_start_int(ap_start_int),
    .ap_loop_init(ap_loop_init),
    .ap_ready_int(ap_ready_int),
    .ap_loop_exit_ready(ap_condition_exit_pp0_iter1_stage0),
    .ap_loop_exit_done(ap_done_int),
    .ap_continue_int(ap_continue_int),
    .ap_done_int(ap_done_int)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue_int == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter2_reg == 1'b1))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b1 == ap_condition_exit_pp0_iter1_stage0)) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_enable_reg_pp0_iter1 <= ap_start_int;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready == 1'b0))) begin
        ap_loop_exit_ready_pp0_iter2_reg <= 1'b0;
    end else if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_loop_exit_ready_pp0_iter2_reg <= ap_loop_exit_ready;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        if ((ap_loop_init == 1'b1)) begin
            loop_index57_fu_60 <= 61'd0;
        end else if (((exitcond83_fu_126_p2 == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
            loop_index57_fu_60 <= empty_fu_114_p2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        loop_index57_load_reg_157 <= loop_index57_fu_60;
        mem_addr_read_reg_162 <= m_axi_mem_RDATA;
        sext_ln182_cast_reg_147 <= sext_ln182_cast_fu_98_p1;
    end
end

always @ (*) begin
    if (((exitcond83_fu_126_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_condition_exit_pp0_iter1_stage0 = 1'b1;
    end else begin
        ap_condition_exit_pp0_iter1_stage0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter2_reg == 1'b1))) begin
        ap_done_int = 1'b1;
    end else begin
        ap_done_int = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_idle_pp0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_start_int == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_ready_int = 1'b1;
    end else begin
        ap_ready_int = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        m_axi_mem_RREADY = 1'b1;
    end else begin
        m_axi_mem_RREADY = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        mem_blk_n_R = m_axi_mem_RVALID;
    end else begin
        mem_blk_n_R = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        node_cluster_assignments_ce1 = 1'b1;
    end else begin
        node_cluster_assignments_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        node_cluster_assignments_we1 = 1'b1;
    end else begin
        node_cluster_assignments_we1 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_pp0_stage0 : begin
            ap_NS_fsm = ap_ST_fsm_pp0_stage0;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_pp0_stage0_11001 = ((m_axi_mem_RVALID == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b1));
end

always @ (*) begin
    ap_block_pp0_stage0_subdone = ((m_axi_mem_RVALID == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b1));
end

assign ap_block_state1_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state2_pp0_stage0_iter1 = (m_axi_mem_RVALID == 1'b0);
end

assign ap_block_state3_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_enable_reg_pp0_iter0 = ap_start_int;

assign ap_loop_exit_ready = ap_condition_exit_pp0_iter1_stage0;

assign empty_fu_114_p2 = (loop_index57_fu_60 + 61'd1);

assign exitcond83_fu_126_p2 = ((empty_fu_114_p2 == sext_ln182_cast_reg_147) ? 1'b1 : 1'b0);

assign loop_index57_cast_fu_136_p1 = loop_index57_load_reg_157;

assign m_axi_mem_ARADDR = 64'd0;

assign m_axi_mem_ARBURST = 2'd0;

assign m_axi_mem_ARCACHE = 4'd0;

assign m_axi_mem_ARID = 1'd0;

assign m_axi_mem_ARLEN = 32'd0;

assign m_axi_mem_ARLOCK = 2'd0;

assign m_axi_mem_ARPROT = 3'd0;

assign m_axi_mem_ARQOS = 4'd0;

assign m_axi_mem_ARREGION = 4'd0;

assign m_axi_mem_ARSIZE = 3'd0;

assign m_axi_mem_ARUSER = 1'd0;

assign m_axi_mem_ARVALID = 1'b0;

assign m_axi_mem_AWADDR = 64'd0;

assign m_axi_mem_AWBURST = 2'd0;

assign m_axi_mem_AWCACHE = 4'd0;

assign m_axi_mem_AWID = 1'd0;

assign m_axi_mem_AWLEN = 32'd0;

assign m_axi_mem_AWLOCK = 2'd0;

assign m_axi_mem_AWPROT = 3'd0;

assign m_axi_mem_AWQOS = 4'd0;

assign m_axi_mem_AWREGION = 4'd0;

assign m_axi_mem_AWSIZE = 3'd0;

assign m_axi_mem_AWUSER = 1'd0;

assign m_axi_mem_AWVALID = 1'b0;

assign m_axi_mem_BREADY = 1'b0;

assign m_axi_mem_WDATA = 64'd0;

assign m_axi_mem_WID = 1'd0;

assign m_axi_mem_WLAST = 1'b0;

assign m_axi_mem_WSTRB = 8'd0;

assign m_axi_mem_WUSER = 1'd0;

assign m_axi_mem_WVALID = 1'b0;

assign node_cluster_assignments_address1 = loop_index57_cast_fu_136_p1;

assign node_cluster_assignments_d1 = mem_addr_read_reg_162;

assign sext_ln182_cast_fu_98_p1 = $signed(sext_ln182);

endmodule //kmeans_top_kmeans_top_Pipeline_3


// Content from kmeans_top_kmeans_Pipeline_3.v
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2022.2 (64-bit)
// Version: 2022.2
// Copyright (C) Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module kmeans_top_kmeans_Pipeline_3 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        centroid_x_coords_next_address0,
        centroid_x_coords_next_ce0,
        centroid_x_coords_next_we0,
        centroid_x_coords_next_d0,
        k_cast2_cast_cast
);

parameter    ap_ST_fsm_pp0_stage0 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
output  [7:0] centroid_x_coords_next_address0;
output   centroid_x_coords_next_ce0;
output   centroid_x_coords_next_we0;
output  [63:0] centroid_x_coords_next_d0;
input  [31:0] k_cast2_cast_cast;

reg ap_idle;
reg centroid_x_coords_next_ce0;
reg centroid_x_coords_next_we0;

(* fsm_encoding = "none" *) reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_enable_reg_pp0_iter0;
reg    ap_enable_reg_pp0_iter1;
reg    ap_idle_pp0;
wire    ap_block_state1_pp0_stage0_iter0;
wire    ap_block_state2_pp0_stage0_iter1;
wire    ap_block_pp0_stage0_subdone;
wire   [0:0] exitcond2_fu_71_p2;
reg    ap_condition_exit_pp0_iter1_stage0;
wire    ap_loop_exit_ready;
reg    ap_ready_int;
wire   [63:0] k_cast2_cast_cast_cast_cast_fu_52_p1;
reg   [63:0] k_cast2_cast_cast_cast_cast_reg_88;
wire    ap_block_pp0_stage0_11001;
wire    ap_block_pp0_stage0;
reg   [63:0] empty_fu_24;
wire   [63:0] empty_71_fu_65_p2;
wire    ap_loop_init;
wire  signed [60:0] k_cast2_cast_cast_cast_fu_48_p1;
reg    ap_done_reg;
wire    ap_continue_int;
reg    ap_done_int;
reg   [0:0] ap_NS_fsm;
wire    ap_enable_pp0;
wire    ap_start_int;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_CS_fsm = 1'd1;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_done_reg = 1'b0;
end

kmeans_top_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(ap_start),
    .ap_ready(ap_ready),
    .ap_done(ap_done),
    .ap_start_int(ap_start_int),
    .ap_loop_init(ap_loop_init),
    .ap_ready_int(ap_ready_int),
    .ap_loop_exit_ready(ap_condition_exit_pp0_iter1_stage0),
    .ap_loop_exit_done(ap_done_int),
    .ap_continue_int(ap_continue_int),
    .ap_done_int(ap_done_int)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue_int == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((ap_loop_exit_ready == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b1 == ap_condition_exit_pp0_iter1_stage0)) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_enable_reg_pp0_iter1 <= ap_start_int;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        if ((ap_loop_init == 1'b1)) begin
            empty_fu_24 <= 64'd0;
        end else if (((exitcond2_fu_71_p2 == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
            empty_fu_24 <= empty_71_fu_65_p2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        k_cast2_cast_cast_cast_cast_reg_88[60 : 0] <= k_cast2_cast_cast_cast_cast_fu_52_p1[60 : 0];
    end
end

always @ (*) begin
    if (((exitcond2_fu_71_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_condition_exit_pp0_iter1_stage0 = 1'b1;
    end else begin
        ap_condition_exit_pp0_iter1_stage0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_loop_exit_ready == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_done_int = 1'b1;
    end else begin
        ap_done_int = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_idle_pp0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_start_int == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_ready_int = 1'b1;
    end else begin
        ap_ready_int = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        centroid_x_coords_next_ce0 = 1'b1;
    end else begin
        centroid_x_coords_next_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        centroid_x_coords_next_we0 = 1'b1;
    end else begin
        centroid_x_coords_next_we0 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_pp0_stage0 : begin
            ap_NS_fsm = ap_ST_fsm_pp0_stage0;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

assign ap_block_state1_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_enable_reg_pp0_iter0 = ap_start_int;

assign ap_loop_exit_ready = ap_condition_exit_pp0_iter1_stage0;

assign centroid_x_coords_next_address0 = empty_fu_24;

assign centroid_x_coords_next_d0 = 64'd0;

assign empty_71_fu_65_p2 = (empty_fu_24 + 64'd1);

assign exitcond2_fu_71_p2 = ((empty_71_fu_65_p2 == k_cast2_cast_cast_cast_cast_reg_88) ? 1'b1 : 1'b0);

assign k_cast2_cast_cast_cast_cast_fu_52_p1 = $unsigned(k_cast2_cast_cast_cast_fu_48_p1);

assign k_cast2_cast_cast_cast_fu_48_p1 = $signed(k_cast2_cast_cast);

always @ (posedge ap_clk) begin
    k_cast2_cast_cast_cast_cast_reg_88[63:61] <= 3'b000;
end

endmodule //kmeans_top_kmeans_Pipeline_3


// Content from kmeans_top_kmeans_top_Pipeline_6.v
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2022.2 (64-bit)
// Version: 2022.2
// Copyright (C) Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module kmeans_top_kmeans_top_Pipeline_6 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        m_axi_mem_AWVALID,
        m_axi_mem_AWREADY,
        m_axi_mem_AWADDR,
        m_axi_mem_AWID,
        m_axi_mem_AWLEN,
        m_axi_mem_AWSIZE,
        m_axi_mem_AWBURST,
        m_axi_mem_AWLOCK,
        m_axi_mem_AWCACHE,
        m_axi_mem_AWPROT,
        m_axi_mem_AWQOS,
        m_axi_mem_AWREGION,
        m_axi_mem_AWUSER,
        m_axi_mem_WVALID,
        m_axi_mem_WREADY,
        m_axi_mem_WDATA,
        m_axi_mem_WSTRB,
        m_axi_mem_WLAST,
        m_axi_mem_WID,
        m_axi_mem_WUSER,
        m_axi_mem_ARVALID,
        m_axi_mem_ARREADY,
        m_axi_mem_ARADDR,
        m_axi_mem_ARID,
        m_axi_mem_ARLEN,
        m_axi_mem_ARSIZE,
        m_axi_mem_ARBURST,
        m_axi_mem_ARLOCK,
        m_axi_mem_ARCACHE,
        m_axi_mem_ARPROT,
        m_axi_mem_ARQOS,
        m_axi_mem_ARREGION,
        m_axi_mem_ARUSER,
        m_axi_mem_RVALID,
        m_axi_mem_RREADY,
        m_axi_mem_RDATA,
        m_axi_mem_RLAST,
        m_axi_mem_RID,
        m_axi_mem_RFIFONUM,
        m_axi_mem_RUSER,
        m_axi_mem_RRESP,
        m_axi_mem_BVALID,
        m_axi_mem_BREADY,
        m_axi_mem_BRESP,
        m_axi_mem_BID,
        m_axi_mem_BUSER,
        p_cast9_cast,
        node_cluster_assignments_address0,
        node_cluster_assignments_ce0,
        node_cluster_assignments_q0,
        sext_ln182
);

parameter    ap_ST_fsm_pp0_stage0 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
output   m_axi_mem_AWVALID;
input   m_axi_mem_AWREADY;
output  [63:0] m_axi_mem_AWADDR;
output  [0:0] m_axi_mem_AWID;
output  [31:0] m_axi_mem_AWLEN;
output  [2:0] m_axi_mem_AWSIZE;
output  [1:0] m_axi_mem_AWBURST;
output  [1:0] m_axi_mem_AWLOCK;
output  [3:0] m_axi_mem_AWCACHE;
output  [2:0] m_axi_mem_AWPROT;
output  [3:0] m_axi_mem_AWQOS;
output  [3:0] m_axi_mem_AWREGION;
output  [0:0] m_axi_mem_AWUSER;
output   m_axi_mem_WVALID;
input   m_axi_mem_WREADY;
output  [63:0] m_axi_mem_WDATA;
output  [7:0] m_axi_mem_WSTRB;
output   m_axi_mem_WLAST;
output  [0:0] m_axi_mem_WID;
output  [0:0] m_axi_mem_WUSER;
output   m_axi_mem_ARVALID;
input   m_axi_mem_ARREADY;
output  [63:0] m_axi_mem_ARADDR;
output  [0:0] m_axi_mem_ARID;
output  [31:0] m_axi_mem_ARLEN;
output  [2:0] m_axi_mem_ARSIZE;
output  [1:0] m_axi_mem_ARBURST;
output  [1:0] m_axi_mem_ARLOCK;
output  [3:0] m_axi_mem_ARCACHE;
output  [2:0] m_axi_mem_ARPROT;
output  [3:0] m_axi_mem_ARQOS;
output  [3:0] m_axi_mem_ARREGION;
output  [0:0] m_axi_mem_ARUSER;
input   m_axi_mem_RVALID;
output   m_axi_mem_RREADY;
input  [63:0] m_axi_mem_RDATA;
input   m_axi_mem_RLAST;
input  [0:0] m_axi_mem_RID;
input  [8:0] m_axi_mem_RFIFONUM;
input  [0:0] m_axi_mem_RUSER;
input  [1:0] m_axi_mem_RRESP;
input   m_axi_mem_BVALID;
output   m_axi_mem_BREADY;
input  [1:0] m_axi_mem_BRESP;
input  [0:0] m_axi_mem_BID;
input  [0:0] m_axi_mem_BUSER;
input  [60:0] p_cast9_cast;
output  [12:0] node_cluster_assignments_address0;
output   node_cluster_assignments_ce0;
input  [63:0] node_cluster_assignments_q0;
input  [31:0] sext_ln182;

reg ap_idle;
reg m_axi_mem_WVALID;
reg node_cluster_assignments_ce0;

(* fsm_encoding = "none" *) reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_enable_reg_pp0_iter0;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter2;
reg    ap_enable_reg_pp0_iter3;
reg    ap_idle_pp0;
wire    ap_block_state1_pp0_stage0_iter0;
wire    ap_block_state2_pp0_stage0_iter1;
wire    ap_block_state3_pp0_stage0_iter2;
wire    ap_block_state4_pp0_stage0_iter3;
reg    ap_block_pp0_stage0_subdone;
wire   [0:0] exitcond78_fu_126_p2;
reg    ap_condition_exit_pp0_iter1_stage0;
wire    ap_loop_exit_ready;
reg    ap_ready_int;
reg    mem_blk_n_W;
wire    ap_block_pp0_stage0;
wire  signed [60:0] sext_ln182_cast_fu_99_p1;
reg  signed [60:0] sext_ln182_cast_reg_149;
reg    ap_block_pp0_stage0_11001;
reg   [63:0] node_cluster_assignments_load_reg_168;
wire   [63:0] loop_index39_cast_fu_121_p1;
wire    ap_block_pp0_stage0_01001;
reg   [60:0] loop_index39_fu_62;
wire   [60:0] empty_fu_115_p2;
wire    ap_loop_init;
reg    ap_done_reg;
wire    ap_continue_int;
reg    ap_done_int;
reg    ap_loop_exit_ready_pp0_iter2_reg;
reg    ap_loop_exit_ready_pp0_iter3_reg;
reg   [0:0] ap_NS_fsm;
wire    ap_enable_pp0;
wire    ap_start_int;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_CS_fsm = 1'd1;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_done_reg = 1'b0;
end

kmeans_top_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(ap_start),
    .ap_ready(ap_ready),
    .ap_done(ap_done),
    .ap_start_int(ap_start_int),
    .ap_loop_init(ap_loop_init),
    .ap_ready_int(ap_ready_int),
    .ap_loop_exit_ready(ap_condition_exit_pp0_iter1_stage0),
    .ap_loop_exit_done(ap_done_int),
    .ap_continue_int(ap_continue_int),
    .ap_done_int(ap_done_int)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue_int == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter3_reg == 1'b1))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b1 == ap_condition_exit_pp0_iter1_stage0)) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_enable_reg_pp0_iter1 <= ap_start_int;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter2_reg == 1'b0))) begin
        ap_loop_exit_ready_pp0_iter3_reg <= 1'b0;
    end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        ap_loop_exit_ready_pp0_iter3_reg <= ap_loop_exit_ready_pp0_iter2_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        if ((ap_loop_init == 1'b1)) begin
            loop_index39_fu_62 <= 61'd0;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (exitcond78_fu_126_p2 == 1'd0))) begin
            loop_index39_fu_62 <= empty_fu_115_p2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_loop_exit_ready_pp0_iter2_reg <= ap_loop_exit_ready;
        sext_ln182_cast_reg_149 <= sext_ln182_cast_fu_99_p1;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        node_cluster_assignments_load_reg_168 <= node_cluster_assignments_q0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (exitcond78_fu_126_p2 == 1'd1))) begin
        ap_condition_exit_pp0_iter1_stage0 = 1'b1;
    end else begin
        ap_condition_exit_pp0_iter1_stage0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter3_reg == 1'b1))) begin
        ap_done_int = 1'b1;
    end else begin
        ap_done_int = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_idle_pp0 == 1'b1) & (ap_start_int == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_ready_int = 1'b1;
    end else begin
        ap_ready_int = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1))) begin
        m_axi_mem_WVALID = 1'b1;
    end else begin
        m_axi_mem_WVALID = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter3 == 1'b1))) begin
        mem_blk_n_W = m_axi_mem_WREADY;
    end else begin
        mem_blk_n_W = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        node_cluster_assignments_ce0 = 1'b1;
    end else begin
        node_cluster_assignments_ce0 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_pp0_stage0 : begin
            ap_NS_fsm = ap_ST_fsm_pp0_stage0;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_01001 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_pp0_stage0_11001 = ((m_axi_mem_WREADY == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b1));
end

always @ (*) begin
    ap_block_pp0_stage0_subdone = ((m_axi_mem_WREADY == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b1));
end

assign ap_block_state1_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_enable_reg_pp0_iter0 = ap_start_int;

assign ap_loop_exit_ready = ap_condition_exit_pp0_iter1_stage0;

assign empty_fu_115_p2 = (loop_index39_fu_62 + 61'd1);

assign exitcond78_fu_126_p2 = ((empty_fu_115_p2 == sext_ln182_cast_reg_149) ? 1'b1 : 1'b0);

assign loop_index39_cast_fu_121_p1 = loop_index39_fu_62;

assign m_axi_mem_ARADDR = 64'd0;

assign m_axi_mem_ARBURST = 2'd0;

assign m_axi_mem_ARCACHE = 4'd0;

assign m_axi_mem_ARID = 1'd0;

assign m_axi_mem_ARLEN = 32'd0;

assign m_axi_mem_ARLOCK = 2'd0;

assign m_axi_mem_ARPROT = 3'd0;

assign m_axi_mem_ARQOS = 4'd0;

assign m_axi_mem_ARREGION = 4'd0;

assign m_axi_mem_ARSIZE = 3'd0;

assign m_axi_mem_ARUSER = 1'd0;

assign m_axi_mem_ARVALID = 1'b0;

assign m_axi_mem_AWADDR = 64'd0;

assign m_axi_mem_AWBURST = 2'd0;

assign m_axi_mem_AWCACHE = 4'd0;

assign m_axi_mem_AWID = 1'd0;

assign m_axi_mem_AWLEN = 32'd0;

assign m_axi_mem_AWLOCK = 2'd0;

assign m_axi_mem_AWPROT = 3'd0;

assign m_axi_mem_AWQOS = 4'd0;

assign m_axi_mem_AWREGION = 4'd0;

assign m_axi_mem_AWSIZE = 3'd0;

assign m_axi_mem_AWUSER = 1'd0;

assign m_axi_mem_AWVALID = 1'b0;

assign m_axi_mem_BREADY = 1'b0;

assign m_axi_mem_RREADY = 1'b0;

assign m_axi_mem_WDATA = node_cluster_assignments_load_reg_168;

assign m_axi_mem_WID = 1'd0;

assign m_axi_mem_WLAST = 1'b0;

assign m_axi_mem_WSTRB = 8'd255;

assign m_axi_mem_WUSER = 1'd0;

assign node_cluster_assignments_address0 = loop_index39_cast_fu_121_p1;

assign sext_ln182_cast_fu_99_p1 = $signed(sext_ln182);

endmodule //kmeans_top_kmeans_top_Pipeline_6


// Content from kmeans_top_mem_m_axi.v
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2022.2 (64-bit)
// Version: 2022.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// ==============================================================
// 67d7842dbbe25473c3c32b93c0da8047785f30d78e8a024de1b57352245f9689

`timescale 1ns/1ps
`default_nettype none

module kmeans_top_mem_m_axi
#(parameter
    CONSERVATIVE            = 0,
    NUM_READ_OUTSTANDING    = 2,
    NUM_WRITE_OUTSTANDING   = 2,
    MAX_READ_BURST_LENGTH   = 16,
    MAX_WRITE_BURST_LENGTH  = 16,
    C_M_AXI_ID_WIDTH        = 1,
    C_M_AXI_ADDR_WIDTH      = 32,
    C_M_AXI_DATA_WIDTH      = 32, // power of 2 & range: 2 to 1024
    C_M_AXI_AWUSER_WIDTH    = 1,
    C_M_AXI_ARUSER_WIDTH    = 1,
    C_M_AXI_WUSER_WIDTH     = 1,
    C_M_AXI_RUSER_WIDTH     = 1,
    C_M_AXI_BUSER_WIDTH     = 1,
    C_TARGET_ADDR           = 32'h00000000,
    C_USER_VALUE            = 1'b0,
    C_PROT_VALUE            = 3'b000,
    C_CACHE_VALUE           = 4'b0011,
    USER_DW                 = 32, // multiple of 8
    USER_AW                 = 32,
    USER_MAXREQS            = 16,
    USER_RFIFONUM_WIDTH     = 6,
    MAXI_BUFFER_IMPL        = "block"
)(
    
    // system signal
    input  wire                               ACLK,
    input  wire                               ARESET,
    input  wire                               ACLK_EN,
    // write address channel
    output wire [C_M_AXI_ID_WIDTH-1:0]        AWID,
    output wire [C_M_AXI_ADDR_WIDTH-1:0]      AWADDR,
    output wire [7:0]                         AWLEN,
    output wire [2:0]                         AWSIZE,
    output wire [1:0]                         AWBURST,
    output wire [1:0]                         AWLOCK,
    output wire [3:0]                         AWCACHE,
    output wire [2:0]                         AWPROT,
    output wire [3:0]                         AWQOS,
    output wire [3:0]                         AWREGION,
    output wire [C_M_AXI_AWUSER_WIDTH-1:0]    AWUSER,
    output wire                               AWVALID,
    input  wire                               AWREADY,
    // write data channel
    output wire [C_M_AXI_ID_WIDTH-1:0]        WID,
    output wire [C_M_AXI_DATA_WIDTH-1:0]      WDATA,
    output wire [C_M_AXI_DATA_WIDTH/8-1:0]    WSTRB,
    output wire                               WLAST,
    output wire [C_M_AXI_WUSER_WIDTH-1:0]     WUSER,
    output wire                               WVALID,
    input  wire                               WREADY,
    // write response channel
    input  wire [C_M_AXI_ID_WIDTH-1:0]        BID,
    input  wire [1:0]                         BRESP,
    input  wire [C_M_AXI_BUSER_WIDTH-1:0]     BUSER,
    input  wire                               BVALID,
    output wire                               BREADY,
    // read address channel
    output wire [C_M_AXI_ID_WIDTH-1:0]        ARID,
    output wire [C_M_AXI_ADDR_WIDTH-1:0]      ARADDR,
    output wire [7:0]                         ARLEN,
    output wire [2:0]                         ARSIZE,
    output wire [1:0]                         ARBURST,
    output wire [1:0]                         ARLOCK,
    output wire [3:0]                         ARCACHE,
    output wire [2:0]                         ARPROT,
    output wire [3:0]                         ARQOS,
    output wire [3:0]                         ARREGION,
    output wire [C_M_AXI_ARUSER_WIDTH-1:0]    ARUSER,
    output wire                               ARVALID,
    input  wire                               ARREADY,
    // read data channel
    input  wire [C_M_AXI_ID_WIDTH-1:0]        RID,
    input  wire [C_M_AXI_DATA_WIDTH-1:0]      RDATA,
    input  wire [1:0]                         RRESP,
    input  wire                               RLAST,
    input  wire [C_M_AXI_RUSER_WIDTH-1:0]     RUSER,
    input  wire                               RVALID,
    output wire                               RREADY,

    // internal bus ports
    // write address
    input  wire [USER_AW-1:0]                 I_AWADDR,
    input  wire [31:0]                        I_AWLEN,
    input  wire                               I_AWVALID,
    output wire                               I_AWREADY,
    // write data
    input  wire [USER_DW-1:0]                 I_WDATA,
    input  wire [USER_DW/8-1:0]               I_WSTRB,
    input  wire                               I_WVALID,
    output wire                               I_WREADY,
    // write response
    output wire                               I_BVALID,
    input  wire                               I_BREADY,
    // read address
    input  wire [USER_AW-1:0]                 I_ARADDR,
    input  wire [31:0]                        I_ARLEN,
    input  wire                               I_ARVALID,
    output wire                               I_ARREADY,
    // read data
    output wire [USER_DW-1:0]                 I_RDATA,
    output wire                               I_RVALID,
    input  wire                               I_RREADY,
    output wire [USER_RFIFONUM_WIDTH-1:0]     I_RFIFONUM);
//------------------------Local signal-------------------

    wire [C_M_AXI_ADDR_WIDTH-1:0]   AWADDR_Dummy;
    wire [31:0]                     AWLEN_Dummy;
    wire                            AWVALID_Dummy;
    wire                            AWREADY_Dummy;
    wire [C_M_AXI_DATA_WIDTH-1:0]   WDATA_Dummy;
    wire [C_M_AXI_DATA_WIDTH/8-1:0] WSTRB_Dummy;
    wire                            WVALID_Dummy;
    wire                            WREADY_Dummy;
    wire                            BVALID_Dummy;
    wire                            BREADY_Dummy;
    wire [C_M_AXI_ADDR_WIDTH-1:0]   ARADDR_Dummy;
    wire [31:0]                     ARLEN_Dummy;
    wire                            ARVALID_Dummy;
    wire                            ARREADY_Dummy;
    wire [C_M_AXI_DATA_WIDTH-1:0]   RDATA_Dummy;
    wire [1:0]                      RLAST_Dummy;
    wire                            RVALID_Dummy;
    wire                            RREADY_Dummy;
    wire                            RBURST_READY_Dummy;
    
//------------------------Instantiation------------------
    // kmeans_top_mem_m_axi_store
    kmeans_top_mem_m_axi_store #(
        .C_TARGET_ADDR           ( C_TARGET_ADDR ),
        .NUM_WRITE_OUTSTANDING   ( NUM_WRITE_OUTSTANDING ),
        .MAX_WRITE_BURST_LENGTH  ( MAX_WRITE_BURST_LENGTH ),
        .BUS_ADDR_WIDTH          ( C_M_AXI_ADDR_WIDTH ),
        .BUS_DATA_WIDTH          ( C_M_AXI_DATA_WIDTH ),
        .USER_DW                 ( USER_DW ),
        .USER_AW                 ( USER_AW ),
        .USER_MAXREQS            ( USER_MAXREQS ),
        .BUFFER_IMPL             ( MAXI_BUFFER_IMPL )
    ) store_unit (
        .ACLK                    ( ACLK ),
        .ARESET                  ( ARESET ),
        .ACLK_EN                 ( ACLK_EN ),
        .out_AXI_AWADDR          ( AWADDR_Dummy ),
        .out_AXI_AWLEN           ( AWLEN_Dummy ),
        .out_AXI_AWVALID         ( AWVALID_Dummy ),
        .in_AXI_AWREADY          ( AWREADY_Dummy ),
        .out_AXI_WDATA           ( WDATA_Dummy ),
        .out_AXI_WSTRB           ( WSTRB_Dummy ),
        .out_AXI_WVALID          ( WVALID_Dummy ),
        .in_AXI_WREADY           ( WREADY_Dummy ),
        .in_AXI_BVALID           ( BVALID_Dummy ),
        .out_AXI_BREADY          ( BREADY_Dummy ),
        .in_HLS_AWADDR           ( I_AWADDR ),
        .in_HLS_AWLEN            ( I_AWLEN ),
        .in_HLS_AWVALID          ( I_AWVALID ),
        .out_HLS_AWREADY         ( I_AWREADY ),
        .in_HLS_WDATA            ( I_WDATA ),
        .in_HLS_WSTRB            ( I_WSTRB ),
        .in_HLS_WVALID           ( I_WVALID ),
        .out_HLS_WREADY          ( I_WREADY ),
        .out_HLS_BVALID          ( I_BVALID ),
        .in_HLS_BREADY           ( I_BREADY ));

    // kmeans_top_mem_m_axi_load
    kmeans_top_mem_m_axi_load #(
        .C_TARGET_ADDR           ( C_TARGET_ADDR ),
        .NUM_READ_OUTSTANDING    ( NUM_READ_OUTSTANDING ),
        .MAX_READ_BURST_LENGTH   ( MAX_READ_BURST_LENGTH ),
        .BUS_ADDR_WIDTH          ( C_M_AXI_ADDR_WIDTH ),
        .BUS_DATA_WIDTH          ( C_M_AXI_DATA_WIDTH ),
        .USER_DW                 ( USER_DW ),
        .USER_AW                 ( USER_AW ),
        .USER_MAXREQS            ( USER_MAXREQS ),
        .USER_RFIFONUM_WIDTH     ( USER_RFIFONUM_WIDTH ),
        .BUFFER_IMPL             ( MAXI_BUFFER_IMPL )
    ) load_unit (
        .ACLK                    ( ACLK ),
        .ARESET                  ( ARESET ),
        .ACLK_EN                 ( ACLK_EN ),
        .out_AXI_ARADDR          ( ARADDR_Dummy ),
        .out_AXI_ARLEN           ( ARLEN_Dummy ),
        .out_AXI_ARVALID         ( ARVALID_Dummy ),
        .in_AXI_ARREADY          ( ARREADY_Dummy ),
        .in_AXI_RDATA            ( RDATA_Dummy ),
        .in_AXI_RLAST            ( RLAST_Dummy ),
        .in_AXI_RVALID           ( RVALID_Dummy ),
        .out_AXI_RREADY          ( RREADY_Dummy ),
        .out_AXI_RBURST_READY    ( RBURST_READY_Dummy),
        .in_HLS_ARADDR           ( I_ARADDR ),
        .in_HLS_ARLEN            ( I_ARLEN ),
        .in_HLS_ARVALID          ( I_ARVALID ),
        .out_HLS_ARREADY         ( I_ARREADY ),
        .out_HLS_RDATA           ( I_RDATA ),
        .out_HLS_RVALID          ( I_RVALID ),
        .in_HLS_RREADY           ( I_RREADY ),
        .out_HLS_RFIFONUM        ( I_RFIFONUM ));

    // kmeans_top_mem_m_axi_write
    kmeans_top_mem_m_axi_write #(
        .CONSERVATIVE            ( CONSERVATIVE),
        .C_M_AXI_ID_WIDTH        ( C_M_AXI_ID_WIDTH ),
        .C_M_AXI_AWUSER_WIDTH    ( C_M_AXI_AWUSER_WIDTH ),
        .C_M_AXI_WUSER_WIDTH     ( C_M_AXI_WUSER_WIDTH ),
        .C_M_AXI_BUSER_WIDTH     ( C_M_AXI_BUSER_WIDTH ),
        .C_USER_VALUE            ( C_USER_VALUE ),
        .C_PROT_VALUE            ( C_PROT_VALUE ),
        .C_CACHE_VALUE           ( C_CACHE_VALUE ),
        .BUS_ADDR_WIDTH          ( C_M_AXI_ADDR_WIDTH ),
        .BUS_DATA_WIDTH          ( C_M_AXI_DATA_WIDTH ),
        .NUM_WRITE_OUTSTANDING   ( NUM_WRITE_OUTSTANDING ),
        .MAX_WRITE_BURST_LENGTH  ( MAX_WRITE_BURST_LENGTH )
    ) bus_write (
        .ACLK                    ( ACLK ),
        .ARESET                  ( ARESET ),
        .ACLK_EN                 ( ACLK_EN ),
        .out_BUS_AWID            ( AWID ),
        .out_BUS_AWSIZE          ( AWSIZE ),
        .out_BUS_AWBURST         ( AWBURST ),
        .out_BUS_AWLOCK          ( AWLOCK ),
        .out_BUS_AWCACHE         ( AWCACHE ),
        .out_BUS_AWPROT          ( AWPROT ),
        .out_BUS_AWQOS           ( AWQOS ),
        .out_BUS_AWREGION        ( AWREGION ),
        .out_BUS_AWUSER          ( AWUSER ),
        .out_BUS_AWADDR          ( AWADDR ),
        .out_BUS_AWLEN           ( AWLEN ),
        
        
        .out_BUS_AWVALID         ( AWVALID ),
        .in_BUS_AWREADY          ( AWREADY ),
        .out_BUS_WID             ( WID),
        .out_BUS_WUSER           ( WUSER),
        .out_BUS_WDATA           ( WDATA ),
        .out_BUS_WSTRB           ( WSTRB ),
        .out_BUS_WLAST           ( WLAST ),
        
        
        .out_BUS_WVALID          ( WVALID ),
        .in_BUS_WREADY           ( WREADY ),
        .in_BUS_BID              ( BID ),
        .in_BUS_BRESP            ( BRESP ),
        .in_BUS_BUSER            ( BUSER ),
        .in_BUS_BVALID           ( BVALID ),
        
        
        .out_BUS_BREADY          ( BREADY ),
        .in_HLS_AWVALID          ( AWVALID_Dummy ),
        .out_HLS_AWREADY         ( AWREADY_Dummy ),
        .in_HLS_AWADDR           ( AWADDR_Dummy ),
        .in_HLS_AWLEN            ( AWLEN_Dummy ),
        .in_HLS_WVALID           ( WVALID_Dummy ),
        .out_HLS_WREADY          ( WREADY_Dummy ),
        .in_HLS_WSTRB            ( WSTRB_Dummy ),
        .in_HLS_WDATA            ( WDATA_Dummy ),
        .out_HLS_BVALID          ( BVALID_Dummy ),
        .in_HLS_BREADY           ( BREADY_Dummy ));

    // kmeans_top_mem_m_axi_read
    kmeans_top_mem_m_axi_read #(
        .C_M_AXI_ID_WIDTH         ( C_M_AXI_ID_WIDTH ),
        .C_M_AXI_ARUSER_WIDTH     ( C_M_AXI_ARUSER_WIDTH ),
        .C_M_AXI_RUSER_WIDTH      ( C_M_AXI_RUSER_WIDTH ),
        .C_USER_VALUE             ( C_USER_VALUE ),
        .C_PROT_VALUE             ( C_PROT_VALUE ),
        .C_CACHE_VALUE            ( C_CACHE_VALUE ),
        .BUS_ADDR_WIDTH           ( C_M_AXI_ADDR_WIDTH ),
        .BUS_DATA_WIDTH           ( C_M_AXI_DATA_WIDTH ),
        .NUM_READ_OUTSTANDING     ( NUM_READ_OUTSTANDING ),
        .MAX_READ_BURST_LENGTH    ( MAX_READ_BURST_LENGTH )
    ) bus_read (
        .ACLK                     ( ACLK ),
        .ARESET                   ( ARESET ),
        .ACLK_EN                  ( ACLK_EN ),
        .out_BUS_ARID             ( ARID ),
        .out_BUS_ARADDR           ( ARADDR ),
        .out_BUS_ARLEN            ( ARLEN ),
        .out_BUS_ARSIZE           ( ARSIZE ),
        .out_BUS_ARBURST          ( ARBURST ),
        .out_BUS_ARLOCK           ( ARLOCK ),
        .out_BUS_ARCACHE          ( ARCACHE ),
        .out_BUS_ARPROT           ( ARPROT ),
        .out_BUS_ARQOS            ( ARQOS ),
        .out_BUS_ARREGION         ( ARREGION ),
        .out_BUS_ARUSER           ( ARUSER ),
        
        
        .out_BUS_ARVALID          ( ARVALID ),
        .in_BUS_ARREADY           ( ARREADY ),
        .in_BUS_RID               ( RID ),
        .in_BUS_RDATA             ( RDATA ),
        .in_BUS_RRESP             ( RRESP ),
        .in_BUS_RLAST             ( RLAST ),
        .in_BUS_RUSER             ( RUSER ),
        .in_BUS_RVALID            ( RVALID ),
        
        
        .out_BUS_RREADY           ( RREADY ),
        .in_HLS_ARVALID           ( ARVALID_Dummy ),
        .out_HLS_ARREADY          ( ARREADY_Dummy ),
        .in_HLS_ARADDR            ( ARADDR_Dummy ),
        .in_HLS_ARLEN             ( ARLEN_Dummy ),
        .out_HLS_RVALID           ( RVALID_Dummy ),
        .in_HLS_RREADY            ( RREADY_Dummy ),
        .in_HLS_RBUST_READY       ( RBURST_READY_Dummy),
        .out_HLS_RDATA            ( RDATA_Dummy ),
        .out_HLS_RLAST            ( RLAST_Dummy ));

    
endmodule
`default_nettype wire// 67d7842dbbe25473c3c32b93c0da8047785f30d78e8a024de1b57352245f9689

`timescale 1ns/1ps

module kmeans_top_mem_m_axi_load
#(parameter
    C_TARGET_ADDR                         = 32'h00000000,
    NUM_READ_OUTSTANDING                  = 2,
    MAX_READ_BURST_LENGTH                 = 16,
    BUS_ADDR_WIDTH                        = 32,
    BUS_DATA_WIDTH                        = 32,
    USER_DW                               = 16,
    USER_AW                               = 32,
    USER_MAXREQS                          = 16,
    USER_RFIFONUM_WIDTH                   = 6,
    BUFFER_IMPL                           = "auto"
)(
    // system signal
    input  wire                           ACLK,
    input  wire                           ARESET,
    input  wire                           ACLK_EN,

    // read address channel
    output wire [BUS_ADDR_WIDTH-1:0]      out_AXI_ARADDR,
    output wire [31:0]                    out_AXI_ARLEN,
    output wire                           out_AXI_ARVALID,
    input  wire                           in_AXI_ARREADY,
    // read data channel
    input  wire [BUS_DATA_WIDTH-1:0]      in_AXI_RDATA,
    input  wire [1:0]                     in_AXI_RLAST,
    input  wire                           in_AXI_RVALID,
    output wire                           out_AXI_RREADY,
    output wire                           out_AXI_RBURST_READY,

    // internal bus ports
    // read address
    input  wire [USER_AW-1:0]             in_HLS_ARADDR,
    input  wire [31:0]                    in_HLS_ARLEN,
    input  wire                           in_HLS_ARVALID,
    output wire                           out_HLS_ARREADY,
    // read data
    output wire [USER_DW-1:0]             out_HLS_RDATA,
    output wire                           out_HLS_RVALID,
    input  wire                           in_HLS_RREADY,
    output wire [USER_RFIFONUM_WIDTH-1:0] out_HLS_RFIFONUM);

//------------------------Parameter----------------------
    localparam
        USER_DATA_WIDTH = calc_data_width(USER_DW),
        USER_DATA_BYTES = USER_DATA_WIDTH / 8,
        USER_ADDR_ALIGN = log2(USER_DATA_BYTES),
        BUS_ADDR_ALIGN  = log2(BUS_DATA_WIDTH/8),
        RBUFF_DEPTH     = NUM_READ_OUTSTANDING * MAX_READ_BURST_LENGTH,
        TARGET_ADDR     = C_TARGET_ADDR & (32'hffffffff << USER_ADDR_ALIGN);

//------------------------Task and function--------------
    function integer calc_data_width;
        input integer x;
        integer y;
    begin
        y = 8;
        while (y < x) y = y * 2;
        calc_data_width = y;
    end
    endfunction

    function integer log2;
        input integer x;
        integer n, m;
    begin
        n = 0;
        m = 1;
        while (m < x) begin
            n = n + 1;
            m = m * 2;
        end
        log2 = n;
    end
    endfunction

//------------------------Local signal-------------------

    wire                           next_rreq;
    wire                           ready_for_rreq;
    wire                           rreq_ready;

    wire [USER_AW-1 : 0]           rreq_addr;
    wire [31:0]                    rreq_len;
    wire                           rreq_valid;

    wire                           valid_length;

    reg  [BUS_ADDR_WIDTH-1 : 0]    tmp_addr;
    reg  [31:0]                    tmp_len;
    reg                            tmp_valid;

    wire                           burst_ready;
    wire                           beat_valid;
    wire                           next_beat;
    wire                           last_beat;
    wire [BUS_DATA_WIDTH-1 : 0]    beat_data;
    wire [log2(RBUFF_DEPTH) : 0]   beat_nvalid;

    reg                            ready_for_outstanding;

//------------------------Instantiation------------------
    kmeans_top_mem_m_axi_fifo #(
        .DATA_WIDTH        (USER_AW + 32),
        .ADDR_WIDTH        (log2(USER_MAXREQS)),
        .DEPTH             (USER_MAXREQS)
    ) fifo_rreq (
        .clk               (ACLK),
        .reset             (ARESET),
        .clk_en            (ACLK_EN),
        .if_full_n         (out_HLS_ARREADY),
        .if_write          (in_HLS_ARVALID),
        .if_din            ({in_HLS_ARLEN, in_HLS_ARADDR}),
        .if_empty_n        (rreq_valid),
        .if_read           (next_rreq),
        .if_dout           ({rreq_len, rreq_addr}),
        .if_num_data_valid ());

    // ===================================================================
    // start of ARADDR PREPROCESSOR
    
    assign next_rreq       = rreq_valid && ready_for_rreq;
    assign ready_for_rreq  = ~tmp_valid || (in_AXI_ARREADY && rreq_ready);

    assign valid_length    = (rreq_len != 32'b0) && !rreq_len[31];

    assign out_AXI_ARLEN   = tmp_len;   // Byte length
    assign out_AXI_ARADDR  = tmp_addr;  // Byte address
    assign out_AXI_ARVALID = tmp_valid && rreq_ready;

    always @(posedge ACLK)
    begin
        if (ARESET) begin
            tmp_len  <= 0;
            tmp_addr <= 0;
        end
        else if (ACLK_EN) begin
            if(next_rreq) begin
                tmp_len  <= (rreq_len << USER_ADDR_ALIGN) - 1;            // byte length
                tmp_addr <= TARGET_ADDR + (rreq_addr << USER_ADDR_ALIGN); // byte address
            end
        end
    end
 
    always @(posedge ACLK) 
    begin
        if (ARESET)
            tmp_valid <= 1'b0;
        else if (ACLK_EN) begin
            if (next_rreq && valid_length)
                tmp_valid <= 1'b1;
            else if (in_AXI_ARREADY && rreq_ready)
                tmp_valid <= 1'b0;
        end
    end

    // end of ARADDR PREPROCESSOR
    // ===================================================================

    kmeans_top_mem_m_axi_fifo #(
        .MEM_STYLE         (BUFFER_IMPL),
        .DATA_WIDTH        (BUS_DATA_WIDTH + 2),
        .ADDR_WIDTH        (log2(RBUFF_DEPTH)),
        .DEPTH             (RBUFF_DEPTH)
    ) buff_rdata (
        .clk               (ACLK),
        .reset             (ARESET),
        .clk_en            (ACLK_EN),
        .if_full_n         (out_AXI_RREADY),
        .if_write          (in_AXI_RVALID),
        .if_din            ({in_AXI_RLAST, in_AXI_RDATA}),
        .if_empty_n        (beat_valid),
        .if_read           (next_beat),
        .if_dout           ({burst_ready, last_beat, beat_data}),
        .if_num_data_valid (beat_nvalid));

    assign out_AXI_RBURST_READY = ready_for_outstanding;

    always @(posedge ACLK) 
    begin
        if (ARESET)
            ready_for_outstanding <= 1'b0;
        else if (ACLK_EN) begin
            if (next_beat)
                ready_for_outstanding <= burst_ready;
            else
                ready_for_outstanding <= 1'b0;
        end
    end
    // ===================================================================
    // start of RDATA PREPROCESSOR
    generate
    if (USER_DATA_WIDTH == BUS_DATA_WIDTH) begin : bus_equal_gen

        assign rreq_ready       = 1'b1;
        assign next_beat        = in_HLS_RREADY;

        assign out_HLS_RDATA    = beat_data[USER_DW-1 : 0];
        assign out_HLS_RVALID   = beat_valid;
        assign out_HLS_RFIFONUM = beat_nvalid;

    end
    else if (USER_DATA_WIDTH < BUS_DATA_WIDTH) begin : bus_wide_gen
        localparam
            TOTAL_SPLIT  = BUS_DATA_WIDTH / USER_DATA_WIDTH,
            SPLIT_ALIGN  = log2(TOTAL_SPLIT);

        wire [USER_AW - 1:0]        tmp_addr_end;

        wire                        offset_full_n;
        wire                        offset_write;
        wire [SPLIT_ALIGN-1 : 0]    start_offset;
        wire [SPLIT_ALIGN-1 : 0]    end_offset;

        wire                        offset_valid;
        wire                        next_offset;
        wire [SPLIT_ALIGN-1 : 0]    head_offset;
        wire [SPLIT_ALIGN-1 : 0]    tail_offset;

        reg                         first_beat;

        wire                        first_data;
        wire                        last_data;
        wire                        ready_for_data;

        reg  [BUS_DATA_WIDTH-1 : 0] data_buf;
        reg                         data_valid;

        reg  [USER_RFIFONUM_WIDTH-1:0] rdata_nvalid; 
        reg  [SPLIT_ALIGN : 0]      data_nvalid;
        wire [SPLIT_ALIGN : 0]      split_nvalid;
        
        wire [SPLIT_ALIGN-1 : 0]    split_cnt;
        reg  [SPLIT_ALIGN-1 : 0]    split_cnt_buf;

        wire                        first_split;
        wire                        next_split;
        wire                        last_split;

        // Recording the offset of start & end address to extract the expect data from beats when USER_DW < BUS_DW.
        kmeans_top_mem_m_axi_fifo #(
            .DATA_WIDTH         (2*SPLIT_ALIGN),
            .ADDR_WIDTH         (log2(NUM_READ_OUTSTANDING)),
            .DEPTH              (NUM_READ_OUTSTANDING)
        ) rreq_offset (
            .clk                (ACLK),
            .reset              (ARESET),
            .clk_en             (ACLK_EN),
            .if_full_n          (offset_full_n),
            .if_write           (offset_write),
            .if_din             ({start_offset, end_offset}),
            .if_empty_n         (offset_valid),
            .if_read            (next_offset),
            .if_dout            ({head_offset, tail_offset}),
            .if_num_data_valid  ());

        assign rreq_ready       = offset_full_n | ~offset_write;
        assign tmp_addr_end     = tmp_addr + tmp_len;

        assign start_offset     = tmp_addr[BUS_ADDR_ALIGN - 1 : 0] >> USER_ADDR_ALIGN;
        assign end_offset       = tmp_addr_end[BUS_ADDR_ALIGN - 1 : 0] >> USER_ADDR_ALIGN;
        assign offset_write     = tmp_valid & in_AXI_ARREADY;

        assign next_offset      = (last_beat & beat_valid) & last_split;
        assign next_beat        = last_split;

        assign out_HLS_RDATA    = data_buf[USER_DW-1 : 0];
        assign out_HLS_RVALID   = data_valid;
        assign out_HLS_RFIFONUM = rdata_nvalid + data_nvalid;

        assign ready_for_data   = ~data_valid | in_HLS_RREADY;
        assign first_data       = first_beat && beat_valid && offset_valid;
        assign last_data        = last_beat && beat_valid && offset_valid;

        assign first_split      = (~first_data) ? (split_cnt == 0 && beat_valid && ready_for_data) : ((split_cnt == head_offset) && ready_for_data);
        assign last_split       = (~last_data)  ? (split_cnt == (TOTAL_SPLIT-1) && ready_for_data) : ((split_cnt == tail_offset) && ready_for_data);
        assign next_split       = (~first_data) ? (split_cnt != 0 && ready_for_data)               : ((split_cnt != head_offset) && ready_for_data);

        assign split_cnt        = (first_data && (split_cnt_buf == 0)) ? head_offset : split_cnt_buf;

        assign split_nvalid     = (first_data && last_data)  ? tail_offset - head_offset + 1 :
                                   first_data                ? TOTAL_SPLIT - head_offset     :
                                   last_data                 ? tail_offset + 1               :
                                   TOTAL_SPLIT;
        always @(posedge ACLK)
        begin
            if (ARESET)
                split_cnt_buf <= 0;
            else if (ACLK_EN) begin 
                if (last_split)
                    split_cnt_buf <= 0;
                else if (first_split || next_split)
                    split_cnt_buf <= split_cnt + 1;
            end
        end

        always @(posedge ACLK)
        begin
            if (ARESET)
                first_beat <= 1'b1;
            else if (ACLK_EN) begin
                if (last_beat && last_split)
                    first_beat <= 1'b1;
                else if (first_beat && last_split)
                    first_beat <= 1'b0;
            end
        end

        always @(posedge ACLK)
        begin
            if (ACLK_EN) begin
                if (first_split & first_data)
                    data_buf <= beat_data >> (head_offset * USER_DATA_WIDTH);
                else if (first_split)
                    data_buf <= beat_data;
                else if (next_split)
                    data_buf <= data_buf >> USER_DATA_WIDTH;
            end
        end

        always @(posedge ACLK)
        begin
            if (ARESET)
                data_valid <= 1'b0;
            else if (ACLK_EN) begin
                if (first_split)
                    data_valid <= 1'b1;
                else if (~(first_split || next_split) && ready_for_data)
                    data_valid <= 1'b0;
            end
        end

        always @(posedge ACLK)
        begin
            if (ARESET)
                data_nvalid <= 0;
            else if (ACLK_EN) begin
                if (first_split)
                    data_nvalid <= split_nvalid;
                else if (next_split)
                    data_nvalid <= data_nvalid - 1;
                else if (~(first_split || next_split) && ready_for_data)
                    data_nvalid <= 0;
            end
        end

        always @(posedge ACLK)
        begin
            if (ARESET)
                rdata_nvalid <= 0;
            else if (ACLK_EN) begin
                if (!beat_valid)
                    rdata_nvalid <= 0;
                else
                    rdata_nvalid <= ((beat_nvalid - 1) << SPLIT_ALIGN);
            end
        end
        
    end
    else begin : bus_narrow_gen
        localparam
            TOTAL_PADS      = USER_DATA_WIDTH / BUS_DATA_WIDTH,
            PAD_ALIGN       = log2(TOTAL_PADS);

        reg [USER_DATA_WIDTH-1 : 0] data_buf;
        reg                         data_valid;
        reg [PAD_ALIGN:0]           data_nvalid;
        wire                        ready_for_data;

        wire [TOTAL_PADS - 1:0]     pad_oh;
        reg  [TOTAL_PADS - 1:0]     pad_oh_reg;

        reg                         first_pad;
        wire                        last_pad;
        wire                        next_pad;

        assign rreq_ready       = 1'b1; 
        assign next_beat        = next_pad;
        
        assign out_HLS_RDATA    = data_buf[USER_DW-1 : 0];
        assign out_HLS_RVALID   = data_valid;
        assign out_HLS_RFIFONUM = beat_nvalid[log2(RBUFF_DEPTH) : PAD_ALIGN] + (beat_nvalid[PAD_ALIGN-1:0] + data_nvalid) >> PAD_ALIGN;
        assign ready_for_data   = ~data_valid | in_HLS_RREADY;

        assign next_pad         = beat_valid && ready_for_data;
        assign last_pad         = pad_oh[TOTAL_PADS - 1];

        always @(posedge ACLK)
        begin
            if (ARESET)
                first_pad <= 1'b1;
            else if (ACLK_EN) begin
                if (next_pad && ~last_pad)
                    first_pad <= 1'b0;
                else if (next_pad && last_pad)
                    first_pad <= 1'b1;
            end
        end

        assign pad_oh = (beat_valid == 0)  ?  0 :
                        (first_pad)        ?  1 :
                        pad_oh_reg;
 
        always @(posedge ACLK)
        begin
            if (ARESET)
                pad_oh_reg <= 0;
            else if (ACLK_EN) begin
                if (next_pad)
                    pad_oh_reg <= {pad_oh[TOTAL_PADS - 2:0], 1'b0};
            end
        end

        genvar  i;
        for (i = 0; i < TOTAL_PADS; i = i + 1) begin : data_gen
            always @(posedge ACLK)
            begin
                if (ACLK_EN) begin
                    if (pad_oh[i] == 1'b1 && ready_for_data)
                        data_buf[i*BUS_DATA_WIDTH +: BUS_DATA_WIDTH] <= beat_data;
                end
            end
        end

        always @(posedge ACLK)
        begin
            if (ARESET)
                data_valid <= 1'b0;
            else if (ACLK_EN) begin
                if (next_beat)
                    data_valid <= 1'b1;
                else if (ready_for_data)
                    data_valid <= 1'b0;
            end
        end

        always @(posedge ACLK)
        begin
            if (ARESET)
                data_nvalid <= 0;
            else if (ACLK_EN) begin
                if (first_pad)
                    data_nvalid <= 1;
                else if (next_pad)
                    data_nvalid <= data_nvalid + 1;
            end
        end

    end
    endgenerate
    // end of RDATA PREPROCESSOR
    // ===================================================================

endmodule


module kmeans_top_mem_m_axi_store
#(parameter
    C_TARGET_ADDR           = 32'h00000000,
    NUM_WRITE_OUTSTANDING   = 2,
    MAX_WRITE_BURST_LENGTH  = 16,
    BUS_ADDR_WIDTH          = 32,
    BUS_DATA_WIDTH          = 32,
    USER_DW                 = 16,
    USER_AW                 = 32,
    USER_MAXREQS            = 16,
    BUFFER_IMPL             = "auto"
)(
    // system signal
    input  wire                        ACLK,
    input  wire                        ARESET,
    input  wire                        ACLK_EN,
    // write address channel
    output wire [BUS_ADDR_WIDTH-1:0]   out_AXI_AWADDR,
    output wire [31:0]                 out_AXI_AWLEN,
    output wire                        out_AXI_AWVALID,
    input  wire                        in_AXI_AWREADY,
    // write data channel
    output wire [BUS_DATA_WIDTH-1:0]   out_AXI_WDATA,
    output wire [BUS_DATA_WIDTH/8-1:0] out_AXI_WSTRB,
    output wire                        out_AXI_WVALID,
    input  wire                        in_AXI_WREADY,
    // write response channel
    input  wire                        in_AXI_BVALID,
    output wire                        out_AXI_BREADY,

    // internal bus ports
    // write address
    input  wire [USER_AW-1:0]          in_HLS_AWADDR,
    input  wire [31:0]                 in_HLS_AWLEN,
    input  wire                        in_HLS_AWVALID,
    output wire                        out_HLS_AWREADY,
    // write data
    input  wire [USER_DW-1:0]          in_HLS_WDATA,
    input  wire [USER_DW/8-1:0]        in_HLS_WSTRB,
    input  wire                        in_HLS_WVALID,
    output wire                        out_HLS_WREADY,
    // write response
    output wire                        out_HLS_BVALID,
    input  wire                        in_HLS_BREADY);

//------------------------Parameter----------------------
    localparam
        USER_DATA_WIDTH = calc_data_width(USER_DW),
        USER_DATA_BYTES = USER_DATA_WIDTH / 8,
        USER_ADDR_ALIGN = log2(USER_DATA_BYTES),
        BUS_DATA_BYTES  = BUS_DATA_WIDTH / 8,
        BUS_ADDR_ALIGN  = log2(BUS_DATA_BYTES),
        // write buffer size 
        WBUFF_DEPTH     = max(MAX_WRITE_BURST_LENGTH * BUS_DATA_WIDTH / USER_DATA_WIDTH, 1),  
        TARGET_ADDR     = C_TARGET_ADDR & (32'hffffffff << USER_ADDR_ALIGN); 

//------------------------Task and function--------------

    function integer max;
        input integer x;
        input integer y;
    begin
        max = (x > y) ? x : y;
    end
    endfunction

    function integer calc_data_width;
        input integer x;
        integer y;
    begin
        y = 8;
        while (y < x) y = y * 2;
        calc_data_width = y;
    end
    endfunction

    function integer log2;
        input integer x;
        integer n, m;
    begin
        n = 0;
        m = 1;
        while (m < x) begin
            n = n + 1;
            m = m * 2;
        end
        log2 = n;
    end
    endfunction

//------------------------Local signal-------------------

    wire                                next_wreq;
    wire                                ready_for_wreq;
    wire                                wreq_ready;

    wire [USER_AW-1 : 0]                wreq_addr;
    wire [31:0]                         wreq_len;
    wire                                wreq_valid;

    wire                                valid_length;

    reg  [USER_AW-1 : 0]                tmp_addr;
    reg  [31:0]                         tmp_len;
    reg                                 tmp_valid;

    wire                                next_wdata;
    wire                                wdata_valid;
    wire [USER_DW-1 : 0]                tmp_wdata;
    wire [USER_DW/8-1 : 0]              tmp_wstrb;

    wire                                wrsp_ready;
    wire                                wrsp_valid;
    wire                                wrsp_read;
    wire                                wrsp_type;

    wire                                ursp_ready;
    wire                                ursp_write;

//------------------------Instantiation------------------
    kmeans_top_mem_m_axi_fifo #(
        .DATA_WIDTH     (USER_AW + 32),
        .ADDR_WIDTH     (log2(USER_MAXREQS)),
        .DEPTH          (USER_MAXREQS)
    ) fifo_wreq (
        .clk            (ACLK),
        .reset          (ARESET),
        .clk_en         (ACLK_EN),
        .if_full_n      (out_HLS_AWREADY),
        .if_write       (in_HLS_AWVALID),
        .if_din         ({in_HLS_AWLEN, in_HLS_AWADDR}),
        .if_empty_n     (wreq_valid),
        .if_read        (next_wreq),
        .if_dout        ({wreq_len, wreq_addr}),
        .if_num_data_valid());

    assign next_wreq = wreq_valid && ready_for_wreq && wrsp_ready;
    assign ready_for_wreq  = ~tmp_valid || (in_AXI_AWREADY && wreq_ready);

    assign valid_length    = (wreq_len != 32'b0) && !wreq_len[31];

    assign out_AXI_AWLEN   = tmp_len;   // Byte length
    assign out_AXI_AWADDR  = tmp_addr;  // Byte address
    assign out_AXI_AWVALID = tmp_valid && wreq_ready;

    always @(posedge ACLK)
    begin
        if (ARESET) begin
            tmp_len  <= 0;
            tmp_addr <= 0;
        end
        else if (ACLK_EN) begin
            if(next_wreq) begin
                tmp_len  <= (wreq_len << USER_ADDR_ALIGN) - 1;
                tmp_addr <= TARGET_ADDR + (wreq_addr << USER_ADDR_ALIGN);
            end
        end
    end
 
    always @(posedge ACLK) 
    begin
        if (ARESET)
            tmp_valid <= 1'b0;
        else if (next_wreq && valid_length)
            tmp_valid <= 1'b1;
        else if (in_AXI_AWREADY && wreq_ready)
            tmp_valid <= 1'b0;
    end

    // ===================================================================

    kmeans_top_mem_m_axi_fifo #(
        .MEM_STYLE         (BUFFER_IMPL),
        .DATA_WIDTH        (USER_DW + USER_DW/8),
        .ADDR_WIDTH        (log2(WBUFF_DEPTH)),
        .DEPTH             (WBUFF_DEPTH)
    ) buff_wdata (
        .clk               (ACLK),
        .reset             (ARESET),
        .clk_en            (ACLK_EN),
        .if_full_n         (out_HLS_WREADY),
        .if_write          (in_HLS_WVALID),
        .if_din            ({in_HLS_WSTRB , in_HLS_WDATA}),
        .if_empty_n        (wdata_valid),
        .if_read           (next_wdata),
        .if_dout           ({tmp_wstrb, tmp_wdata}),
        .if_num_data_valid ());

    generate
    if (USER_DATA_WIDTH == BUS_DATA_WIDTH) begin : bus_equal_gen
        assign next_wdata       = in_AXI_WREADY;
        assign out_AXI_WVALID   = wdata_valid;
        assign out_AXI_WDATA    = tmp_wdata;
        assign out_AXI_WSTRB    = tmp_wstrb;

        assign wreq_ready   = 1'b1;

    end
    else if (USER_DATA_WIDTH < BUS_DATA_WIDTH) begin : bus_wide_gen
        localparam
            TOTAL_PADS      = BUS_DATA_WIDTH / USER_DATA_WIDTH,
            PAD_ALIGN       = log2(TOTAL_PADS),
            BEAT_LEN_WIDTH  = 32 - BUS_ADDR_ALIGN;

        function [TOTAL_PADS-1 : 0] decoder;
            input [PAD_ALIGN-1 : 0] din;
            reg  [TOTAL_PADS-1 : 0] dout;
            integer i;
        begin
            dout = {TOTAL_PADS{1'b0}};
            i = 0;
            while (i < din) begin
                dout[i] = 1'b1;
                i = i + 1;
            end
            decoder = dout;
        end
        endfunction

        wire [USER_AW - 1:0]        tmp_addr_end;

        wire                        offset_full_n;
        wire                        offset_write;
        wire [PAD_ALIGN-1 : 0]      start_offset;
        wire [PAD_ALIGN-1 : 0]      end_offset;
        wire [BEAT_LEN_WIDTH-1 : 0] beat_total;

        wire                        offset_valid;
        wire                        next_offset;
        wire [PAD_ALIGN-1 : 0]      head_offset;
        wire [PAD_ALIGN-1 : 0]      tail_offset;

        wire [BEAT_LEN_WIDTH-1 : 0] beat_len;
        reg  [BEAT_LEN_WIDTH-1:0]   len_cnt;

        wire [TOTAL_PADS - 1:0]     add_head;
        wire [TOTAL_PADS - 1:0]     add_tail;
        wire [TOTAL_PADS - 1:0]     pad_oh;
        reg  [TOTAL_PADS - 1:0]     pad_oh_reg;

        reg [TOTAL_PADS-1 : 0]     head_pad_sel;
        reg [0 : TOTAL_PADS-1]     tail_pad_sel; // reverse
        wire                        ready_for_data;
        wire                        next_pad;
        reg                         first_pad;
        wire                        last_pad;
        wire                        first_beat;
        wire                        last_beat;
        wire                        next_beat;

        reg  [BUS_DATA_WIDTH - 1:0] data_buf;
        reg  [BUS_DATA_BYTES - 1:0] strb_buf;
        reg                         data_valid;

        // Recording the offset of start & end address to align beats from data USER_DW < BUS_DW.
        kmeans_top_mem_m_axi_fifo #(
            .DATA_WIDTH             (2*PAD_ALIGN + BEAT_LEN_WIDTH),
            .ADDR_WIDTH             (log2(NUM_WRITE_OUTSTANDING)),
            .DEPTH                  (NUM_WRITE_OUTSTANDING)
        ) wreq_offset (
            .clk                    (ACLK),
            .reset                  (ARESET),
            .clk_en                 (ACLK_EN),
            .if_full_n              (offset_full_n),
            .if_write               (offset_write),
            .if_din                 ({start_offset, end_offset, beat_total}),
            .if_empty_n             (offset_valid),
            .if_read                (next_offset),
            .if_dout                ({head_offset, tail_offset, beat_len}),
            .if_num_data_valid      ());

        assign wreq_ready   = offset_full_n | ~offset_write;
        assign tmp_addr_end = tmp_addr + tmp_len;

        assign start_offset   = tmp_addr[BUS_ADDR_ALIGN-1 : 0] >> USER_ADDR_ALIGN;
        assign end_offset     = ~tmp_addr_end[BUS_ADDR_ALIGN-1 : 0] >> USER_ADDR_ALIGN;
        assign beat_total     = (tmp_len + tmp_addr[BUS_ADDR_ALIGN-1 : 0]) >> BUS_ADDR_ALIGN;

        assign offset_write   = tmp_valid & in_AXI_AWREADY;

        assign out_AXI_WDATA  = data_buf;
        assign out_AXI_WSTRB  = strb_buf;
        assign out_AXI_WVALID = data_valid;

        assign next_wdata     = next_pad;
        assign next_offset    = last_beat && next_beat;
        assign ready_for_data = ~data_valid || in_AXI_WREADY;

        assign first_beat     = (len_cnt == 0) && offset_valid;
        assign last_beat      = (len_cnt == beat_len) && offset_valid;
        assign next_beat      = offset_valid && last_pad && ready_for_data;

        assign next_pad       = offset_valid && wdata_valid && ready_for_data;
        assign last_pad       = (last_beat) ? pad_oh[TOTAL_PADS-tail_offset-1] : pad_oh[TOTAL_PADS-1];

        // assign head_pad_sel   = decoder(head_offset);
        // assign tail_pad_sel   = decoder(tail_offset);

        always @(*) begin
            integer i;
            head_pad_sel = {TOTAL_PADS{1'b0}};
            for (i = 0; i < TOTAL_PADS; i = i + 1) begin
                if (i < head_offset)
                    head_pad_sel[i] = 1'b1;
                else
                    head_pad_sel[i] = 1'b0;
            end
        end

        always @(*) begin
            integer i;
            tail_pad_sel = {TOTAL_PADS{1'b0}};
            for (i = 0; i < TOTAL_PADS; i = i + 1) begin
                if (i < tail_offset)
                    tail_pad_sel[i] = 1'b1;
                else
                    tail_pad_sel[i] = 1'b0;
            end

        end

        always @(posedge ACLK)
        begin
            if (ARESET)
                len_cnt <= 0;
            else if (ACLK_EN) begin
                if (next_offset)
                    len_cnt <= 0;
                else if (next_beat)
                    len_cnt <= len_cnt + 1;
            end
        end

        always @(posedge ACLK)
        begin
            if (ARESET)
                first_pad <= 1'b1;
            else if (ACLK_EN) begin
                if (next_pad && ~last_pad)
                    first_pad <= 1'b0;
                else if (next_pad && last_pad)
                    first_pad <= 1'b1;
            end
        end 
        
        assign pad_oh = (~wdata_valid)            ? 0                :
                        (first_pad && first_beat) ? 1 << head_offset :
                        (first_pad)?                1                :
                        pad_oh_reg;

        always @(posedge ACLK)
        begin
            if (ARESET)
                pad_oh_reg <= 0;
            else if (ACLK_EN) begin
                if (next_pad)
                    pad_oh_reg <= {pad_oh[TOTAL_PADS - 2:0], 1'b0};
            end
        end

        genvar  i;
        for (i = 0; i < TOTAL_PADS; i = i + 1) begin : data_gen
            assign add_head[i] = head_pad_sel[i] && first_beat;
            assign add_tail[i] = tail_pad_sel[i] && last_beat;

            always @(posedge ACLK)
            begin
                if (ARESET)
                    data_buf[i*USER_DATA_WIDTH +: USER_DATA_WIDTH] <= {USER_DATA_WIDTH{1'b0}};
                else if (ACLK_EN) begin
                    if ((add_head[i] || add_tail[i]) && ready_for_data)
                        data_buf[i*USER_DATA_WIDTH +: USER_DATA_WIDTH] <= {USER_DATA_WIDTH{1'b0}};
                    else if (pad_oh[i] == 1'b1 && ready_for_data)
                        data_buf[i*USER_DATA_WIDTH +: USER_DATA_WIDTH] <= tmp_wdata;
                end
            end

            always @(posedge ACLK)
            begin
                if (ARESET)
                    strb_buf[i*USER_DATA_BYTES +: USER_DATA_BYTES] <= {USER_DATA_BYTES{1'b0}};
                else if (ACLK_EN) begin
                    if ((add_head[i] || add_tail[i]) && ready_for_data)
                        strb_buf[i*USER_DATA_BYTES +: USER_DATA_BYTES] <= {USER_DATA_BYTES{1'b0}};
                    else if (pad_oh[i] == 1'b1 && ready_for_data)
                        strb_buf[i*USER_DATA_BYTES +: USER_DATA_BYTES] <= tmp_wstrb;
                end
            end

        end

        always @(posedge ACLK)
        begin
            if (ARESET)
                data_valid <= 1'b0;
            else if (ACLK_EN) begin
                if (next_beat)
                    data_valid <= 1'b1;
                else if (ready_for_data)
                    data_valid <= 1'b0;
            end
        end

    end
    else begin : bus_narrow_gen
        localparam
            TOTAL_SPLIT       = USER_DATA_WIDTH / BUS_DATA_WIDTH,
            SPLIT_ALIGN       = log2(TOTAL_SPLIT),
            BEAT_LEN_WIDTH    = 32 - BUS_ADDR_ALIGN;


        wire [USER_AW - 1:0]        tmp_addr_end;

        wire                        offset_full_n;
        wire                        offset_write;
        wire  [BEAT_LEN_WIDTH-1 : 0] beat_total;

        wire                        offset_valid;
        wire                        next_offset;

        wire [BEAT_LEN_WIDTH-1 : 0] beat_len;
        reg  [BEAT_LEN_WIDTH-1 : 0] len_cnt;

        wire                        ready_for_data;
        reg  [BUS_DATA_WIDTH - 1:0] data_buf;
        reg  [BUS_DATA_BYTES - 1:0] strb_buf;
        reg                         data_valid;

        reg [SPLIT_ALIGN-1 : 0]     split_cnt;

        wire                        first_split;
        wire                        next_split;
        wire                        last_split;

        // Recording the offset of start & end address to align beats from data USER_DW < BUS_DW.
        kmeans_top_mem_m_axi_fifo #(
            .DATA_WIDTH        (BEAT_LEN_WIDTH),
            .ADDR_WIDTH        (log2(NUM_WRITE_OUTSTANDING)),
            .DEPTH             (NUM_WRITE_OUTSTANDING)
        ) wreq_offset (
            .clk               (ACLK),
            .reset             (ARESET),
            .clk_en            (ACLK_EN),
            .if_full_n         (offset_full_n),
            .if_write          (offset_write),
            .if_din            (beat_total),
            .if_empty_n        (offset_valid),
            .if_read           (next_offset),
            .if_dout           (beat_len),
            .if_num_data_valid ());

        assign wreq_ready     = offset_full_n | ~offset_write;
        assign beat_total     = (tmp_len + tmp_addr[BUS_ADDR_ALIGN-1 : 0]) >> BUS_ADDR_ALIGN;

        assign offset_write   = tmp_valid & in_AXI_AWREADY;

        assign out_AXI_WDATA  = data_buf[BUS_DATA_WIDTH - 1:0];
        assign out_AXI_WSTRB  = strb_buf[BUS_DATA_BYTES - 1:0];
        assign out_AXI_WVALID = data_valid;

        assign next_wdata     = first_split;
        assign next_offset    = (len_cnt == beat_len) && offset_valid && last_split;
        assign ready_for_data = ~data_valid | in_AXI_WREADY;

        assign first_split    = (split_cnt == 0) && wdata_valid && offset_valid && ready_for_data;
        assign last_split     = (split_cnt == (TOTAL_SPLIT - 1)) && ready_for_data;
        assign next_split     = (split_cnt != 0) && ready_for_data;
        
        always @(posedge ACLK)
        begin
            if (ARESET)
                split_cnt <= 0;
            else if (ACLK_EN) begin
                if (last_split)
                    split_cnt <= 0;
                else if (first_split || next_split)
                    split_cnt <= split_cnt + 1;
            end
        end

        always @(posedge ACLK)
        begin
            if (ARESET)
                len_cnt <= 0;
            else if (ACLK_EN) begin
                if (next_offset)
                    len_cnt <= 0;
                else if (next_wdata || next_split)
                    len_cnt <= len_cnt + 1;
            end
        end
 
        always @(posedge ACLK)
        begin
            if (ACLK_EN) begin
                if (next_wdata)
                    data_buf <= tmp_wdata;
                else if (next_split)
                    data_buf <= data_buf >> BUS_DATA_WIDTH;
            end
        end

        always @(posedge ACLK)
        begin
            if (ARESET)
                strb_buf <= 0;
            else if (ACLK_EN) begin
                if (next_wdata)
                    strb_buf <= tmp_wstrb;
                else if (next_split)
                    strb_buf <= strb_buf >> BUS_DATA_BYTES;
            end
        end

        always @(posedge ACLK)
        begin
            if (ARESET)
                data_valid <= 0;
            else if (ACLK_EN) begin
                if (next_wdata)
                    data_valid <= 1;
                else if (~(first_split || next_split) && ready_for_data)
                    data_valid <= 0;
            end
        end
    end
    endgenerate

    // ===================================================================

    // generate response for all request (including request with invalid length)
    kmeans_top_mem_m_axi_fifo #(
        .DATA_WIDTH        (1),
        .ADDR_WIDTH        (log2(NUM_WRITE_OUTSTANDING)),
        .DEPTH             (NUM_WRITE_OUTSTANDING)
    ) fifo_wrsp (
        .clk               (ACLK),
        .reset             (ARESET),
        .clk_en            (ACLK_EN),
        .if_full_n         (wrsp_ready),
        .if_write          (next_wreq),
        .if_din            (valid_length),
        .if_empty_n        (wrsp_valid),
        .if_read           (wrsp_read),
        .if_dout           (wrsp_type), // 1 - valid length request, 0 - invalid length request
        .if_num_data_valid ());

    kmeans_top_mem_m_axi_fifo #(
        .DATA_WIDTH        (1),
        .ADDR_WIDTH        (log2(USER_MAXREQS)),
        .DEPTH             (USER_MAXREQS)
    ) user_resp (
        .clk               (ACLK),
        .reset             (ARESET),
        .clk_en            (ACLK_EN),
        .if_full_n         (ursp_ready),
        .if_write          (ursp_write),
        .if_din            (1'b1),
        .if_empty_n        (out_HLS_BVALID),
        .if_read           (in_HLS_BREADY),
        .if_dout           (),
        .if_num_data_valid ());

    assign ursp_write  = wrsp_valid && (!wrsp_type || in_AXI_BVALID);
    assign wrsp_read   = ursp_ready && ursp_write;

    assign out_AXI_BREADY = wrsp_type && ursp_ready;

endmodule

// 67d7842dbbe25473c3c32b93c0da8047785f30d78e8a024de1b57352245f9689

`timescale 1ns/1ps

//


module kmeans_top_mem_m_axi_read
#(parameter
    C_M_AXI_ID_WIDTH          = 1,
    C_M_AXI_ARUSER_WIDTH      = 1,
    C_M_AXI_RUSER_WIDTH       = 1,
    C_USER_VALUE              = 1'b0,
    C_PROT_VALUE              = 3'b000,
    C_CACHE_VALUE             = 4'b0011,
    BUS_ADDR_WIDTH            = 32,
    BUS_DATA_WIDTH            = 32,
    NUM_READ_OUTSTANDING      = 2,
    MAX_READ_BURST_LENGTH     = 16
)(
    // system signal
    input  wire                            ACLK,
    input  wire                            ARESET,
    input  wire                            ACLK_EN,
    // read address channel
    output wire [C_M_AXI_ID_WIDTH-1:0]     out_BUS_ARID,
    output wire [BUS_ADDR_WIDTH-1:0]       out_BUS_ARADDR,
    output wire [7:0]                      out_BUS_ARLEN,
    output wire [2:0]                      out_BUS_ARSIZE,
    output wire [1:0]                      out_BUS_ARBURST,
    output wire [1:0]                      out_BUS_ARLOCK,
    output wire [3:0]                      out_BUS_ARCACHE,
    output wire [2:0]                      out_BUS_ARPROT,
    output wire [3:0]                      out_BUS_ARQOS,
    output wire [3:0]                      out_BUS_ARREGION,
    output wire [C_M_AXI_ARUSER_WIDTH-1:0] out_BUS_ARUSER,
    output wire                            out_BUS_ARVALID,
    input  wire                            in_BUS_ARREADY,
    // read data channel
    input  wire [C_M_AXI_ID_WIDTH-1:0]     in_BUS_RID,
    input  wire [BUS_DATA_WIDTH-1:0]       in_BUS_RDATA,
    input  wire [1:0]                      in_BUS_RRESP,
    input  wire                            in_BUS_RLAST,
    input  wire [C_M_AXI_RUSER_WIDTH-1:0]  in_BUS_RUSER,
    input  wire                            in_BUS_RVALID,
    output wire                            out_BUS_RREADY,

    // HLS internal read request channel
    input  wire [BUS_ADDR_WIDTH-1:0]       in_HLS_ARADDR,
    input  wire [31:0]                     in_HLS_ARLEN,
    input  wire                            in_HLS_ARVALID,
    output wire                            out_HLS_ARREADY,
    output wire [BUS_DATA_WIDTH-1:0]       out_HLS_RDATA,
    output wire [1:0]                      out_HLS_RLAST,
    output wire                            out_HLS_RVALID,
    input  wire                            in_HLS_RREADY,
    input  wire                            in_HLS_RBUST_READY);

//------------------------Parameter----------------------
    localparam
        BUS_DATA_BYTES  = BUS_DATA_WIDTH / 8,
        BUS_ADDR_ALIGN  = log2(BUS_DATA_BYTES),
        NUM_READ_WIDTH  = log2(MAX_READ_BURST_LENGTH),
        RBUFFER_AWIDTH  = log2(MAX_READ_BURST_LENGTH*NUM_READ_OUTSTANDING),
        BOUNDARY_BEATS  = {12-BUS_ADDR_ALIGN{1'b1}};

//------------------------Task and function--------------
    function integer calc_data_width;
        input integer x;
        integer y;
    begin
        y = 8;
        while (y < x) y = y * 2;
        calc_data_width = y;
    end
    endfunction

    function integer log2;
        input integer x;
        integer n, m;
    begin
        n = 0;
        m = 1;
        while (m < x) begin
            n = n + 1;
            m = m * 2;
        end
        log2 = n;
    end
    endfunction

//------------------------Local signal-------------------
    // AR channel
    wire                                rreq_valid;
    wire [BUS_ADDR_WIDTH - 1:0]         tmp_addr;
    wire [31:0]                         tmp_len;
    wire [7:0]                          arlen_tmp;
    wire [BUS_ADDR_WIDTH - 1:0]         araddr_tmp;
    reg  [BUS_ADDR_WIDTH - 1:0]         start_addr;
    reg  [BUS_ADDR_WIDTH - 1:0]         end_addr;
    wire [BUS_ADDR_WIDTH - 1:0]         sect_addr;
    reg  [BUS_ADDR_WIDTH - 1:0]         sect_addr_buf;
    wire [11 - BUS_ADDR_ALIGN:0]        start_to_4k;
    wire [11 - BUS_ADDR_ALIGN:0]        sect_len;
    reg  [11 - BUS_ADDR_ALIGN:0]        sect_len_buf;
    reg  [11 - BUS_ADDR_ALIGN:0]        beat_len;
    reg  [BUS_ADDR_WIDTH - 13:0]        sect_cnt;
    wire                                ar2r_info;
    wire                                fifo_rctl_r;
    wire                                fifo_burst_w;
    reg                                 ARVALID_Dummy;
    wire                                ready_for_sect;
    wire                                next_rreq;
    wire                                ready_for_rreq;
    reg                                 rreq_handling;
    wire                                first_sect;
    wire                                last_sect;
    reg                                 last_sect_buf;
    wire                                next_sect;
    // R channel
    wire [BUS_DATA_WIDTH-1:0]           tmp_data;
    wire                                tmp_last;
    wire                                data_valid;
    wire                                data_ready;
    wire                                next_ctrl;
    wire                                need_rlast;
    wire                                burst_valid;
    wire                                last_burst;
    wire                                fifo_rctl_ready;
    wire                                next_burst;
    wire                                burst_end;

//------------------------AR channel begin---------------
//------------------------Instantiation------------------
    kmeans_top_mem_m_axi_reg_slice #(
        .DATA_WIDTH     (BUS_ADDR_WIDTH + 32)
    ) rs_rreq (
        .clk            (ACLK),
        .reset          (ARESET),
        .s_data         ({in_HLS_ARLEN, in_HLS_ARADDR}),
        .s_valid        (in_HLS_ARVALID),
        .s_ready        (out_HLS_ARREADY),
        .m_data         ({tmp_len, tmp_addr}),
        .m_valid        (rreq_valid),
        .m_ready        (next_rreq));

//------------------------Body---------------------------   
    assign ready_for_rreq = last_sect & next_sect | ~rreq_handling;
    assign next_rreq      = rreq_valid & ready_for_rreq;

    always @(posedge ACLK)
    begin
        if (ARESET) begin
            start_addr <= 0;
            end_addr   <= 0;
            beat_len   <= 0;
        end
        else if (ACLK_EN) begin
            if(next_rreq) begin
                start_addr <= tmp_addr;
                end_addr   <= tmp_addr + tmp_len;
                beat_len   <= (tmp_len[11:0] + tmp_addr[BUS_ADDR_ALIGN-1:0]) >> BUS_ADDR_ALIGN;
            end
        end
    end

    always @(posedge ACLK)
    begin
        if (ARESET)
            rreq_handling <= 1'b0;
        else if (ACLK_EN) begin
            if (rreq_valid && ~rreq_handling)
                rreq_handling <= 1'b1;
            else if (~rreq_valid && last_sect && next_sect)
                rreq_handling <= 1'b0;
        end
    end

    assign first_sect = (sect_cnt == start_addr[BUS_ADDR_WIDTH-1:12]);
    assign last_sect  = (sect_cnt == end_addr[BUS_ADDR_WIDTH-1:12]);
    assign next_sect  = rreq_handling & ready_for_sect;

    assign sect_addr  = (first_sect)? start_addr : {sect_cnt, {12{1'b0}}};
    assign start_to_4k = BOUNDARY_BEATS - start_addr[11:BUS_ADDR_ALIGN];
    assign sect_len    = ( first_sect &&  last_sect)? beat_len :
                         ( first_sect && ~last_sect)? start_to_4k:
                         (~first_sect &&  last_sect)? end_addr[11:BUS_ADDR_ALIGN] :
                                                      BOUNDARY_BEATS;

    always @(posedge ACLK)
    begin
        if (ARESET)
            sect_cnt <= 0;
        else if (ACLK_EN) begin
            if (next_rreq)
                sect_cnt <= tmp_addr[BUS_ADDR_WIDTH-1:12];
            else if (next_sect)
                sect_cnt <= sect_cnt + 1;
        end
    end

    always @(posedge ACLK)
    begin
        if (ARESET) begin
            sect_addr_buf <= 0;
            sect_len_buf <= 0;
            last_sect_buf <= 1'b0;
        end
        else if (ACLK_EN) begin
            if (next_sect) begin
                sect_addr_buf <= sect_addr;
                sect_len_buf <= sect_len;
                last_sect_buf <= last_sect;
            end
        end
    end

    assign out_BUS_ARID     = 0;
    assign out_BUS_ARSIZE   = BUS_ADDR_ALIGN;
    assign out_BUS_ARBURST  = 2'b01;
    assign out_BUS_ARLOCK   = 2'b00;
    assign out_BUS_ARCACHE  = C_CACHE_VALUE;
    assign out_BUS_ARPROT   = C_PROT_VALUE;
    assign out_BUS_ARUSER   = C_USER_VALUE;
    assign out_BUS_ARQOS    = 4'b0000;
    assign out_BUS_ARREGION = 4'b0000;

    generate
    if (BUS_DATA_BYTES >= 4096/MAX_READ_BURST_LENGTH) begin : must_one_burst
        assign out_BUS_ARADDR  = {sect_addr_buf[BUS_ADDR_WIDTH - 1:BUS_ADDR_ALIGN], {BUS_ADDR_ALIGN{1'b0}}};
        assign out_BUS_ARLEN   = sect_len_buf;
        assign out_BUS_ARVALID = ARVALID_Dummy;

        assign ready_for_sect = ~(ARVALID_Dummy && ~in_BUS_ARREADY) && fifo_rctl_ready;

        always @(posedge ACLK)
        begin
            if (ARESET)
                ARVALID_Dummy <= 1'b0;
            else if (ACLK_EN) begin
                if (next_sect)
                    ARVALID_Dummy <= 1'b1;
                else if (~next_sect && in_BUS_ARREADY)
                    ARVALID_Dummy <= 1'b0;
            end
        end

        assign fifo_rctl_r  = next_sect;
        assign ar2r_info    = last_sect;

        assign fifo_burst_w = next_sect;
        assign araddr_tmp   = sect_addr[BUS_ADDR_WIDTH - 1:0];
        assign arlen_tmp    = sect_len;
    end
    else begin : could_multi_bursts
        reg  [BUS_ADDR_WIDTH - 1:0]                     araddr_buf;
        reg  [7:0]                                      arlen_buf;
        reg  [11 - NUM_READ_WIDTH - BUS_ADDR_ALIGN:0]   loop_cnt;
        reg                                             sect_handling;
        wire                                            last_loop;
        wire                                            next_loop;
        wire                                            ready_for_loop;

        assign out_BUS_ARADDR  = araddr_buf;
        assign out_BUS_ARLEN   = arlen_buf;
        assign out_BUS_ARVALID = ARVALID_Dummy;

        assign last_loop      = (loop_cnt == sect_len_buf[11 - BUS_ADDR_ALIGN : NUM_READ_WIDTH]);
        assign next_loop      = sect_handling && ready_for_loop;
        assign ready_for_loop = ~(ARVALID_Dummy && ~in_BUS_ARREADY) && fifo_rctl_ready;
        assign ready_for_sect = ~(sect_handling && ~(last_loop && next_loop));

        always @(posedge ACLK)
        begin
            if (ARESET)
                sect_handling <= 1'b0;
            else if (ACLK_EN) begin
                if (rreq_handling && ~sect_handling)
                    sect_handling <= 1'b1;
                else if (~rreq_handling && last_loop && next_loop)
                    sect_handling <= 1'b0;
            end
        end

        always @(posedge ACLK)
        begin
            if (ARESET)
                loop_cnt <= 0;
            else if (ACLK_EN) begin
                if (next_sect)
                    loop_cnt <= 0;
                else if (next_loop)
                    loop_cnt <= loop_cnt + 1;
            end
        end

        assign araddr_tmp = (loop_cnt == 0)? sect_addr_buf[BUS_ADDR_WIDTH - 1:0] : (araddr_buf + ((arlen_buf + 1) << BUS_ADDR_ALIGN));
        assign arlen_tmp  = (NUM_READ_WIDTH == 0) ? 0 :
                            (last_loop)? sect_len_buf[NUM_READ_WIDTH - 1:0] : { NUM_READ_WIDTH{1'b1} };
        always @(posedge ACLK)
        begin
            if (ARESET) begin
                araddr_buf <= 0;
                arlen_buf <= 0;
            end
            else if (ACLK_EN) begin
                if (next_loop) begin
                    araddr_buf <= {araddr_tmp[BUS_ADDR_WIDTH - 1:BUS_ADDR_ALIGN], {BUS_ADDR_ALIGN{1'b0}}};
                    arlen_buf <= arlen_tmp;
                end
            end
        end

        always @(posedge ACLK)
        begin
            if (ARESET)
                ARVALID_Dummy <= 1'b0;
            else if (ACLK_EN) begin
                if (next_loop)
                    ARVALID_Dummy <= 1'b1;
                else if (~next_loop && in_BUS_ARREADY)
                    ARVALID_Dummy <= 1'b0;
            end
        end

        assign fifo_rctl_r  = next_loop;
        assign ar2r_info    = last_loop && last_sect_buf;

        assign fifo_burst_w = next_loop;
    end
    endgenerate
//------------------------AR channel end-----------------

//------------------------R channel begin----------------
//------------------------Instantiation------------------
    kmeans_top_mem_m_axi_reg_slice #(
        .DATA_WIDTH     (BUS_DATA_WIDTH + 1)
    ) rs_rdata (
        .clk            (ACLK),
        .reset          (ARESET),
        .s_data         ({in_BUS_RLAST, in_BUS_RDATA}),
        .s_valid        (in_BUS_RVALID),
        .s_ready        (out_BUS_RREADY),
        .m_data         ({tmp_last, tmp_data}),
        .m_valid        (data_valid),
        .m_ready        (data_ready));

    kmeans_top_mem_m_axi_fifo #(
        .DATA_WIDTH     (1),
        .ADDR_WIDTH     (log2(NUM_READ_OUTSTANDING)),
        .DEPTH          (NUM_READ_OUTSTANDING)
    ) fifo_rctl (
        .clk            (ACLK),
        .reset          (ARESET),
        .clk_en         (ACLK_EN),
        .if_full_n      (fifo_rctl_ready),
        .if_write       (fifo_rctl_r),
        .if_din         (ar2r_info),
        .if_empty_n     (need_rlast),
        .if_read        (next_ctrl),
        .if_dout        (),
        .if_num_data_valid());

    kmeans_top_mem_m_axi_fifo #(
        .DATA_WIDTH     (1),
        .ADDR_WIDTH     (log2(NUM_READ_OUTSTANDING)),
        .DEPTH          (NUM_READ_OUTSTANDING)
    ) fifo_burst (
        .clk            (ACLK),
        .reset          (ARESET),
        .clk_en         (ACLK_EN),
        .if_full_n      (),
        .if_write       (fifo_rctl_r),
        .if_din         (ar2r_info),
        .if_empty_n     (burst_valid),
        .if_read        (next_burst),
        .if_dout        (last_burst),
        .if_num_data_valid());

//------------------------Body---------------------------
    assign next_ctrl      = in_HLS_RBUST_READY && need_rlast;
    assign next_burst     = burst_end && data_valid && data_ready;

    assign burst_end      = tmp_last === 1'b1;
    assign out_HLS_RLAST  = {burst_end, burst_end && last_burst && burst_valid};
    assign out_HLS_RDATA  = tmp_data;
    assign out_HLS_RVALID = data_valid;
    assign data_ready     = in_HLS_RREADY;
//------------------------R channel end------------------
endmodule

module kmeans_top_mem_m_axi_write
#(parameter
    CONSERVATIVE              = 0,
    C_M_AXI_ID_WIDTH          = 1,
    C_M_AXI_AWUSER_WIDTH      = 1,
    C_M_AXI_WUSER_WIDTH       = 1,
    C_M_AXI_BUSER_WIDTH       = 1,
    C_USER_VALUE              = 1'b0,
    C_PROT_VALUE              = 3'b000,
    C_CACHE_VALUE             = 4'b0011,
    BUS_ADDR_WIDTH            = 32,
    BUS_DATA_WIDTH            = 32,
    NUM_WRITE_OUTSTANDING     = 2,
    MAX_WRITE_BURST_LENGTH    = 16
)(
    // system signal
    input  wire                             ACLK,
    input  wire                             ARESET,
    input  wire                             ACLK_EN,
    // write address channel
    output wire [C_M_AXI_ID_WIDTH-1:0]      out_BUS_AWID,
    output wire [2:0]                       out_BUS_AWSIZE,
    output wire [1:0]                       out_BUS_AWBURST,
    output wire [1:0]                       out_BUS_AWLOCK,
    output wire [3:0]                       out_BUS_AWCACHE,
    output wire [2:0]                       out_BUS_AWPROT,
    output wire [3:0]                       out_BUS_AWQOS,
    output wire [3:0]                       out_BUS_AWREGION,
    output wire [C_M_AXI_AWUSER_WIDTH-1:0]  out_BUS_AWUSER,
    output wire [BUS_ADDR_WIDTH-1:0]        out_BUS_AWADDR,
    output wire [7:0]                       out_BUS_AWLEN,
    output wire                             out_BUS_AWVALID,
    input  wire                             in_BUS_AWREADY,
    // write data channel
    output wire [C_M_AXI_ID_WIDTH-1:0]      out_BUS_WID,
    output wire [C_M_AXI_WUSER_WIDTH-1:0]   out_BUS_WUSER,
    output wire [BUS_DATA_WIDTH-1:0]        out_BUS_WDATA,
    output wire [BUS_DATA_WIDTH/8-1:0]      out_BUS_WSTRB,
    output wire                             out_BUS_WLAST,
    output wire                             out_BUS_WVALID,
    input  wire                             in_BUS_WREADY,
    // write response channel
    input  wire [C_M_AXI_ID_WIDTH-1:0]      in_BUS_BID,
    input  wire [1:0]                       in_BUS_BRESP,
    input  wire [C_M_AXI_BUSER_WIDTH-1:0]   in_BUS_BUSER,
    input  wire                             in_BUS_BVALID,
    output wire                             out_BUS_BREADY,
    // write request
    input  wire [BUS_ADDR_WIDTH-1:0]        in_HLS_AWADDR,
    input  wire [31:0]                      in_HLS_AWLEN,
    input  wire                             in_HLS_AWVALID,
    output wire                             out_HLS_AWREADY,

    input  wire [BUS_DATA_WIDTH-1:0]        in_HLS_WDATA,
    input  wire [BUS_DATA_WIDTH/8-1:0]      in_HLS_WSTRB,
    input  wire                             in_HLS_WVALID,
    output wire                             out_HLS_WREADY,
    output wire                             out_HLS_BVALID,
    input  wire                             in_HLS_BREADY);

//------------------------Parameter----------------------
    localparam
        BUS_DATA_BYTES  = BUS_DATA_WIDTH / 8,
        BUS_ADDR_ALIGN  = log2(BUS_DATA_BYTES),
        NUM_WRITE_WIDTH = log2(MAX_WRITE_BURST_LENGTH),
        BOUNDARY_BEATS  = {12-BUS_ADDR_ALIGN{1'b1}};

//------------------------Task and function--------------
    function integer calc_data_width;
        input integer x;
        integer y;
    begin
        y = 8;
        while (y < x) y = y * 2;
        calc_data_width = y;
    end
    endfunction

    function integer log2;
        input integer x;
        integer n, m;
    begin
        n = 0;
        m = 1;
        while (m < x) begin
            n = n + 1;
            m = m * 2;
        end
        log2 = n;
    end
    endfunction

//------------------------Local signal-------------------
    // AW channel
    wire                                wreq_valid;
    wire [BUS_ADDR_WIDTH - 1:0]         tmp_addr;
    wire [31:0]                         tmp_len;
    wire [7:0]                          awlen_tmp;
    wire [BUS_ADDR_WIDTH - 1:0]         awaddr_tmp;
    reg  [BUS_ADDR_WIDTH - 1:0]         start_addr;
    reg  [BUS_ADDR_WIDTH - 1:0]         end_addr;
    wire [BUS_ADDR_WIDTH - 1:0]         sect_addr;
    reg  [BUS_ADDR_WIDTH - 1:0]         sect_addr_buf;
    wire [11 - BUS_ADDR_ALIGN:0]        start_to_4k;
    wire [11 - BUS_ADDR_ALIGN:0]        sect_len;
    reg  [11 - BUS_ADDR_ALIGN:0]        sect_len_buf;
    reg  [11 - BUS_ADDR_ALIGN:0]        beat_len;
    wire                                aw2b_info;
    reg  [BUS_ADDR_WIDTH - 13:0]        sect_cnt;
    wire                                fifo_burst_w;
    wire                                fifo_resp_w;

    wire [BUS_ADDR_WIDTH - 1:0]         AWADDR_Dummy;
    wire [7:0]                          AWLEN_Dummy;
    reg                                 AWVALID_Dummy;
    wire                                AWREADY_Dummy;
    wire                                ready_for_sect;
    wire                                next_wreq;
    wire                                ready_for_wreq;
    reg                                 wreq_handling;
    wire                                first_sect;
    reg                                 last_sect_buf;
    wire                                last_sect;
    wire                                next_sect;
    // W channel
    wire                                next_data;
    wire                                data_valid;
    wire                                data_ready;
    reg  [BUS_DATA_WIDTH - 1:0]         data_buf;
    reg  [BUS_DATA_BYTES - 1:0]         strb_buf;
    wire                                ready_for_data;

    reg  [7:0]                          len_cnt;
    wire [7:0]                          burst_len;
    wire                                fifo_burst_ready;
    wire                                next_burst;
    wire                                burst_valid;
    reg                                 WVALID_Dummy;
    wire                                WREADY_Dummy;
    reg                                 WLAST_Dummy;
    //B channel
    wire                                next_resp;
    wire                                last_resp;
    wire                                fifo_resp_ready;
    wire                                need_wrsp;
    wire                                resp_valid;
    wire                                resp_ready;

//------------------------AW channel begin---------------
//------------------------Instantiation------------------
    kmeans_top_mem_m_axi_reg_slice #(
        .DATA_WIDTH     (BUS_ADDR_WIDTH + 32)
    ) rs_wreq (
        .clk            (ACLK),
        .reset          (ARESET),
        .s_data         ({in_HLS_AWLEN, in_HLS_AWADDR}),
        .s_valid        (in_HLS_AWVALID),
        .s_ready        (out_HLS_AWREADY),
        .m_data         ({tmp_len, tmp_addr}),
        .m_valid        (wreq_valid),
        .m_ready        (next_wreq));

//------------------------Body---------------------------
    assign ready_for_wreq = last_sect & next_sect | ~wreq_handling;
    assign next_wreq      = wreq_valid & ready_for_wreq;

    always @(posedge ACLK)
    begin
        if (ARESET) begin
            start_addr <= 0;
            end_addr   <= 0;
            beat_len   <= 0;
        end
        else if (ACLK_EN) begin
            if (next_wreq) begin
                start_addr <= tmp_addr;
                end_addr   <= tmp_addr + tmp_len;
                beat_len   <= (tmp_len[11:0] + tmp_addr[BUS_ADDR_ALIGN-1:0]) >> BUS_ADDR_ALIGN;
            end
        end
    end

    always @(posedge ACLK)
    begin
        if (ARESET)
            wreq_handling <= 1'b0;
        else if (ACLK_EN) begin
            if (wreq_valid && ~wreq_handling)
                wreq_handling <= 1'b1;
            else if (~wreq_valid && last_sect && next_sect)
                wreq_handling <= 1'b0;
        end
    end

    // 4k boundary
    assign first_sect = (sect_cnt == start_addr[BUS_ADDR_WIDTH-1:12]);
    assign last_sect  = (sect_cnt == end_addr[BUS_ADDR_WIDTH-1:12]);
    assign next_sect  = wreq_handling && ready_for_sect;

    assign sect_addr  = (first_sect)? start_addr : {sect_cnt, {12{1'b0}}};

    assign start_to_4k = BOUNDARY_BEATS - start_addr[11:BUS_ADDR_ALIGN];
    assign sect_len    = ( first_sect &&  last_sect)? beat_len :
                         ( first_sect && ~last_sect)? start_to_4k:
                         (~first_sect &&  last_sect)? end_addr[11:BUS_ADDR_ALIGN] :
                                                      BOUNDARY_BEATS;

    always @(posedge ACLK)
    begin
        if (ARESET)
            sect_cnt <= 0;
        else if (ACLK_EN) begin
            if (next_wreq)
                sect_cnt <= tmp_addr[BUS_ADDR_WIDTH-1:12];
            else if (next_sect)
                sect_cnt <= sect_cnt + 1;
        end
    end

    always @(posedge ACLK)
    begin
        if (ARESET) begin
            sect_addr_buf <= 0;
            sect_len_buf <= 0;
            last_sect_buf <= 1'b0;
        end
        else if (ACLK_EN) begin
            if (next_sect) begin
                sect_addr_buf <= sect_addr;
                sect_len_buf <= sect_len;
                last_sect_buf <= last_sect;
            end
        end
    end

    // burst converter
    assign out_BUS_AWID     = 0;
    assign out_BUS_AWSIZE   = BUS_ADDR_ALIGN;
    assign out_BUS_AWBURST  = 2'b01;
    assign out_BUS_AWLOCK   = 2'b00;
    assign out_BUS_AWCACHE  = C_CACHE_VALUE;
    assign out_BUS_AWPROT   = C_PROT_VALUE;
    assign out_BUS_AWUSER   = C_USER_VALUE;
    assign out_BUS_AWQOS    = 4'b0000;
    assign out_BUS_AWREGION = 4'b0000;

    generate
    if (BUS_DATA_BYTES >= 4096/MAX_WRITE_BURST_LENGTH) begin : must_one_burst
        assign AWADDR_Dummy   = {sect_addr_buf[BUS_ADDR_WIDTH - 1:BUS_ADDR_ALIGN], {BUS_ADDR_ALIGN{1'b0}}};
        assign AWLEN_Dummy    = sect_len_buf;

        assign ready_for_sect = ~(AWVALID_Dummy && ~AWREADY_Dummy) && fifo_burst_ready && fifo_resp_ready;

        always @(posedge ACLK)
        begin
            if (ARESET)
                AWVALID_Dummy <= 1'b0;
            else if (ACLK_EN) begin
                if (next_sect)
                    AWVALID_Dummy <= 1'b1;
                else if (~next_sect && AWREADY_Dummy)
                    AWVALID_Dummy <= 1'b0;
            end
        end

        assign fifo_resp_w = next_sect;
        assign aw2b_info   = last_sect;

        assign fifo_burst_w = next_sect;
        assign awaddr_tmp   = sect_addr[BUS_ADDR_WIDTH - 1:0];
        assign awlen_tmp    = sect_len;
    end
    else begin : could_multi_bursts
        reg  [BUS_ADDR_WIDTH - 1:0]                         awaddr_buf;
        reg  [7:0]                                          awlen_buf;
        reg  [11 - NUM_WRITE_WIDTH - BUS_ADDR_ALIGN : 0]    loop_cnt;
        reg                                                 sect_handling;
        wire                                                last_loop;
        wire                                                next_loop;
        wire                                                ready_for_loop;

        assign AWADDR_Dummy   = awaddr_buf;
        assign AWLEN_Dummy    = awlen_buf;

        assign last_loop      = (loop_cnt == sect_len_buf[11 - BUS_ADDR_ALIGN : NUM_WRITE_WIDTH]);
        assign next_loop      = sect_handling && ready_for_loop;
        assign ready_for_loop = ~(AWVALID_Dummy && ~AWREADY_Dummy) && fifo_burst_ready && fifo_resp_ready;
        assign ready_for_sect = ~(sect_handling && ~(last_loop && next_loop));

        always @(posedge ACLK)
        begin
            if (ARESET)
                sect_handling <= 1'b0;
            else if (ACLK_EN) begin
                if (wreq_handling && ~sect_handling)
                    sect_handling <= 1'b1;
                else if (~wreq_handling && last_loop && next_loop)
                    sect_handling <= 1'b0;
            end
        end

        always @(posedge ACLK)
        begin
            if (ARESET)
                loop_cnt <= 0;
            else if (ACLK_EN) begin
                if (next_sect)
                    loop_cnt <= 0;
                else if (next_loop)
                    loop_cnt <= loop_cnt + 1;
            end
        end

        assign awaddr_tmp = (loop_cnt == 0)? sect_addr_buf[BUS_ADDR_WIDTH - 1:0] : (awaddr_buf + ((awlen_buf + 1) << BUS_ADDR_ALIGN));
        assign awlen_tmp  = (NUM_WRITE_WIDTH == 0)? 0 :
                    (last_loop)? sect_len_buf[NUM_WRITE_WIDTH - 1:0] : { NUM_WRITE_WIDTH{1'b1} };
        always @(posedge ACLK)
        begin
            if (ARESET) begin
                awaddr_buf <= 0;
                awlen_buf <= 0;
            end
            else if (ACLK_EN) begin
                if (next_loop) begin
                    awaddr_buf <= {awaddr_tmp[BUS_ADDR_WIDTH - 1:BUS_ADDR_ALIGN], {BUS_ADDR_ALIGN{1'b0}}};
                    awlen_buf <= awlen_tmp;
                end
            end
        end

        always @(posedge ACLK)
        begin
            if (ARESET)
                AWVALID_Dummy <= 1'b0;
            else if (ACLK_EN) begin
                if (next_loop)
                    AWVALID_Dummy <= 1'b1;
                else if (~next_loop && AWREADY_Dummy)
                    AWVALID_Dummy <= 1'b0;
            end
        end

        assign fifo_resp_w = next_loop;
        assign fifo_burst_w = next_loop;
        assign aw2b_info = last_loop && last_sect_buf;
    end
    endgenerate
//------------------------AW channel end-----------------

//------------------------W channel begin----------------
//------------------------Instantiation------------------

    kmeans_top_mem_m_axi_fifo #(
        .DATA_WIDTH     (8),
        .ADDR_WIDTH     (log2(NUM_WRITE_OUTSTANDING)),
        .DEPTH          (NUM_WRITE_OUTSTANDING)
    ) fifo_burst (
        .clk            (ACLK),
        .reset          (ARESET),
        .clk_en         (ACLK_EN),
        .if_full_n      (fifo_burst_ready),
        .if_write       (fifo_burst_w),
        .if_din         (awlen_tmp),
        .if_empty_n     (burst_valid),
        .if_read        (next_burst),
        .if_dout        (burst_len),
        .if_num_data_valid());

//------------------------Body---------------------------

    assign out_BUS_WUSER    = C_USER_VALUE;
    assign out_BUS_WID      = 0;
    assign out_HLS_WREADY   = data_ready;

    assign data_valid       = in_HLS_WVALID;
    assign data_ready       = burst_valid && ready_for_data;
    assign next_data        = data_ready && data_valid;
    assign next_burst       = (len_cnt == burst_len) && next_data;
    assign ready_for_data   = ~WVALID_Dummy || WREADY_Dummy;

    always @(posedge ACLK)
    begin
        if (ARESET) begin
            strb_buf <= 0;
            data_buf <= 0;
        end
        if (ACLK_EN) begin
            if (next_data) begin
                data_buf <= in_HLS_WDATA;
                strb_buf <= in_HLS_WSTRB;
            end
        end
    end

    always @(posedge ACLK)
    begin
        if (ARESET)
            WVALID_Dummy <= 1'b0;
        else if (ACLK_EN) begin
            if (next_data)
                WVALID_Dummy <= 1'b1;
            else if (ready_for_data)
                WVALID_Dummy <= 1'b0;
        end
    end

    always @(posedge ACLK)
    begin
        if (ARESET)
            WLAST_Dummy <= 0;
        else if (ACLK_EN) begin
            if (next_burst)
                WLAST_Dummy <= 1;
            else if (ready_for_data)
                WLAST_Dummy <= 0;
        end
    end

    always @(posedge ACLK)
    begin
        if (ARESET)
            len_cnt <= 0;
        else if (ACLK_EN) begin
            if (next_burst)
                len_cnt <= 0;
            else if (next_data)
                len_cnt <= len_cnt + 1;
        end
    end
//------------------------W channel end------------------

    // Write throttling unit
    kmeans_top_mem_m_axi_throttle #(
        .CONSERVATIVE(CONSERVATIVE),
        .USED_FIX(0),
        .ADDR_WIDTH(BUS_ADDR_WIDTH),
        .DATA_WIDTH(BUS_DATA_WIDTH),
        .DEPTH(MAX_WRITE_BURST_LENGTH),
        .MAXREQS(NUM_WRITE_OUTSTANDING),
        .AVERAGE_MODE(0)
    ) wreq_throttle (
        .clk(ACLK),
        .reset(ARESET),
        .clk_en(ACLK_EN),
        // internal 
        .in_TOP_AWADDR(AWADDR_Dummy),
        .in_TOP_AWLEN(AWLEN_Dummy),
        .in_TOP_AWVALID(AWVALID_Dummy),
        .out_TOP_AWREADY(AWREADY_Dummy),

        .in_TOP_WDATA(data_buf),
        .in_TOP_WSTRB(strb_buf),
        .in_TOP_WLAST(WLAST_Dummy),
        .in_TOP_WVALID(WVALID_Dummy),
        .out_TOP_WREADY(WREADY_Dummy),

        // AXI BUS
        .out_BUS_AWADDR(out_BUS_AWADDR),
        .out_BUS_AWLEN(out_BUS_AWLEN),
        .out_BUS_AWVALID(out_BUS_AWVALID),
        .in_BUS_AWREADY(in_BUS_AWREADY),

        .out_BUS_WDATA(out_BUS_WDATA),
        .out_BUS_WSTRB(out_BUS_WSTRB),
        .out_BUS_WLAST(out_BUS_WLAST),
        .out_BUS_WVALID(out_BUS_WVALID),
        .in_BUS_WREADY(in_BUS_WREADY)
    );
    
//------------------------B channel begin----------------
//------------------------Instantiation------------------
    kmeans_top_mem_m_axi_reg_slice #(
        .DATA_WIDTH     (1)
    ) rs_resp (
        .clk            (ACLK),
        .reset          (ARESET),
        .s_data         (1'b1),
        .s_valid        (in_BUS_BVALID),
        .s_ready        (out_BUS_BREADY),
        .m_data         (),
        .m_valid        (resp_valid),
        .m_ready        (resp_ready));

    kmeans_top_mem_m_axi_fifo #(
        .DATA_WIDTH     (1),
        .ADDR_WIDTH     (log2(NUM_WRITE_OUTSTANDING)),
        .DEPTH          (NUM_WRITE_OUTSTANDING)
    ) fifo_resp (
        .clk            (ACLK),
        .reset          (ARESET),
        .clk_en         (ACLK_EN),
        .if_full_n      (fifo_resp_ready),
        .if_write       (fifo_resp_w),
        .if_din         (aw2b_info),
        .if_empty_n     (need_wrsp),
        .if_read        (next_resp),
        .if_dout        (last_resp),
        .if_num_data_valid());
//------------------------Body---------------------------

    assign resp_ready = need_wrsp && (in_HLS_BREADY || (last_resp === 1'b0));
    assign next_resp  = resp_ready && resp_valid;

    assign out_HLS_BVALID = resp_valid && (last_resp === 1'b1 ) ;

//------------------------B channel end------------------
endmodule

module kmeans_top_mem_m_axi_throttle
#(parameter
    CONSERVATIVE   = 0,
    USED_FIX       = 0,
    FIX_VALUE      = 4,
    ADDR_WIDTH     = 32,
    DATA_WIDTH     = 32,
    DEPTH          = 16,
    MAXREQS        = 16,
    AVERAGE_MODE   = 0 
)(
    input  wire                      clk,
    input  wire                      reset,
    input  wire                      clk_en,

    input  wire [ADDR_WIDTH-1:0]     in_TOP_AWADDR,
    input  wire [7:0]                in_TOP_AWLEN,
    input  wire                      in_TOP_AWVALID,
    output wire                      out_TOP_AWREADY,
    input  wire [DATA_WIDTH-1:0]     in_TOP_WDATA,
    input  wire [DATA_WIDTH/8-1:0]   in_TOP_WSTRB,
    input  wire                      in_TOP_WLAST,
    input  wire                      in_TOP_WVALID,
    output wire                      out_TOP_WREADY,

    output wire [ADDR_WIDTH-1:0]     out_BUS_AWADDR,
    output wire [7:0]                out_BUS_AWLEN,
    output wire                      out_BUS_AWVALID,
    input  wire                      in_BUS_AWREADY,
    output wire [DATA_WIDTH-1:0]     out_BUS_WDATA,
    output wire [DATA_WIDTH/8-1:0]   out_BUS_WSTRB,
    output wire                      out_BUS_WLAST,
    output wire                      out_BUS_WVALID,
    input  wire                      in_BUS_WREADY);

    function integer log2;
        input integer x;
        integer n, m;
    begin
        n = 0;
        m = 1;
        while (m < x) begin
            n = n + 1;
            m = m * 2;
        end
        log2 = n;
    end
    endfunction
// aggressive mode
    generate
    if (CONSERVATIVE == 0) begin
        localparam threshold = (USED_FIX)? FIX_VALUE-1 : 0;

        wire                req_en;
        wire                handshake;
        wire  [7:0]         load_init;
        reg   [8:0]         throttl_cnt;

        // AW Channel
        assign out_BUS_AWADDR = in_TOP_AWADDR;
        assign out_BUS_AWLEN  = in_TOP_AWLEN;

        // W Channel
        assign out_BUS_WDATA  = in_TOP_WDATA;
        assign out_BUS_WSTRB  = in_TOP_WSTRB;
        assign out_BUS_WLAST  = in_TOP_WLAST;
        assign out_BUS_WVALID = in_TOP_WVALID & (throttl_cnt > 0);
        assign out_TOP_WREADY = in_BUS_WREADY & (throttl_cnt > 0);

        if (USED_FIX) begin
            assign load_init = FIX_VALUE-1;
            assign handshake = 1'b1;
        end else if (AVERAGE_MODE) begin
            assign load_init = in_TOP_AWLEN;
            assign handshake = 1'b1;
        end else begin
            assign load_init = in_TOP_AWLEN;
            assign handshake = out_BUS_WVALID & in_BUS_WREADY;
        end

        assign out_BUS_AWVALID = in_TOP_AWVALID & req_en;
        assign out_TOP_AWREADY = in_BUS_AWREADY & req_en;
        assign req_en = (throttl_cnt == 0) | (throttl_cnt == 1 & handshake);

        always @(posedge clk)
        begin
            if (reset)
                throttl_cnt <= 0;
            else if (clk_en) begin
                if (in_TOP_AWLEN >= threshold && req_en && in_TOP_AWVALID && in_BUS_AWREADY)
                    throttl_cnt <= load_init + 1'b1; //load
                else if (throttl_cnt > 0 && handshake)
                    throttl_cnt <= throttl_cnt - 1'b1;
            end
        end

    end
// conservative mode
    else begin
        localparam CNT_WIDTH = ((DEPTH < 4)? 2 : log2(DEPTH)) + 1;

        // Instantiation for reg slice for AW channel
        wire                        rs_req_ready;
        wire                        rs_req_valid;
        wire [ADDR_WIDTH + 7 : 0]   rs_req_in;
        wire [ADDR_WIDTH + 7 : 0]   rs_req_out;

        kmeans_top_mem_m_axi_reg_slice #(
            .DATA_WIDTH     (ADDR_WIDTH + 8)
        ) rs_req (
            .clk            (clk),
            .reset          (reset),
            .s_data         (rs_req_in),
            .s_valid        (rs_req_valid),
            .s_ready        (rs_req_ready),
            .m_data         (rs_req_out),
            .m_valid        (out_BUS_AWVALID),
            .m_ready        (in_BUS_AWREADY));

        wire  [DATA_WIDTH + DATA_WIDTH/8 : 0]   data_in;
        wire  [DATA_WIDTH + DATA_WIDTH/8 : 0]   data_out;
        wire  [ADDR_WIDTH + 7 : 0]              req_in;
        reg                                     req_en;
        wire                                    data_en;
        wire                                    fifo_valid;
        wire                                    read_fifo;
        wire                                    req_fifo_valid;
        wire                                    read_req;
        wire                                    data_push;
        wire                                    data_pop;
        reg                                     flying_req;
        reg   [CNT_WIDTH-1 : 0]                 last_cnt;

        //AW Channel
        assign req_in   = {in_TOP_AWLEN, in_TOP_AWADDR};
        assign out_BUS_AWADDR = rs_req_out[ADDR_WIDTH-1 : 0];
        assign out_BUS_AWLEN  = rs_req_out[ADDR_WIDTH+7 : ADDR_WIDTH];
        assign rs_req_valid = req_fifo_valid & req_en;

        assign read_req      = rs_req_ready & req_en;

        always @(*)
        begin
            if (~flying_req & data_en)
                req_en <= 1;
            else if (flying_req & (out_BUS_WLAST & data_pop) & (last_cnt[CNT_WIDTH-1:1] != 0))
                req_en <= 1;
            else
                req_en <= 0;
        end

        always @(posedge clk)
        begin
            if (reset)
                flying_req <= 0;
            else if (clk_en) begin
                if (rs_req_valid & rs_req_ready)
                    flying_req <= 1;
                else if (out_BUS_WLAST & data_pop)
                    flying_req <= 0;
            end
        end

        kmeans_top_mem_m_axi_fifo #(
            .DATA_WIDTH     (ADDR_WIDTH + 8),
            .ADDR_WIDTH     (log2(MAXREQS)),
            .DEPTH          (MAXREQS)
        ) req_fifo (
            .clk            (clk),
            .reset          (reset),
            .clk_en         (clk_en),
            .if_full_n      (out_TOP_AWREADY),
            .if_write       (in_TOP_AWVALID),
            .if_din         (req_in),
            .if_empty_n     (req_fifo_valid),
            .if_read        (read_req),
            .if_dout        (rs_req_in),
            .if_num_data_valid());

        //W Channel
        assign data_in  = {in_TOP_WLAST, in_TOP_WSTRB, in_TOP_WDATA};
        assign out_BUS_WDATA = data_out[DATA_WIDTH-1 : 0];
        assign out_BUS_WSTRB = data_out[DATA_WIDTH+DATA_WIDTH/8-1 : DATA_WIDTH];
        assign out_BUS_WLAST = data_out[DATA_WIDTH+DATA_WIDTH/8];
        assign out_BUS_WVALID = fifo_valid & data_en & flying_req;

        assign data_en   = last_cnt != 0;
        assign data_push = in_TOP_WVALID & out_TOP_WREADY;
        assign data_pop  = fifo_valid & read_fifo;
        assign read_fifo = in_BUS_WREADY & data_en & flying_req;

        always @(posedge clk)
        begin
            if (reset)
                last_cnt <= 0;
            else if (clk_en) begin
                if ((in_TOP_WLAST & data_push) && ~(out_BUS_WLAST & data_pop))
                    last_cnt <= last_cnt + 1;
                else if (~(in_TOP_WLAST & data_push) && (out_BUS_WLAST & data_pop))
                    last_cnt <= last_cnt - 1;
            end
        end
            
        kmeans_top_mem_m_axi_fifo #(
            .DATA_WIDTH     (DATA_WIDTH + DATA_WIDTH/8 + 1),
            .ADDR_WIDTH     (log2(DEPTH)),
            .DEPTH          (DEPTH)
        ) data_fifo (
            .clk            (clk),
            .reset          (reset),
            .clk_en         (clk_en),
            .if_full_n      (out_TOP_WREADY),
            .if_write       (in_TOP_WVALID),
            .if_din         (data_in),
            .if_empty_n     (fifo_valid),
            .if_read        (read_fifo),
            .if_dout        (data_out),
            .if_num_data_valid());

        end
    endgenerate

endmodule


module kmeans_top_mem_m_axi_reg_slice
#(parameter
    DATA_WIDTH = 8
) (
    // system signals
    input  wire                  clk,
    input  wire                  reset,
    // slave side
    input  wire [DATA_WIDTH-1:0] s_data,
    input  wire                  s_valid,
    output wire                  s_ready,
    // master side
    output wire [DATA_WIDTH-1:0] m_data,
    output wire                  m_valid,
    input  wire                  m_ready);
    //------------------------Parameter----------------------
    // state
    localparam [1:0]
        ZERO = 2'b10,
        ONE  = 2'b11,
        TWO  = 2'b01;
    //------------------------Local signal-------------------
    reg  [DATA_WIDTH-1:0] data_p1;
    reg  [DATA_WIDTH-1:0] data_p2;
    wire         load_p1;
    wire         load_p2;
    wire         load_p1_from_p2;
    reg          s_ready_t;
    reg  [1:0]   state;
    reg  [1:0]   next;
    //------------------------Body---------------------------
    assign s_ready = s_ready_t;
    assign m_data  = data_p1;
    assign m_valid = state[0];

    assign load_p1 = (state == ZERO && s_valid) ||
                    (state == ONE && s_valid && m_ready) ||
                    (state == TWO && m_ready);
    assign load_p2 = s_valid & s_ready;
    assign load_p1_from_p2 = (state == TWO);

    // data_p1
    always @(posedge clk) begin
        if (load_p1) begin
            if (load_p1_from_p2)
                data_p1 <= data_p2;
            else
                data_p1 <= s_data;
        end
    end

    // data_p2
    always @(posedge clk) begin
        if (load_p2) data_p2 <= s_data;
    end

    // s_ready_t
    always @(posedge clk) begin
        if (reset)
            s_ready_t <= 1'b0;
        else if (state == ZERO)
            s_ready_t <= 1'b1;
        else if (state == ONE && next == TWO)
            s_ready_t <= 1'b0;
        else if (state == TWO && next == ONE)
            s_ready_t <= 1'b1;
    end

    // state
    always @(posedge clk) begin
        if (reset)
            state <= ZERO;
        else
            state <= next;
    end

    // next
    always @(*) begin
        case (state)
            ZERO:
                if (s_valid & s_ready)
                    next = ONE;
                else
                    next = ZERO;
            ONE:
                if (~s_valid & m_ready)
                    next = ZERO;
                else if (s_valid & ~m_ready)
                    next = TWO;
                else
                    next = ONE;
            TWO:
                if (m_ready)
                    next = ONE;
                else
                    next = TWO;
            default:
                next = ZERO;
        endcase
    end
endmodule

module kmeans_top_mem_m_axi_fifo
#(parameter
    MEM_STYLE   = "shiftreg",
    DATA_WIDTH = 32,
    ADDR_WIDTH = 5,
    DEPTH      = 32
) (
    // system signal
    input  wire                  clk,
    input  wire                  reset,
    input  wire                  clk_en,

    // write
    output wire                  if_full_n,
    input  wire                  if_write,
    input  wire [DATA_WIDTH-1:0] if_din,

    // read
    output wire                  if_empty_n,
    input  wire                  if_read,
    output wire [DATA_WIDTH-1:0] if_dout,
    output wire [ADDR_WIDTH:0]   if_num_data_valid);

//------------------------Local signal-------------------

    wire                  push;
    wire                  pop;
    reg                   full_n = 1'b1;
    reg                   empty_n = 1'b0;
    reg                   dout_vld = 1'b0;
    reg  [ADDR_WIDTH:0]   mOutPtr = 1'b0;

//------------------------Instantiation------------------
    generate 
    if ((MEM_STYLE == "shiftreg") || (DEPTH == 1)) begin
        reg  [ADDR_WIDTH-1:0] raddr = 1'b0;

        kmeans_top_mem_m_axi_srl
        #(  .DATA_WIDTH     (DATA_WIDTH),
            .ADDR_WIDTH     (ADDR_WIDTH),
            .DEPTH          (DEPTH))
        U_fifo_srl(
            .clk            (clk),
            .reset          (reset),
            .clk_en         (clk_en),
            .we             (push),
            .din            (if_din),
            .raddr          (raddr),
            .re             (pop),
            .dout           (if_dout)
        );

        // raddr
        always @(posedge clk) begin
            if (reset == 1'b1)
                raddr <= 1'b0;
            else if (clk_en) begin
                if (push & ~pop & empty_n)
                    raddr <= raddr + 1'b1;
                else if (~push & pop && raddr != 0)
                    raddr <= raddr - 1'b1;
            end
        end

    end else begin
        reg  [ADDR_WIDTH-1:0] waddr = 1'b0;
        reg  [ADDR_WIDTH-1:0] raddr = 1'b0;
        wire [ADDR_WIDTH-1:0] wnext;
        wire [ADDR_WIDTH-1:0] rnext;

        kmeans_top_mem_m_axi_mem
        #(  .MEM_STYLE      (MEM_STYLE),
            .DATA_WIDTH     (DATA_WIDTH),
            .ADDR_WIDTH     (ADDR_WIDTH),
            .DEPTH          (DEPTH))
        U_fifo_mem(
            .clk            (clk),
            .reset          (reset),
            .clk_en         (clk_en),
            .we             (push),
            .waddr          (waddr),
            .din            (if_din),
            .raddr          (rnext),
            .re             (pop),
            .dout           (if_dout)
        );

        assign wnext =  !push                ? waddr :
                        (waddr == DEPTH - 2) ? 1'b0  :
                        waddr + 1'b1;
        assign rnext =  !pop                 ? raddr :
                        (raddr == DEPTH - 2) ? 1'b0  :
                        raddr + 1'b1;

        // waddr
        always @(posedge clk) begin
            if (reset == 1'b1)
                waddr <= 1'b0;
            else if (clk_en)
                waddr <= wnext;
        end

        // raddr
        always @(posedge clk) begin
            if (reset == 1'b1)
                raddr <= 1'b0;
            else if (clk_en)
                raddr <= rnext;
        end
    end
    endgenerate

//------------------------Body---------------------------
    assign if_num_data_valid = dout_vld ? mOutPtr + 1'b1 : 'b0;

    generate if (DEPTH == 1) begin
        assign if_full_n  = !dout_vld;
        assign if_empty_n = dout_vld;
        assign push = !dout_vld & if_write;
        assign pop  = !dout_vld & if_write;
    
    end else begin

        assign if_full_n  = full_n;
        assign if_empty_n = dout_vld;
        assign push = full_n & if_write;
        assign pop  = empty_n & (if_read | ~dout_vld);

        // mOutPtr
        always @(posedge clk) begin
            if (reset == 1'b1)
                mOutPtr <= 'b0;
            else if (clk_en)
                if (push & ~pop)
                    mOutPtr <= mOutPtr + 1'b1;
                else if (~push & pop)
                    mOutPtr <= mOutPtr - 1'b1;
        end

        // full_n
        always @(posedge clk) begin
            if (reset == 1'b1)
                full_n <= 1'b1;
            else if (clk_en)
                if (push & ~pop)
                    full_n <= (mOutPtr != DEPTH - 2);
                else if (~push & pop)
                    full_n <= 1'b1;
        end

        // empty_n
        always @(posedge clk)
        begin
            if (reset)
                empty_n <= 1'b0;
            else if (clk_en) begin
                if (push & ~pop)
                    empty_n <= 1'b1;
                else if (~push & pop)
                    empty_n <= (mOutPtr != 1'b1);
            end
        end
    end
    endgenerate

    // dout_vld
    always @(posedge clk) begin
        if (reset == 1'b1)
            dout_vld <= 1'b0;
        else if (clk_en)
            if (pop)
                dout_vld <= 1'b1;
            else if (if_read)
                dout_vld <= 1'b0;
    end

endmodule

module kmeans_top_mem_m_axi_srl
#(parameter
        DATA_WIDTH  = 32,
        ADDR_WIDTH  = 6,
        DEPTH       = 63
    )(
        input  wire                  clk,
        input  wire                  reset,
        input  wire                  clk_en,
        input  wire                  we,
        input  wire [DATA_WIDTH-1:0] din,
        input  wire [ADDR_WIDTH-1:0] raddr,
        input  wire                  re,
        output reg  [DATA_WIDTH-1:0] dout
    );

    generate
    if (DEPTH > 1) begin
        reg  [DATA_WIDTH-1:0] mem[0:DEPTH-2];

        integer i;
        always @(posedge clk)
        begin
            if (clk_en & we) begin
                for (i = 0; i < DEPTH - 2; i = i + 1) begin
                    mem[i+1] <= mem[i];
                end
                mem[0] <= din;
            end
        end

        always @(posedge clk)
        begin
            if (reset)
                dout <= 0;
            else if (clk_en & re) begin
                dout <= mem[raddr];
            end
        end
    end
    else begin
        always @(posedge clk)
        begin
            if (reset)
                dout <= 0;
            else if (clk_en & we) begin
                dout <= din;
            end
        end
    end
    endgenerate

endmodule

module kmeans_top_mem_m_axi_mem
#(parameter
    MEM_STYLE   = "auto",
    DATA_WIDTH  = 32,
    ADDR_WIDTH  = 6,
    DEPTH       = 63
)(
    input  wire                  clk,
    input  wire                  reset,
    input  wire                  clk_en,
    input  wire                  we,
    input  wire [ADDR_WIDTH-1:0] waddr,
    input  wire [DATA_WIDTH-1:0] din,
    input  wire [ADDR_WIDTH-1:0] raddr,
    input  wire                  re,
    output reg  [DATA_WIDTH-1:0] dout);

    (* ram_style = MEM_STYLE, rw_addr_collision = "yes" *)
    reg  [DATA_WIDTH-1:0] mem[0:DEPTH-2];
    reg  [ADDR_WIDTH-1:0] raddr_reg;

    //write to ram
    always @(posedge clk) begin
        if (clk_en & we)
            mem[waddr] <= din;
    end

    //buffer the raddr
    always @(posedge clk) begin
        if (clk_en)
            raddr_reg <= raddr;
    end

    //read from ram
    always @(posedge clk) begin
        if (reset)
            dout <= 0;
        else if (clk_en & re)
            dout <= mem[raddr_reg];
    end
endmodule


// Content from kmeans_top_kmeans_Pipeline_2.v
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2022.2 (64-bit)
// Version: 2022.2
// Copyright (C) Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module kmeans_top_kmeans_Pipeline_2 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        cluster_cardinality_next_address0,
        cluster_cardinality_next_ce0,
        cluster_cardinality_next_we0,
        cluster_cardinality_next_d0,
        p_cast3_cast
);

parameter    ap_ST_fsm_pp0_stage0 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
output  [7:0] cluster_cardinality_next_address0;
output   cluster_cardinality_next_ce0;
output   cluster_cardinality_next_we0;
output  [15:0] cluster_cardinality_next_d0;
input  [33:0] p_cast3_cast;

reg ap_idle;
reg cluster_cardinality_next_ce0;
reg cluster_cardinality_next_we0;

(* fsm_encoding = "none" *) reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_enable_reg_pp0_iter0;
reg    ap_enable_reg_pp0_iter1;
reg    ap_idle_pp0;
wire    ap_block_state1_pp0_stage0_iter0;
wire    ap_block_state2_pp0_stage0_iter1;
wire    ap_block_pp0_stage0_subdone;
wire   [0:0] empty_74_fu_69_p2;
reg    ap_condition_exit_pp0_iter1_stage0;
wire    ap_loop_exit_ready;
reg    ap_ready_int;
wire   [63:0] p_cast3_cast_cast_cast_fu_50_p1;
reg   [63:0] p_cast3_cast_cast_cast_reg_86;
wire    ap_block_pp0_stage0_11001;
wire    ap_block_pp0_stage0;
reg   [63:0] empty_fu_22;
wire   [63:0] empty_73_fu_63_p2;
wire    ap_loop_init;
wire  signed [62:0] p_cast3_cast_cast_fu_46_p1;
reg    ap_done_reg;
wire    ap_continue_int;
reg    ap_done_int;
reg   [0:0] ap_NS_fsm;
wire    ap_enable_pp0;
wire    ap_start_int;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_CS_fsm = 1'd1;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_done_reg = 1'b0;
end

kmeans_top_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(ap_start),
    .ap_ready(ap_ready),
    .ap_done(ap_done),
    .ap_start_int(ap_start_int),
    .ap_loop_init(ap_loop_init),
    .ap_ready_int(ap_ready_int),
    .ap_loop_exit_ready(ap_condition_exit_pp0_iter1_stage0),
    .ap_loop_exit_done(ap_done_int),
    .ap_continue_int(ap_continue_int),
    .ap_done_int(ap_done_int)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue_int == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((ap_loop_exit_ready == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b1 == ap_condition_exit_pp0_iter1_stage0)) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_enable_reg_pp0_iter1 <= ap_start_int;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        if ((ap_loop_init == 1'b1)) begin
            empty_fu_22 <= 64'd0;
        end else if (((empty_74_fu_69_p2 == 1'd1) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
            empty_fu_22 <= empty_73_fu_63_p2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        p_cast3_cast_cast_cast_reg_86[62 : 0] <= p_cast3_cast_cast_cast_fu_50_p1[62 : 0];
    end
end

always @ (*) begin
    if (((empty_74_fu_69_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_condition_exit_pp0_iter1_stage0 = 1'b1;
    end else begin
        ap_condition_exit_pp0_iter1_stage0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_loop_exit_ready == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_done_int = 1'b1;
    end else begin
        ap_done_int = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_idle_pp0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_start_int == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_ready_int = 1'b1;
    end else begin
        ap_ready_int = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        cluster_cardinality_next_ce0 = 1'b1;
    end else begin
        cluster_cardinality_next_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        cluster_cardinality_next_we0 = 1'b1;
    end else begin
        cluster_cardinality_next_we0 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_pp0_stage0 : begin
            ap_NS_fsm = ap_ST_fsm_pp0_stage0;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

assign ap_block_state1_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_enable_reg_pp0_iter0 = ap_start_int;

assign ap_loop_exit_ready = ap_condition_exit_pp0_iter1_stage0;

assign cluster_cardinality_next_address0 = empty_fu_22;

assign cluster_cardinality_next_d0 = 16'd0;

assign empty_73_fu_63_p2 = (empty_fu_22 + 64'd1);

assign empty_74_fu_69_p2 = ((empty_73_fu_63_p2 < p_cast3_cast_cast_cast_reg_86) ? 1'b1 : 1'b0);

assign p_cast3_cast_cast_cast_fu_50_p1 = $unsigned(p_cast3_cast_cast_fu_46_p1);

assign p_cast3_cast_cast_fu_46_p1 = $signed(p_cast3_cast);

always @ (posedge ap_clk) begin
    p_cast3_cast_cast_cast_reg_86[63] <= 1'b0;
end

endmodule //kmeans_top_kmeans_Pipeline_2


// Content from kmeans_top_kmeans_top_Pipeline_1.v
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2022.2 (64-bit)
// Version: 2022.2
// Copyright (C) Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module kmeans_top_kmeans_top_Pipeline_1 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        m_axi_mem_AWVALID,
        m_axi_mem_AWREADY,
        m_axi_mem_AWADDR,
        m_axi_mem_AWID,
        m_axi_mem_AWLEN,
        m_axi_mem_AWSIZE,
        m_axi_mem_AWBURST,
        m_axi_mem_AWLOCK,
        m_axi_mem_AWCACHE,
        m_axi_mem_AWPROT,
        m_axi_mem_AWQOS,
        m_axi_mem_AWREGION,
        m_axi_mem_AWUSER,
        m_axi_mem_WVALID,
        m_axi_mem_WREADY,
        m_axi_mem_WDATA,
        m_axi_mem_WSTRB,
        m_axi_mem_WLAST,
        m_axi_mem_WID,
        m_axi_mem_WUSER,
        m_axi_mem_ARVALID,
        m_axi_mem_ARREADY,
        m_axi_mem_ARADDR,
        m_axi_mem_ARID,
        m_axi_mem_ARLEN,
        m_axi_mem_ARSIZE,
        m_axi_mem_ARBURST,
        m_axi_mem_ARLOCK,
        m_axi_mem_ARCACHE,
        m_axi_mem_ARPROT,
        m_axi_mem_ARQOS,
        m_axi_mem_ARREGION,
        m_axi_mem_ARUSER,
        m_axi_mem_RVALID,
        m_axi_mem_RREADY,
        m_axi_mem_RDATA,
        m_axi_mem_RLAST,
        m_axi_mem_RID,
        m_axi_mem_RFIFONUM,
        m_axi_mem_RUSER,
        m_axi_mem_RRESP,
        m_axi_mem_BVALID,
        m_axi_mem_BREADY,
        m_axi_mem_BRESP,
        m_axi_mem_BID,
        m_axi_mem_BUSER,
        p_cast_cast,
        node_x_coords_address1,
        node_x_coords_ce1,
        node_x_coords_we1,
        node_x_coords_d1,
        sext_ln182
);

parameter    ap_ST_fsm_pp0_stage0 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
output   m_axi_mem_AWVALID;
input   m_axi_mem_AWREADY;
output  [63:0] m_axi_mem_AWADDR;
output  [0:0] m_axi_mem_AWID;
output  [31:0] m_axi_mem_AWLEN;
output  [2:0] m_axi_mem_AWSIZE;
output  [1:0] m_axi_mem_AWBURST;
output  [1:0] m_axi_mem_AWLOCK;
output  [3:0] m_axi_mem_AWCACHE;
output  [2:0] m_axi_mem_AWPROT;
output  [3:0] m_axi_mem_AWQOS;
output  [3:0] m_axi_mem_AWREGION;
output  [0:0] m_axi_mem_AWUSER;
output   m_axi_mem_WVALID;
input   m_axi_mem_WREADY;
output  [63:0] m_axi_mem_WDATA;
output  [7:0] m_axi_mem_WSTRB;
output   m_axi_mem_WLAST;
output  [0:0] m_axi_mem_WID;
output  [0:0] m_axi_mem_WUSER;
output   m_axi_mem_ARVALID;
input   m_axi_mem_ARREADY;
output  [63:0] m_axi_mem_ARADDR;
output  [0:0] m_axi_mem_ARID;
output  [31:0] m_axi_mem_ARLEN;
output  [2:0] m_axi_mem_ARSIZE;
output  [1:0] m_axi_mem_ARBURST;
output  [1:0] m_axi_mem_ARLOCK;
output  [3:0] m_axi_mem_ARCACHE;
output  [2:0] m_axi_mem_ARPROT;
output  [3:0] m_axi_mem_ARQOS;
output  [3:0] m_axi_mem_ARREGION;
output  [0:0] m_axi_mem_ARUSER;
input   m_axi_mem_RVALID;
output   m_axi_mem_RREADY;
input  [63:0] m_axi_mem_RDATA;
input   m_axi_mem_RLAST;
input  [0:0] m_axi_mem_RID;
input  [8:0] m_axi_mem_RFIFONUM;
input  [0:0] m_axi_mem_RUSER;
input  [1:0] m_axi_mem_RRESP;
input   m_axi_mem_BVALID;
output   m_axi_mem_BREADY;
input  [1:0] m_axi_mem_BRESP;
input  [0:0] m_axi_mem_BID;
input  [0:0] m_axi_mem_BUSER;
input  [60:0] p_cast_cast;
output  [12:0] node_x_coords_address1;
output   node_x_coords_ce1;
output   node_x_coords_we1;
output  [63:0] node_x_coords_d1;
input  [31:0] sext_ln182;

reg ap_idle;
reg m_axi_mem_RREADY;
reg node_x_coords_ce1;
reg node_x_coords_we1;

(* fsm_encoding = "none" *) reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_enable_reg_pp0_iter0;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter2;
reg    ap_idle_pp0;
wire    ap_block_state1_pp0_stage0_iter0;
reg    ap_block_state2_pp0_stage0_iter1;
wire    ap_block_state3_pp0_stage0_iter2;
reg    ap_block_pp0_stage0_subdone;
wire   [0:0] exitcond85_fu_126_p2;
reg    ap_condition_exit_pp0_iter1_stage0;
wire    ap_loop_exit_ready;
reg    ap_ready_int;
reg    mem_blk_n_R;
wire    ap_block_pp0_stage0;
wire  signed [60:0] sext_ln182_cast_fu_98_p1;
reg  signed [60:0] sext_ln182_cast_reg_147;
reg    ap_block_pp0_stage0_11001;
reg   [60:0] loop_index69_load_reg_157;
reg   [63:0] mem_addr_read_reg_162;
wire   [63:0] loop_index69_cast_fu_136_p1;
reg   [60:0] loop_index69_fu_60;
wire   [60:0] empty_fu_114_p2;
wire    ap_loop_init;
reg    ap_done_reg;
wire    ap_continue_int;
reg    ap_done_int;
reg    ap_loop_exit_ready_pp0_iter2_reg;
reg   [0:0] ap_NS_fsm;
wire    ap_enable_pp0;
wire    ap_start_int;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_CS_fsm = 1'd1;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_done_reg = 1'b0;
end

kmeans_top_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(ap_start),
    .ap_ready(ap_ready),
    .ap_done(ap_done),
    .ap_start_int(ap_start_int),
    .ap_loop_init(ap_loop_init),
    .ap_ready_int(ap_ready_int),
    .ap_loop_exit_ready(ap_condition_exit_pp0_iter1_stage0),
    .ap_loop_exit_done(ap_done_int),
    .ap_continue_int(ap_continue_int),
    .ap_done_int(ap_done_int)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue_int == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter2_reg == 1'b1))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b1 == ap_condition_exit_pp0_iter1_stage0)) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_enable_reg_pp0_iter1 <= ap_start_int;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready == 1'b0))) begin
        ap_loop_exit_ready_pp0_iter2_reg <= 1'b0;
    end else if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_loop_exit_ready_pp0_iter2_reg <= ap_loop_exit_ready;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        if ((ap_loop_init == 1'b1)) begin
            loop_index69_fu_60 <= 61'd0;
        end else if (((exitcond85_fu_126_p2 == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
            loop_index69_fu_60 <= empty_fu_114_p2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        loop_index69_load_reg_157 <= loop_index69_fu_60;
        mem_addr_read_reg_162 <= m_axi_mem_RDATA;
        sext_ln182_cast_reg_147 <= sext_ln182_cast_fu_98_p1;
    end
end

always @ (*) begin
    if (((exitcond85_fu_126_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_condition_exit_pp0_iter1_stage0 = 1'b1;
    end else begin
        ap_condition_exit_pp0_iter1_stage0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter2_reg == 1'b1))) begin
        ap_done_int = 1'b1;
    end else begin
        ap_done_int = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_idle_pp0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_start_int == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_ready_int = 1'b1;
    end else begin
        ap_ready_int = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        m_axi_mem_RREADY = 1'b1;
    end else begin
        m_axi_mem_RREADY = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        mem_blk_n_R = m_axi_mem_RVALID;
    end else begin
        mem_blk_n_R = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        node_x_coords_ce1 = 1'b1;
    end else begin
        node_x_coords_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        node_x_coords_we1 = 1'b1;
    end else begin
        node_x_coords_we1 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_pp0_stage0 : begin
            ap_NS_fsm = ap_ST_fsm_pp0_stage0;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_pp0_stage0_11001 = ((m_axi_mem_RVALID == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b1));
end

always @ (*) begin
    ap_block_pp0_stage0_subdone = ((m_axi_mem_RVALID == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b1));
end

assign ap_block_state1_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state2_pp0_stage0_iter1 = (m_axi_mem_RVALID == 1'b0);
end

assign ap_block_state3_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_enable_reg_pp0_iter0 = ap_start_int;

assign ap_loop_exit_ready = ap_condition_exit_pp0_iter1_stage0;

assign empty_fu_114_p2 = (loop_index69_fu_60 + 61'd1);

assign exitcond85_fu_126_p2 = ((empty_fu_114_p2 == sext_ln182_cast_reg_147) ? 1'b1 : 1'b0);

assign loop_index69_cast_fu_136_p1 = loop_index69_load_reg_157;

assign m_axi_mem_ARADDR = 64'd0;

assign m_axi_mem_ARBURST = 2'd0;

assign m_axi_mem_ARCACHE = 4'd0;

assign m_axi_mem_ARID = 1'd0;

assign m_axi_mem_ARLEN = 32'd0;

assign m_axi_mem_ARLOCK = 2'd0;

assign m_axi_mem_ARPROT = 3'd0;

assign m_axi_mem_ARQOS = 4'd0;

assign m_axi_mem_ARREGION = 4'd0;

assign m_axi_mem_ARSIZE = 3'd0;

assign m_axi_mem_ARUSER = 1'd0;

assign m_axi_mem_ARVALID = 1'b0;

assign m_axi_mem_AWADDR = 64'd0;

assign m_axi_mem_AWBURST = 2'd0;

assign m_axi_mem_AWCACHE = 4'd0;

assign m_axi_mem_AWID = 1'd0;

assign m_axi_mem_AWLEN = 32'd0;

assign m_axi_mem_AWLOCK = 2'd0;

assign m_axi_mem_AWPROT = 3'd0;

assign m_axi_mem_AWQOS = 4'd0;

assign m_axi_mem_AWREGION = 4'd0;

assign m_axi_mem_AWSIZE = 3'd0;

assign m_axi_mem_AWUSER = 1'd0;

assign m_axi_mem_AWVALID = 1'b0;

assign m_axi_mem_BREADY = 1'b0;

assign m_axi_mem_WDATA = 64'd0;

assign m_axi_mem_WID = 1'd0;

assign m_axi_mem_WLAST = 1'b0;

assign m_axi_mem_WSTRB = 8'd0;

assign m_axi_mem_WUSER = 1'd0;

assign m_axi_mem_WVALID = 1'b0;

assign node_x_coords_address1 = loop_index69_cast_fu_136_p1;

assign node_x_coords_d1 = mem_addr_read_reg_162;

assign sext_ln182_cast_fu_98_p1 = $signed(sext_ln182);

endmodule //kmeans_top_kmeans_top_Pipeline_1


// Content from kmeans_top_kmeans_centroid_x_coords_next_RAM_AUTO_1R1W.v
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2022.2 (64-bit)
// Version: 2022.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module kmeans_top_kmeans_centroid_x_coords_next_RAM_AUTO_1R1W (
     
    address0, ce0,
    d0, we0, 
    q0, 
     
    reset, clk);

parameter DataWidth = 64;
parameter AddressWidth = 8;
parameter AddressRange = 256;
 
input[AddressWidth-1:0] address0;
input ce0;
input[DataWidth-1:0] d0;
input we0; 
output reg[DataWidth-1:0] q0; 

input reset;
input clk;

(* ram_style = "auto"  *)reg [DataWidth-1:0] ram[0:AddressRange-1];


 





//read first
always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram[address0] <= d0; 
        q0 <= ram[address0];

    end
end 
 
 

endmodule



// Content from kmeans_top_mul_64s_64s_64_1_1.v
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2022.2 (64-bit)
// Version: 2022.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// ==============================================================

`timescale 1 ns / 1 ps

module kmeans_top_mul_64s_64s_64_1_1(din0, din1, dout);
parameter ID = 1;
parameter NUM_STAGE = 0;
parameter din0_WIDTH = 14;
parameter din1_WIDTH = 12;
parameter dout_WIDTH = 26;
input [din0_WIDTH - 1 : 0] din0; 
input [din1_WIDTH - 1 : 0] din1; 
output [dout_WIDTH - 1 : 0] dout;

assign dout = $signed(din0) * $signed(din1);
endmodule


// Content from kmeans_top_kmeans_top_Pipeline_4.v
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2022.2 (64-bit)
// Version: 2022.2
// Copyright (C) Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module kmeans_top_kmeans_top_Pipeline_4 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        m_axi_mem_AWVALID,
        m_axi_mem_AWREADY,
        m_axi_mem_AWADDR,
        m_axi_mem_AWID,
        m_axi_mem_AWLEN,
        m_axi_mem_AWSIZE,
        m_axi_mem_AWBURST,
        m_axi_mem_AWLOCK,
        m_axi_mem_AWCACHE,
        m_axi_mem_AWPROT,
        m_axi_mem_AWQOS,
        m_axi_mem_AWREGION,
        m_axi_mem_AWUSER,
        m_axi_mem_WVALID,
        m_axi_mem_WREADY,
        m_axi_mem_WDATA,
        m_axi_mem_WSTRB,
        m_axi_mem_WLAST,
        m_axi_mem_WID,
        m_axi_mem_WUSER,
        m_axi_mem_ARVALID,
        m_axi_mem_ARREADY,
        m_axi_mem_ARADDR,
        m_axi_mem_ARID,
        m_axi_mem_ARLEN,
        m_axi_mem_ARSIZE,
        m_axi_mem_ARBURST,
        m_axi_mem_ARLOCK,
        m_axi_mem_ARCACHE,
        m_axi_mem_ARPROT,
        m_axi_mem_ARQOS,
        m_axi_mem_ARREGION,
        m_axi_mem_ARUSER,
        m_axi_mem_RVALID,
        m_axi_mem_RREADY,
        m_axi_mem_RDATA,
        m_axi_mem_RLAST,
        m_axi_mem_RID,
        m_axi_mem_RFIFONUM,
        m_axi_mem_RUSER,
        m_axi_mem_RRESP,
        m_axi_mem_BVALID,
        m_axi_mem_BREADY,
        m_axi_mem_BRESP,
        m_axi_mem_BID,
        m_axi_mem_BUSER,
        p_cast1_cast,
        centroid_x_coords_address0,
        centroid_x_coords_ce0,
        centroid_x_coords_we0,
        centroid_x_coords_d0,
        sext_ln185
);

parameter    ap_ST_fsm_pp0_stage0 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
output   m_axi_mem_AWVALID;
input   m_axi_mem_AWREADY;
output  [63:0] m_axi_mem_AWADDR;
output  [0:0] m_axi_mem_AWID;
output  [31:0] m_axi_mem_AWLEN;
output  [2:0] m_axi_mem_AWSIZE;
output  [1:0] m_axi_mem_AWBURST;
output  [1:0] m_axi_mem_AWLOCK;
output  [3:0] m_axi_mem_AWCACHE;
output  [2:0] m_axi_mem_AWPROT;
output  [3:0] m_axi_mem_AWQOS;
output  [3:0] m_axi_mem_AWREGION;
output  [0:0] m_axi_mem_AWUSER;
output   m_axi_mem_WVALID;
input   m_axi_mem_WREADY;
output  [63:0] m_axi_mem_WDATA;
output  [7:0] m_axi_mem_WSTRB;
output   m_axi_mem_WLAST;
output  [0:0] m_axi_mem_WID;
output  [0:0] m_axi_mem_WUSER;
output   m_axi_mem_ARVALID;
input   m_axi_mem_ARREADY;
output  [63:0] m_axi_mem_ARADDR;
output  [0:0] m_axi_mem_ARID;
output  [31:0] m_axi_mem_ARLEN;
output  [2:0] m_axi_mem_ARSIZE;
output  [1:0] m_axi_mem_ARBURST;
output  [1:0] m_axi_mem_ARLOCK;
output  [3:0] m_axi_mem_ARCACHE;
output  [2:0] m_axi_mem_ARPROT;
output  [3:0] m_axi_mem_ARQOS;
output  [3:0] m_axi_mem_ARREGION;
output  [0:0] m_axi_mem_ARUSER;
input   m_axi_mem_RVALID;
output   m_axi_mem_RREADY;
input  [63:0] m_axi_mem_RDATA;
input   m_axi_mem_RLAST;
input  [0:0] m_axi_mem_RID;
input  [8:0] m_axi_mem_RFIFONUM;
input  [0:0] m_axi_mem_RUSER;
input  [1:0] m_axi_mem_RRESP;
input   m_axi_mem_BVALID;
output   m_axi_mem_BREADY;
input  [1:0] m_axi_mem_BRESP;
input  [0:0] m_axi_mem_BID;
input  [0:0] m_axi_mem_BUSER;
input  [60:0] p_cast1_cast;
output  [7:0] centroid_x_coords_address0;
output   centroid_x_coords_ce0;
output   centroid_x_coords_we0;
output  [63:0] centroid_x_coords_d0;
input  [31:0] sext_ln185;

reg ap_idle;
reg m_axi_mem_RREADY;
reg centroid_x_coords_ce0;
reg centroid_x_coords_we0;

(* fsm_encoding = "none" *) reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_enable_reg_pp0_iter0;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter2;
reg    ap_idle_pp0;
wire    ap_block_state1_pp0_stage0_iter0;
reg    ap_block_state2_pp0_stage0_iter1;
wire    ap_block_state3_pp0_stage0_iter2;
reg    ap_block_pp0_stage0_subdone;
wire   [0:0] exitcond82_fu_114_p2;
reg    ap_condition_exit_pp0_iter1_stage0;
wire    ap_loop_exit_ready;
reg    ap_ready_int;
reg    mem_blk_n_R;
wire    ap_block_pp0_stage0;
wire  signed [60:0] sext_ln185_cast_fu_86_p1;
reg  signed [60:0] sext_ln185_cast_reg_135;
reg    ap_block_pp0_stage0_11001;
reg   [60:0] loop_index51_load_reg_145;
reg   [63:0] mem_addr_read_reg_150;
wire   [63:0] loop_index51_cast_fu_124_p1;
reg   [60:0] loop_index51_fu_52;
wire   [60:0] empty_fu_102_p2;
wire    ap_loop_init;
reg    ap_done_reg;
wire    ap_continue_int;
reg    ap_done_int;
reg    ap_loop_exit_ready_pp0_iter2_reg;
reg   [0:0] ap_NS_fsm;
wire    ap_enable_pp0;
wire    ap_start_int;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_CS_fsm = 1'd1;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_done_reg = 1'b0;
end

kmeans_top_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(ap_start),
    .ap_ready(ap_ready),
    .ap_done(ap_done),
    .ap_start_int(ap_start_int),
    .ap_loop_init(ap_loop_init),
    .ap_ready_int(ap_ready_int),
    .ap_loop_exit_ready(ap_condition_exit_pp0_iter1_stage0),
    .ap_loop_exit_done(ap_done_int),
    .ap_continue_int(ap_continue_int),
    .ap_done_int(ap_done_int)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue_int == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter2_reg == 1'b1))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b1 == ap_condition_exit_pp0_iter1_stage0)) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_enable_reg_pp0_iter1 <= ap_start_int;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready == 1'b0))) begin
        ap_loop_exit_ready_pp0_iter2_reg <= 1'b0;
    end else if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_loop_exit_ready_pp0_iter2_reg <= ap_loop_exit_ready;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        if ((ap_loop_init == 1'b1)) begin
            loop_index51_fu_52 <= 61'd0;
        end else if (((exitcond82_fu_114_p2 == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
            loop_index51_fu_52 <= empty_fu_102_p2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        loop_index51_load_reg_145 <= loop_index51_fu_52;
        mem_addr_read_reg_150 <= m_axi_mem_RDATA;
        sext_ln185_cast_reg_135 <= sext_ln185_cast_fu_86_p1;
    end
end

always @ (*) begin
    if (((exitcond82_fu_114_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_condition_exit_pp0_iter1_stage0 = 1'b1;
    end else begin
        ap_condition_exit_pp0_iter1_stage0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter2_reg == 1'b1))) begin
        ap_done_int = 1'b1;
    end else begin
        ap_done_int = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_idle_pp0 == 1'b1) & (ap_start_int == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_ready_int = 1'b1;
    end else begin
        ap_ready_int = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        centroid_x_coords_ce0 = 1'b1;
    end else begin
        centroid_x_coords_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        centroid_x_coords_we0 = 1'b1;
    end else begin
        centroid_x_coords_we0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        m_axi_mem_RREADY = 1'b1;
    end else begin
        m_axi_mem_RREADY = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        mem_blk_n_R = m_axi_mem_RVALID;
    end else begin
        mem_blk_n_R = 1'b1;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_pp0_stage0 : begin
            ap_NS_fsm = ap_ST_fsm_pp0_stage0;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_pp0_stage0_11001 = ((m_axi_mem_RVALID == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b1));
end

always @ (*) begin
    ap_block_pp0_stage0_subdone = ((m_axi_mem_RVALID == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b1));
end

assign ap_block_state1_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_state2_pp0_stage0_iter1 = (m_axi_mem_RVALID == 1'b0);
end

assign ap_block_state3_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_enable_reg_pp0_iter0 = ap_start_int;

assign ap_loop_exit_ready = ap_condition_exit_pp0_iter1_stage0;

assign centroid_x_coords_address0 = loop_index51_cast_fu_124_p1;

assign centroid_x_coords_d0 = mem_addr_read_reg_150;

assign empty_fu_102_p2 = (loop_index51_fu_52 + 61'd1);

assign exitcond82_fu_114_p2 = ((empty_fu_102_p2 == sext_ln185_cast_reg_135) ? 1'b1 : 1'b0);

assign loop_index51_cast_fu_124_p1 = loop_index51_load_reg_145;

assign m_axi_mem_ARADDR = 64'd0;

assign m_axi_mem_ARBURST = 2'd0;

assign m_axi_mem_ARCACHE = 4'd0;

assign m_axi_mem_ARID = 1'd0;

assign m_axi_mem_ARLEN = 32'd0;

assign m_axi_mem_ARLOCK = 2'd0;

assign m_axi_mem_ARPROT = 3'd0;

assign m_axi_mem_ARQOS = 4'd0;

assign m_axi_mem_ARREGION = 4'd0;

assign m_axi_mem_ARSIZE = 3'd0;

assign m_axi_mem_ARUSER = 1'd0;

assign m_axi_mem_ARVALID = 1'b0;

assign m_axi_mem_AWADDR = 64'd0;

assign m_axi_mem_AWBURST = 2'd0;

assign m_axi_mem_AWCACHE = 4'd0;

assign m_axi_mem_AWID = 1'd0;

assign m_axi_mem_AWLEN = 32'd0;

assign m_axi_mem_AWLOCK = 2'd0;

assign m_axi_mem_AWPROT = 3'd0;

assign m_axi_mem_AWQOS = 4'd0;

assign m_axi_mem_AWREGION = 4'd0;

assign m_axi_mem_AWSIZE = 3'd0;

assign m_axi_mem_AWUSER = 1'd0;

assign m_axi_mem_AWVALID = 1'b0;

assign m_axi_mem_BREADY = 1'b0;

assign m_axi_mem_WDATA = 64'd0;

assign m_axi_mem_WID = 1'd0;

assign m_axi_mem_WLAST = 1'b0;

assign m_axi_mem_WSTRB = 8'd0;

assign m_axi_mem_WUSER = 1'd0;

assign m_axi_mem_WVALID = 1'b0;

assign sext_ln185_cast_fu_86_p1 = $signed(sext_ln185);

endmodule //kmeans_top_kmeans_top_Pipeline_4


// Content from kmeans_top_kmeans_top_Pipeline_12.v
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2022.2 (64-bit)
// Version: 2022.2
// Copyright (C) Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module kmeans_top_kmeans_top_Pipeline_12 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        m_axi_mem_AWVALID,
        m_axi_mem_AWREADY,
        m_axi_mem_AWADDR,
        m_axi_mem_AWID,
        m_axi_mem_AWLEN,
        m_axi_mem_AWSIZE,
        m_axi_mem_AWBURST,
        m_axi_mem_AWLOCK,
        m_axi_mem_AWCACHE,
        m_axi_mem_AWPROT,
        m_axi_mem_AWQOS,
        m_axi_mem_AWREGION,
        m_axi_mem_AWUSER,
        m_axi_mem_WVALID,
        m_axi_mem_WREADY,
        m_axi_mem_WDATA,
        m_axi_mem_WSTRB,
        m_axi_mem_WLAST,
        m_axi_mem_WID,
        m_axi_mem_WUSER,
        m_axi_mem_ARVALID,
        m_axi_mem_ARREADY,
        m_axi_mem_ARADDR,
        m_axi_mem_ARID,
        m_axi_mem_ARLEN,
        m_axi_mem_ARSIZE,
        m_axi_mem_ARBURST,
        m_axi_mem_ARLOCK,
        m_axi_mem_ARCACHE,
        m_axi_mem_ARPROT,
        m_axi_mem_ARQOS,
        m_axi_mem_ARREGION,
        m_axi_mem_ARUSER,
        m_axi_mem_RVALID,
        m_axi_mem_RREADY,
        m_axi_mem_RDATA,
        m_axi_mem_RLAST,
        m_axi_mem_RID,
        m_axi_mem_RFIFONUM,
        m_axi_mem_RUSER,
        m_axi_mem_RRESP,
        m_axi_mem_BVALID,
        m_axi_mem_BREADY,
        m_axi_mem_BRESP,
        m_axi_mem_BID,
        m_axi_mem_BUSER,
        p_cast7_cast,
        centroid_x_coords_address0,
        centroid_x_coords_ce0,
        centroid_x_coords_q0,
        sext_ln185
);

parameter    ap_ST_fsm_pp0_stage0 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
output   m_axi_mem_AWVALID;
input   m_axi_mem_AWREADY;
output  [63:0] m_axi_mem_AWADDR;
output  [0:0] m_axi_mem_AWID;
output  [31:0] m_axi_mem_AWLEN;
output  [2:0] m_axi_mem_AWSIZE;
output  [1:0] m_axi_mem_AWBURST;
output  [1:0] m_axi_mem_AWLOCK;
output  [3:0] m_axi_mem_AWCACHE;
output  [2:0] m_axi_mem_AWPROT;
output  [3:0] m_axi_mem_AWQOS;
output  [3:0] m_axi_mem_AWREGION;
output  [0:0] m_axi_mem_AWUSER;
output   m_axi_mem_WVALID;
input   m_axi_mem_WREADY;
output  [63:0] m_axi_mem_WDATA;
output  [7:0] m_axi_mem_WSTRB;
output   m_axi_mem_WLAST;
output  [0:0] m_axi_mem_WID;
output  [0:0] m_axi_mem_WUSER;
output   m_axi_mem_ARVALID;
input   m_axi_mem_ARREADY;
output  [63:0] m_axi_mem_ARADDR;
output  [0:0] m_axi_mem_ARID;
output  [31:0] m_axi_mem_ARLEN;
output  [2:0] m_axi_mem_ARSIZE;
output  [1:0] m_axi_mem_ARBURST;
output  [1:0] m_axi_mem_ARLOCK;
output  [3:0] m_axi_mem_ARCACHE;
output  [2:0] m_axi_mem_ARPROT;
output  [3:0] m_axi_mem_ARQOS;
output  [3:0] m_axi_mem_ARREGION;
output  [0:0] m_axi_mem_ARUSER;
input   m_axi_mem_RVALID;
output   m_axi_mem_RREADY;
input  [63:0] m_axi_mem_RDATA;
input   m_axi_mem_RLAST;
input  [0:0] m_axi_mem_RID;
input  [8:0] m_axi_mem_RFIFONUM;
input  [0:0] m_axi_mem_RUSER;
input  [1:0] m_axi_mem_RRESP;
input   m_axi_mem_BVALID;
output   m_axi_mem_BREADY;
input  [1:0] m_axi_mem_BRESP;
input  [0:0] m_axi_mem_BID;
input  [0:0] m_axi_mem_BUSER;
input  [60:0] p_cast7_cast;
output  [7:0] centroid_x_coords_address0;
output   centroid_x_coords_ce0;
input  [63:0] centroid_x_coords_q0;
input  [31:0] sext_ln185;

reg ap_idle;
reg m_axi_mem_WVALID;
reg centroid_x_coords_ce0;

(* fsm_encoding = "none" *) reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_enable_reg_pp0_iter0;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter2;
reg    ap_enable_reg_pp0_iter3;
reg    ap_idle_pp0;
wire    ap_block_state1_pp0_stage0_iter0;
wire    ap_block_state2_pp0_stage0_iter1;
wire    ap_block_state3_pp0_stage0_iter2;
wire    ap_block_state4_pp0_stage0_iter3;
reg    ap_block_pp0_stage0_subdone;
wire   [0:0] exitcond74_fu_118_p2;
reg    ap_condition_exit_pp0_iter1_stage0;
wire    ap_loop_exit_ready;
reg    ap_ready_int;
reg    mem_blk_n_W;
wire    ap_block_pp0_stage0;
wire  signed [60:0] sext_ln185_cast_fu_91_p1;
reg  signed [60:0] sext_ln185_cast_reg_141;
reg    ap_block_pp0_stage0_11001;
reg   [63:0] centroid_x_coords_load_reg_160;
wire   [63:0] loop_index3_cast_fu_113_p1;
wire    ap_block_pp0_stage0_01001;
reg   [60:0] loop_index3_fu_54;
wire   [60:0] empty_fu_107_p2;
wire    ap_loop_init;
reg    ap_done_reg;
wire    ap_continue_int;
reg    ap_done_int;
reg    ap_loop_exit_ready_pp0_iter2_reg;
reg    ap_loop_exit_ready_pp0_iter3_reg;
reg   [0:0] ap_NS_fsm;
wire    ap_enable_pp0;
wire    ap_start_int;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_CS_fsm = 1'd1;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_done_reg = 1'b0;
end

kmeans_top_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(ap_start),
    .ap_ready(ap_ready),
    .ap_done(ap_done),
    .ap_start_int(ap_start_int),
    .ap_loop_init(ap_loop_init),
    .ap_ready_int(ap_ready_int),
    .ap_loop_exit_ready(ap_condition_exit_pp0_iter1_stage0),
    .ap_loop_exit_done(ap_done_int),
    .ap_continue_int(ap_continue_int),
    .ap_done_int(ap_done_int)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue_int == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter3_reg == 1'b1))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b1 == ap_condition_exit_pp0_iter1_stage0)) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_enable_reg_pp0_iter1 <= ap_start_int;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter2_reg == 1'b0))) begin
        ap_loop_exit_ready_pp0_iter3_reg <= 1'b0;
    end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        ap_loop_exit_ready_pp0_iter3_reg <= ap_loop_exit_ready_pp0_iter2_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        if ((ap_loop_init == 1'b1)) begin
            loop_index3_fu_54 <= 61'd0;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (exitcond74_fu_118_p2 == 1'd0))) begin
            loop_index3_fu_54 <= empty_fu_107_p2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_loop_exit_ready_pp0_iter2_reg <= ap_loop_exit_ready;
        sext_ln185_cast_reg_141 <= sext_ln185_cast_fu_91_p1;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        centroid_x_coords_load_reg_160 <= centroid_x_coords_q0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (exitcond74_fu_118_p2 == 1'd1))) begin
        ap_condition_exit_pp0_iter1_stage0 = 1'b1;
    end else begin
        ap_condition_exit_pp0_iter1_stage0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter3_reg == 1'b1))) begin
        ap_done_int = 1'b1;
    end else begin
        ap_done_int = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_idle_pp0 == 1'b1) & (ap_start_int == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_ready_int = 1'b1;
    end else begin
        ap_ready_int = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        centroid_x_coords_ce0 = 1'b1;
    end else begin
        centroid_x_coords_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1))) begin
        m_axi_mem_WVALID = 1'b1;
    end else begin
        m_axi_mem_WVALID = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter3 == 1'b1))) begin
        mem_blk_n_W = m_axi_mem_WREADY;
    end else begin
        mem_blk_n_W = 1'b1;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_pp0_stage0 : begin
            ap_NS_fsm = ap_ST_fsm_pp0_stage0;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_01001 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_pp0_stage0_11001 = ((m_axi_mem_WREADY == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b1));
end

always @ (*) begin
    ap_block_pp0_stage0_subdone = ((m_axi_mem_WREADY == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b1));
end

assign ap_block_state1_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_enable_reg_pp0_iter0 = ap_start_int;

assign ap_loop_exit_ready = ap_condition_exit_pp0_iter1_stage0;

assign centroid_x_coords_address0 = loop_index3_cast_fu_113_p1;

assign empty_fu_107_p2 = (loop_index3_fu_54 + 61'd1);

assign exitcond74_fu_118_p2 = ((empty_fu_107_p2 == sext_ln185_cast_reg_141) ? 1'b1 : 1'b0);

assign loop_index3_cast_fu_113_p1 = loop_index3_fu_54;

assign m_axi_mem_ARADDR = 64'd0;

assign m_axi_mem_ARBURST = 2'd0;

assign m_axi_mem_ARCACHE = 4'd0;

assign m_axi_mem_ARID = 1'd0;

assign m_axi_mem_ARLEN = 32'd0;

assign m_axi_mem_ARLOCK = 2'd0;

assign m_axi_mem_ARPROT = 3'd0;

assign m_axi_mem_ARQOS = 4'd0;

assign m_axi_mem_ARREGION = 4'd0;

assign m_axi_mem_ARSIZE = 3'd0;

assign m_axi_mem_ARUSER = 1'd0;

assign m_axi_mem_ARVALID = 1'b0;

assign m_axi_mem_AWADDR = 64'd0;

assign m_axi_mem_AWBURST = 2'd0;

assign m_axi_mem_AWCACHE = 4'd0;

assign m_axi_mem_AWID = 1'd0;

assign m_axi_mem_AWLEN = 32'd0;

assign m_axi_mem_AWLOCK = 2'd0;

assign m_axi_mem_AWPROT = 3'd0;

assign m_axi_mem_AWQOS = 4'd0;

assign m_axi_mem_AWREGION = 4'd0;

assign m_axi_mem_AWSIZE = 3'd0;

assign m_axi_mem_AWUSER = 1'd0;

assign m_axi_mem_AWVALID = 1'b0;

assign m_axi_mem_BREADY = 1'b0;

assign m_axi_mem_RREADY = 1'b0;

assign m_axi_mem_WDATA = centroid_x_coords_load_reg_160;

assign m_axi_mem_WID = 1'd0;

assign m_axi_mem_WLAST = 1'b0;

assign m_axi_mem_WSTRB = 8'd255;

assign m_axi_mem_WUSER = 1'd0;

assign sext_ln185_cast_fu_91_p1 = $signed(sext_ln185);

endmodule //kmeans_top_kmeans_top_Pipeline_12


// Content from kmeans_top_kmeans_top_Pipeline_8.v
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2022.2 (64-bit)
// Version: 2022.2
// Copyright (C) Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module kmeans_top_kmeans_top_Pipeline_8 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        m_axi_mem_AWVALID,
        m_axi_mem_AWREADY,
        m_axi_mem_AWADDR,
        m_axi_mem_AWID,
        m_axi_mem_AWLEN,
        m_axi_mem_AWSIZE,
        m_axi_mem_AWBURST,
        m_axi_mem_AWLOCK,
        m_axi_mem_AWCACHE,
        m_axi_mem_AWPROT,
        m_axi_mem_AWQOS,
        m_axi_mem_AWREGION,
        m_axi_mem_AWUSER,
        m_axi_mem_WVALID,
        m_axi_mem_WREADY,
        m_axi_mem_WDATA,
        m_axi_mem_WSTRB,
        m_axi_mem_WLAST,
        m_axi_mem_WID,
        m_axi_mem_WUSER,
        m_axi_mem_ARVALID,
        m_axi_mem_ARREADY,
        m_axi_mem_ARADDR,
        m_axi_mem_ARID,
        m_axi_mem_ARLEN,
        m_axi_mem_ARSIZE,
        m_axi_mem_ARBURST,
        m_axi_mem_ARLOCK,
        m_axi_mem_ARCACHE,
        m_axi_mem_ARPROT,
        m_axi_mem_ARQOS,
        m_axi_mem_ARREGION,
        m_axi_mem_ARUSER,
        m_axi_mem_RVALID,
        m_axi_mem_RREADY,
        m_axi_mem_RDATA,
        m_axi_mem_RLAST,
        m_axi_mem_RID,
        m_axi_mem_RFIFONUM,
        m_axi_mem_RUSER,
        m_axi_mem_RRESP,
        m_axi_mem_BVALID,
        m_axi_mem_BREADY,
        m_axi_mem_BRESP,
        m_axi_mem_BID,
        m_axi_mem_BUSER,
        p_cast13_cast,
        centroid_y_coords_address0,
        centroid_y_coords_ce0,
        centroid_y_coords_q0,
        sext_ln185
);

parameter    ap_ST_fsm_pp0_stage0 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
output   m_axi_mem_AWVALID;
input   m_axi_mem_AWREADY;
output  [63:0] m_axi_mem_AWADDR;
output  [0:0] m_axi_mem_AWID;
output  [31:0] m_axi_mem_AWLEN;
output  [2:0] m_axi_mem_AWSIZE;
output  [1:0] m_axi_mem_AWBURST;
output  [1:0] m_axi_mem_AWLOCK;
output  [3:0] m_axi_mem_AWCACHE;
output  [2:0] m_axi_mem_AWPROT;
output  [3:0] m_axi_mem_AWQOS;
output  [3:0] m_axi_mem_AWREGION;
output  [0:0] m_axi_mem_AWUSER;
output   m_axi_mem_WVALID;
input   m_axi_mem_WREADY;
output  [63:0] m_axi_mem_WDATA;
output  [7:0] m_axi_mem_WSTRB;
output   m_axi_mem_WLAST;
output  [0:0] m_axi_mem_WID;
output  [0:0] m_axi_mem_WUSER;
output   m_axi_mem_ARVALID;
input   m_axi_mem_ARREADY;
output  [63:0] m_axi_mem_ARADDR;
output  [0:0] m_axi_mem_ARID;
output  [31:0] m_axi_mem_ARLEN;
output  [2:0] m_axi_mem_ARSIZE;
output  [1:0] m_axi_mem_ARBURST;
output  [1:0] m_axi_mem_ARLOCK;
output  [3:0] m_axi_mem_ARCACHE;
output  [2:0] m_axi_mem_ARPROT;
output  [3:0] m_axi_mem_ARQOS;
output  [3:0] m_axi_mem_ARREGION;
output  [0:0] m_axi_mem_ARUSER;
input   m_axi_mem_RVALID;
output   m_axi_mem_RREADY;
input  [63:0] m_axi_mem_RDATA;
input   m_axi_mem_RLAST;
input  [0:0] m_axi_mem_RID;
input  [8:0] m_axi_mem_RFIFONUM;
input  [0:0] m_axi_mem_RUSER;
input  [1:0] m_axi_mem_RRESP;
input   m_axi_mem_BVALID;
output   m_axi_mem_BREADY;
input  [1:0] m_axi_mem_BRESP;
input  [0:0] m_axi_mem_BID;
input  [0:0] m_axi_mem_BUSER;
input  [60:0] p_cast13_cast;
output  [7:0] centroid_y_coords_address0;
output   centroid_y_coords_ce0;
input  [63:0] centroid_y_coords_q0;
input  [31:0] sext_ln185;

reg ap_idle;
reg m_axi_mem_WVALID;
reg centroid_y_coords_ce0;

(* fsm_encoding = "none" *) reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_enable_reg_pp0_iter0;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter2;
reg    ap_enable_reg_pp0_iter3;
reg    ap_idle_pp0;
wire    ap_block_state1_pp0_stage0_iter0;
wire    ap_block_state2_pp0_stage0_iter1;
wire    ap_block_state3_pp0_stage0_iter2;
wire    ap_block_state4_pp0_stage0_iter3;
reg    ap_block_pp0_stage0_subdone;
wire   [0:0] exitcond80_fu_118_p2;
reg    ap_condition_exit_pp0_iter1_stage0;
wire    ap_loop_exit_ready;
reg    ap_ready_int;
reg    mem_blk_n_W;
wire    ap_block_pp0_stage0;
wire  signed [60:0] sext_ln185_cast_fu_91_p1;
reg  signed [60:0] sext_ln185_cast_reg_141;
reg    ap_block_pp0_stage0_11001;
reg   [63:0] centroid_y_coords_load_reg_160;
wire   [63:0] loop_index27_cast_fu_113_p1;
wire    ap_block_pp0_stage0_01001;
reg   [60:0] loop_index27_fu_54;
wire   [60:0] empty_fu_107_p2;
wire    ap_loop_init;
reg    ap_done_reg;
wire    ap_continue_int;
reg    ap_done_int;
reg    ap_loop_exit_ready_pp0_iter2_reg;
reg    ap_loop_exit_ready_pp0_iter3_reg;
reg   [0:0] ap_NS_fsm;
wire    ap_enable_pp0;
wire    ap_start_int;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_CS_fsm = 1'd1;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_done_reg = 1'b0;
end

kmeans_top_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(ap_start),
    .ap_ready(ap_ready),
    .ap_done(ap_done),
    .ap_start_int(ap_start_int),
    .ap_loop_init(ap_loop_init),
    .ap_ready_int(ap_ready_int),
    .ap_loop_exit_ready(ap_condition_exit_pp0_iter1_stage0),
    .ap_loop_exit_done(ap_done_int),
    .ap_continue_int(ap_continue_int),
    .ap_done_int(ap_done_int)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue_int == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter3_reg == 1'b1))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b1 == ap_condition_exit_pp0_iter1_stage0)) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_enable_reg_pp0_iter1 <= ap_start_int;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter2_reg == 1'b0))) begin
        ap_loop_exit_ready_pp0_iter3_reg <= 1'b0;
    end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        ap_loop_exit_ready_pp0_iter3_reg <= ap_loop_exit_ready_pp0_iter2_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        if ((ap_loop_init == 1'b1)) begin
            loop_index27_fu_54 <= 61'd0;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (exitcond80_fu_118_p2 == 1'd0))) begin
            loop_index27_fu_54 <= empty_fu_107_p2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_loop_exit_ready_pp0_iter2_reg <= ap_loop_exit_ready;
        sext_ln185_cast_reg_141 <= sext_ln185_cast_fu_91_p1;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        centroid_y_coords_load_reg_160 <= centroid_y_coords_q0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (exitcond80_fu_118_p2 == 1'd1))) begin
        ap_condition_exit_pp0_iter1_stage0 = 1'b1;
    end else begin
        ap_condition_exit_pp0_iter1_stage0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter3_reg == 1'b1))) begin
        ap_done_int = 1'b1;
    end else begin
        ap_done_int = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_idle_pp0 == 1'b1) & (ap_start_int == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_ready_int = 1'b1;
    end else begin
        ap_ready_int = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        centroid_y_coords_ce0 = 1'b1;
    end else begin
        centroid_y_coords_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter3 == 1'b1))) begin
        m_axi_mem_WVALID = 1'b1;
    end else begin
        m_axi_mem_WVALID = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter3 == 1'b1))) begin
        mem_blk_n_W = m_axi_mem_WREADY;
    end else begin
        mem_blk_n_W = 1'b1;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_pp0_stage0 : begin
            ap_NS_fsm = ap_ST_fsm_pp0_stage0;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_01001 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_pp0_stage0_11001 = ((m_axi_mem_WREADY == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b1));
end

always @ (*) begin
    ap_block_pp0_stage0_subdone = ((m_axi_mem_WREADY == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b1));
end

assign ap_block_state1_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage0_iter3 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_enable_reg_pp0_iter0 = ap_start_int;

assign ap_loop_exit_ready = ap_condition_exit_pp0_iter1_stage0;

assign centroid_y_coords_address0 = loop_index27_cast_fu_113_p1;

assign empty_fu_107_p2 = (loop_index27_fu_54 + 61'd1);

assign exitcond80_fu_118_p2 = ((empty_fu_107_p2 == sext_ln185_cast_reg_141) ? 1'b1 : 1'b0);

assign loop_index27_cast_fu_113_p1 = loop_index27_fu_54;

assign m_axi_mem_ARADDR = 64'd0;

assign m_axi_mem_ARBURST = 2'd0;

assign m_axi_mem_ARCACHE = 4'd0;

assign m_axi_mem_ARID = 1'd0;

assign m_axi_mem_ARLEN = 32'd0;

assign m_axi_mem_ARLOCK = 2'd0;

assign m_axi_mem_ARPROT = 3'd0;

assign m_axi_mem_ARQOS = 4'd0;

assign m_axi_mem_ARREGION = 4'd0;

assign m_axi_mem_ARSIZE = 3'd0;

assign m_axi_mem_ARUSER = 1'd0;

assign m_axi_mem_ARVALID = 1'b0;

assign m_axi_mem_AWADDR = 64'd0;

assign m_axi_mem_AWBURST = 2'd0;

assign m_axi_mem_AWCACHE = 4'd0;

assign m_axi_mem_AWID = 1'd0;

assign m_axi_mem_AWLEN = 32'd0;

assign m_axi_mem_AWLOCK = 2'd0;

assign m_axi_mem_AWPROT = 3'd0;

assign m_axi_mem_AWQOS = 4'd0;

assign m_axi_mem_AWREGION = 4'd0;

assign m_axi_mem_AWSIZE = 3'd0;

assign m_axi_mem_AWUSER = 1'd0;

assign m_axi_mem_AWVALID = 1'b0;

assign m_axi_mem_BREADY = 1'b0;

assign m_axi_mem_RREADY = 1'b0;

assign m_axi_mem_WDATA = centroid_y_coords_load_reg_160;

assign m_axi_mem_WID = 1'd0;

assign m_axi_mem_WLAST = 1'b0;

assign m_axi_mem_WSTRB = 8'd255;

assign m_axi_mem_WUSER = 1'd0;

assign sext_ln185_cast_fu_91_p1 = $signed(sext_ln185);

endmodule //kmeans_top_kmeans_top_Pipeline_8


// Content from kmeans_top_kmeans_Pipeline_VITIS_LOOP_73_3.v
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2022.2 (64-bit)
// Version: 2022.2
// Copyright (C) Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module kmeans_top_kmeans_Pipeline_VITIS_LOOP_73_3 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        node_x_coords_address0,
        node_x_coords_ce0,
        node_x_coords_q0,
        node_x_coords_address1,
        node_x_coords_ce1,
        node_x_coords_q1,
        zext_ln69,
        node_y_coords_address0,
        node_y_coords_ce0,
        node_y_coords_q0,
        node_y_coords_address1,
        node_y_coords_ce1,
        node_y_coords_q1,
        k,
        centroid_y_coords_address0,
        centroid_y_coords_ce0,
        centroid_y_coords_q0,
        centroid_y_coords_address1,
        centroid_y_coords_ce1,
        centroid_y_coords_q1,
        centroid_x_coords_address0,
        centroid_x_coords_ce0,
        centroid_x_coords_q0,
        centroid_x_coords_address1,
        centroid_x_coords_ce1,
        centroid_x_coords_q1,
        min_dist_index_out,
        min_dist_index_out_ap_vld
);

parameter    ap_ST_fsm_pp0_stage0 = 2'd1;
parameter    ap_ST_fsm_pp0_stage1 = 2'd2;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
output  [12:0] node_x_coords_address0;
output   node_x_coords_ce0;
input  [63:0] node_x_coords_q0;
output  [12:0] node_x_coords_address1;
output   node_x_coords_ce1;
input  [63:0] node_x_coords_q1;
input  [12:0] zext_ln69;
output  [12:0] node_y_coords_address0;
output   node_y_coords_ce0;
input  [63:0] node_y_coords_q0;
output  [12:0] node_y_coords_address1;
output   node_y_coords_ce1;
input  [63:0] node_y_coords_q1;
input  [31:0] k;
output  [7:0] centroid_y_coords_address0;
output   centroid_y_coords_ce0;
input  [63:0] centroid_y_coords_q0;
output  [7:0] centroid_y_coords_address1;
output   centroid_y_coords_ce1;
input  [63:0] centroid_y_coords_q1;
output  [7:0] centroid_x_coords_address0;
output   centroid_x_coords_ce0;
input  [63:0] centroid_x_coords_q0;
output  [7:0] centroid_x_coords_address1;
output   centroid_x_coords_ce1;
input  [63:0] centroid_x_coords_q1;
output  [31:0] min_dist_index_out;
output   min_dist_index_out_ap_vld;

reg ap_idle;
reg[12:0] node_x_coords_address0;
reg node_x_coords_ce0;
reg[12:0] node_x_coords_address1;
reg node_x_coords_ce1;
reg[12:0] node_y_coords_address0;
reg node_y_coords_ce0;
reg[12:0] node_y_coords_address1;
reg node_y_coords_ce1;
reg[7:0] centroid_y_coords_address0;
reg centroid_y_coords_ce0;
reg[7:0] centroid_y_coords_address1;
reg centroid_y_coords_ce1;
reg[7:0] centroid_x_coords_address0;
reg centroid_x_coords_ce0;
reg[7:0] centroid_x_coords_address1;
reg centroid_x_coords_ce1;
reg min_dist_index_out_ap_vld;

(* fsm_encoding = "none" *) reg   [1:0] ap_CS_fsm;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter2;
reg    ap_idle_pp0;
wire    ap_CS_fsm_pp0_stage1;
wire    ap_block_state2_pp0_stage1_iter0;
wire    ap_block_state4_pp0_stage1_iter1;
wire    ap_block_state6_pp0_stage1_iter2;
wire    ap_block_pp0_stage1_subdone;
reg   [0:0] icmp_ln73_reg_408;
reg    ap_condition_exit_pp0_iter0_stage1;
wire    ap_loop_exit_ready;
reg    ap_ready_int;
reg  signed [63:0] cond68_reg_169;
reg  signed [63:0] cond87_reg_179;
wire    ap_block_state1_pp0_stage0_iter0;
wire    ap_block_state3_pp0_stage0_iter1;
wire    ap_block_state5_pp0_stage0_iter2;
wire    ap_block_pp0_stage0_11001;
reg   [12:0] node_x_coords_addr_reg_391;
reg   [12:0] node_y_coords_addr_reg_397;
wire   [31:0] j_cast_fu_219_p1;
reg   [31:0] j_cast_reg_403;
reg   [31:0] j_cast_reg_403_pp0_iter1_reg;
reg   [31:0] j_cast_reg_403_pp0_iter2_reg;
wire   [0:0] icmp_ln73_fu_223_p2;
reg   [0:0] icmp_ln73_reg_408_pp0_iter1_reg;
reg   [7:0] centroid_x_coords_addr_reg_412;
reg   [7:0] centroid_y_coords_addr_reg_418;
wire   [0:0] icmp_ln77_fu_240_p2;
reg   [0:0] icmp_ln77_reg_424;
wire    ap_block_pp0_stage1_11001;
wire   [0:0] icmp_ln79_fu_246_p2;
reg   [0:0] icmp_ln79_reg_428;
wire   [0:0] icmp_ln81_fu_252_p2;
reg   [0:0] icmp_ln81_reg_432;
wire   [0:0] icmp_ln83_fu_258_p2;
reg   [0:0] icmp_ln83_reg_436;
wire   [63:0] sub_ln79_fu_264_p2;
wire   [63:0] sub_ln78_fu_270_p2;
wire   [63:0] sub_ln81_fu_276_p2;
wire   [63:0] sub_ln80_fu_282_p2;
wire   [63:0] sub_ln83_fu_288_p2;
wire   [63:0] sub_ln82_fu_294_p2;
wire   [63:0] sub_ln85_fu_300_p2;
wire   [63:0] sub_ln84_fu_306_p2;
wire   [63:0] mul_ln79_fu_312_p2;
reg   [63:0] mul_ln79_reg_480;
wire   [63:0] mul_ln83_fu_318_p2;
reg   [63:0] mul_ln83_reg_485;
reg    ap_enable_reg_pp0_iter0_reg;
wire  signed [63:0] ap_phi_reg_pp0_iter0_cond_reg_151;
reg  signed [63:0] ap_phi_reg_pp0_iter1_cond_reg_151;
wire  signed [63:0] ap_phi_reg_pp0_iter0_cond48_reg_160;
reg  signed [63:0] ap_phi_reg_pp0_iter1_cond48_reg_160;
wire  signed [63:0] ap_phi_reg_pp0_iter0_cond68_reg_169;
reg  signed [63:0] ap_phi_reg_pp0_iter1_cond68_reg_169;
wire  signed [63:0] ap_phi_reg_pp0_iter0_cond87_reg_179;
reg  signed [63:0] ap_phi_reg_pp0_iter1_cond87_reg_179;
wire   [63:0] zext_ln69_cast_fu_189_p1;
wire    ap_block_pp0_stage0;
wire   [63:0] trunc_ln87_cast_fu_229_p1;
reg   [31:0] min_dist_index_fu_48;
wire   [31:0] min_dist_index_1_fu_340_p3;
wire    ap_block_pp0_stage1;
wire    ap_loop_init;
reg   [63:0] min_dist_fu_52;
wire   [63:0] min_dist_1_fu_347_p3;
reg   [30:0] j_fu_56;
wire   [30:0] add_ln73_fu_213_p2;
reg   [30:0] ap_sig_allocacmp_j_1;
wire    ap_block_pp0_stage1_01001;
wire   [63:0] centroid_dist_fu_330_p2;
wire   [0:0] icmp_ln87_fu_334_p2;
reg    ap_done_reg;
wire    ap_continue_int;
reg    ap_done_int;
reg    ap_loop_exit_ready_pp0_iter1_reg;
reg   [1:0] ap_NS_fsm;
wire    ap_block_pp0_stage0_subdone;
reg    ap_idle_pp0_1to2;
reg    ap_done_pending_pp0;
wire    ap_enable_pp0;
wire    ap_start_int;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_CS_fsm = 2'd1;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter0_reg = 1'b0;
#0 ap_done_reg = 1'b0;
end

kmeans_top_mul_64s_64s_64_1_1 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 64 ),
    .din1_WIDTH( 64 ),
    .dout_WIDTH( 64 ))
mul_64s_64s_64_1_1_U30(
    .din0(ap_phi_reg_pp0_iter1_cond48_reg_160),
    .din1(ap_phi_reg_pp0_iter1_cond_reg_151),
    .dout(mul_ln79_fu_312_p2)
);

kmeans_top_mul_64s_64s_64_1_1 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 64 ),
    .din1_WIDTH( 64 ),
    .dout_WIDTH( 64 ))
mul_64s_64s_64_1_1_U31(
    .din0(cond87_reg_179),
    .din1(cond68_reg_169),
    .dout(mul_ln83_fu_318_p2)
);

kmeans_top_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(ap_start),
    .ap_ready(ap_ready),
    .ap_done(ap_done),
    .ap_start_int(ap_start_int),
    .ap_loop_init(ap_loop_init),
    .ap_ready_int(ap_ready_int),
    .ap_loop_exit_ready(ap_condition_exit_pp0_iter0_stage1),
    .ap_loop_exit_done(ap_done_int),
    .ap_continue_int(ap_continue_int),
    .ap_done_int(ap_done_int)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue_int == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((ap_loop_exit_ready_pp0_iter1_reg == 1'b1) & (1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0_reg <= 1'b0;
    end else begin
        if ((1'b1 == ap_CS_fsm_pp0_stage0)) begin
            ap_enable_reg_pp0_iter0_reg <= ap_start_int;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b1 == ap_condition_exit_pp0_iter0_stage1)) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln73_reg_408 == 1'd1) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln79_reg_428 == 1'd0))) begin
        ap_phi_reg_pp0_iter1_cond48_reg_160 <= sub_ln81_fu_276_p2;
    end else if (((icmp_ln73_reg_408 == 1'd1) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln79_reg_428 == 1'd1))) begin
        ap_phi_reg_pp0_iter1_cond48_reg_160 <= sub_ln80_fu_282_p2;
    end else if (((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
        ap_phi_reg_pp0_iter1_cond48_reg_160 <= ap_phi_reg_pp0_iter0_cond48_reg_160;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln73_reg_408 == 1'd1) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln81_reg_432 == 1'd0))) begin
        ap_phi_reg_pp0_iter1_cond68_reg_169 <= sub_ln83_fu_288_p2;
    end else if (((icmp_ln73_reg_408 == 1'd1) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln81_reg_432 == 1'd1))) begin
        ap_phi_reg_pp0_iter1_cond68_reg_169 <= sub_ln82_fu_294_p2;
    end else if (((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
        ap_phi_reg_pp0_iter1_cond68_reg_169 <= ap_phi_reg_pp0_iter0_cond68_reg_169;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln73_reg_408 == 1'd1) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln83_reg_436 == 1'd0))) begin
        ap_phi_reg_pp0_iter1_cond87_reg_179 <= sub_ln85_fu_300_p2;
    end else if (((icmp_ln73_reg_408 == 1'd1) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln83_reg_436 == 1'd1))) begin
        ap_phi_reg_pp0_iter1_cond87_reg_179 <= sub_ln84_fu_306_p2;
    end else if (((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
        ap_phi_reg_pp0_iter1_cond87_reg_179 <= ap_phi_reg_pp0_iter0_cond87_reg_179;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln73_reg_408 == 1'd1) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln77_reg_424 == 1'd0))) begin
        ap_phi_reg_pp0_iter1_cond_reg_151 <= sub_ln79_fu_264_p2;
    end else if (((icmp_ln73_reg_408 == 1'd1) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln77_reg_424 == 1'd1))) begin
        ap_phi_reg_pp0_iter1_cond_reg_151 <= sub_ln78_fu_270_p2;
    end else if (((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
        ap_phi_reg_pp0_iter1_cond_reg_151 <= ap_phi_reg_pp0_iter0_cond_reg_151;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        if (((ap_enable_reg_pp0_iter0 == 1'b1) & (icmp_ln73_fu_223_p2 == 1'd1))) begin
            j_fu_56 <= add_ln73_fu_213_p2;
        end else if ((ap_loop_init == 1'b1)) begin
            j_fu_56 <= 31'd0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_loop_init == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        min_dist_fu_52 <= 64'd18446744073709551615;
    end else if (((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
        min_dist_fu_52 <= min_dist_1_fu_347_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_loop_init == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        min_dist_index_fu_48 <= 32'd0;
    end else if (((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter2 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
        min_dist_index_fu_48 <= min_dist_index_1_fu_340_p3;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
        ap_loop_exit_ready_pp0_iter1_reg <= ap_loop_exit_ready;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln73_fu_223_p2 == 1'd1))) begin
        centroid_x_coords_addr_reg_412 <= trunc_ln87_cast_fu_229_p1;
        centroid_y_coords_addr_reg_418 <= trunc_ln87_cast_fu_229_p1;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
        cond68_reg_169 <= ap_phi_reg_pp0_iter1_cond68_reg_169;
        cond87_reg_179 <= ap_phi_reg_pp0_iter1_cond87_reg_179;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        icmp_ln73_reg_408 <= icmp_ln73_fu_223_p2;
        icmp_ln73_reg_408_pp0_iter1_reg <= icmp_ln73_reg_408;
        j_cast_reg_403[30 : 0] <= j_cast_fu_219_p1[30 : 0];
        j_cast_reg_403_pp0_iter1_reg[30 : 0] <= j_cast_reg_403[30 : 0];
        j_cast_reg_403_pp0_iter2_reg[30 : 0] <= j_cast_reg_403_pp0_iter1_reg[30 : 0];
        mul_ln83_reg_485 <= mul_ln83_fu_318_p2;
        node_x_coords_addr_reg_391 <= zext_ln69_cast_fu_189_p1;
        node_y_coords_addr_reg_397 <= zext_ln69_cast_fu_189_p1;
    end
end

always @ (posedge ap_clk) begin
    if (((icmp_ln73_reg_408 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
        icmp_ln77_reg_424 <= icmp_ln77_fu_240_p2;
        icmp_ln79_reg_428 <= icmp_ln79_fu_246_p2;
        icmp_ln81_reg_432 <= icmp_ln81_fu_252_p2;
        icmp_ln83_reg_436 <= icmp_ln83_fu_258_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln73_reg_408_pp0_iter1_reg == 1'd1))) begin
        mul_ln79_reg_480 <= mul_ln79_fu_312_p2;
    end
end

always @ (*) begin
    if (((icmp_ln73_reg_408 == 1'd0) & (1'b0 == ap_block_pp0_stage1_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
        ap_condition_exit_pp0_iter0_stage1 = 1'b1;
    end else begin
        ap_condition_exit_pp0_iter0_stage1 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_loop_exit_ready_pp0_iter1_reg == 1'b1) & (1'b0 == ap_block_pp0_stage1_subdone) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
        ap_done_int = 1'b1;
    end else begin
        ap_done_int = ap_done_reg;
    end
end

always @ (*) begin
    if (~((ap_loop_exit_ready == 1'b0) & (ap_loop_exit_ready_pp0_iter1_reg == 1'b0))) begin
        ap_done_pending_pp0 = 1'b1;
    end else begin
        ap_done_pending_pp0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_pp0_stage0)) begin
        ap_enable_reg_pp0_iter0 = ap_start_int;
    end else begin
        ap_enable_reg_pp0_iter0 = ap_enable_reg_pp0_iter0_reg;
    end
end

always @ (*) begin
    if (((ap_start_int == 1'b0) & (ap_idle_pp0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0))) begin
        ap_idle_pp0_1to2 = 1'b1;
    end else begin
        ap_idle_pp0_1to2 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage1_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
        ap_ready_int = 1'b1;
    end else begin
        ap_ready_int = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (ap_loop_init == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_sig_allocacmp_j_1 = 31'd0;
    end else begin
        ap_sig_allocacmp_j_1 = j_fu_56;
    end
end

always @ (*) begin
    if ((((icmp_ln73_reg_408 == 1'd1) & (1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln79_fu_246_p2 == 1'd1)) | ((icmp_ln73_reg_408 == 1'd1) & (1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln79_fu_246_p2 == 1'd0)))) begin
        centroid_x_coords_address0 = centroid_x_coords_addr_reg_412;
    end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        centroid_x_coords_address0 = trunc_ln87_cast_fu_229_p1;
    end else begin
        centroid_x_coords_address0 = 'bx;
    end
end

always @ (*) begin
    if ((((icmp_ln73_reg_408 == 1'd1) & (1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln77_fu_240_p2 == 1'd1)) | ((icmp_ln73_reg_408 == 1'd1) & (1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln77_fu_240_p2 == 1'd0)))) begin
        centroid_x_coords_address1 = centroid_x_coords_addr_reg_412;
    end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        centroid_x_coords_address1 = trunc_ln87_cast_fu_229_p1;
    end else begin
        centroid_x_coords_address1 = 'bx;
    end
end

always @ (*) begin
    if ((((icmp_ln73_reg_408 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln79_fu_246_p2 == 1'd1)) | ((icmp_ln73_reg_408 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln79_fu_246_p2 == 1'd0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        centroid_x_coords_ce0 = 1'b1;
    end else begin
        centroid_x_coords_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((icmp_ln73_reg_408 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln77_fu_240_p2 == 1'd1)) | ((icmp_ln73_reg_408 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln77_fu_240_p2 == 1'd0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        centroid_x_coords_ce1 = 1'b1;
    end else begin
        centroid_x_coords_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((((icmp_ln73_reg_408 == 1'd1) & (1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln83_fu_258_p2 == 1'd1)) | ((icmp_ln73_reg_408 == 1'd1) & (1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln83_fu_258_p2 == 1'd0)))) begin
        centroid_y_coords_address0 = centroid_y_coords_addr_reg_418;
    end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        centroid_y_coords_address0 = trunc_ln87_cast_fu_229_p1;
    end else begin
        centroid_y_coords_address0 = 'bx;
    end
end

always @ (*) begin
    if ((((icmp_ln73_reg_408 == 1'd1) & (1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln81_fu_252_p2 == 1'd1)) | ((icmp_ln73_reg_408 == 1'd1) & (1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln81_fu_252_p2 == 1'd0)))) begin
        centroid_y_coords_address1 = centroid_y_coords_addr_reg_418;
    end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        centroid_y_coords_address1 = trunc_ln87_cast_fu_229_p1;
    end else begin
        centroid_y_coords_address1 = 'bx;
    end
end

always @ (*) begin
    if ((((icmp_ln73_reg_408 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln83_fu_258_p2 == 1'd1)) | ((icmp_ln73_reg_408 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln83_fu_258_p2 == 1'd0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        centroid_y_coords_ce0 = 1'b1;
    end else begin
        centroid_y_coords_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((icmp_ln73_reg_408 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln81_fu_252_p2 == 1'd1)) | ((icmp_ln73_reg_408 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln81_fu_252_p2 == 1'd0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        centroid_y_coords_ce1 = 1'b1;
    end else begin
        centroid_y_coords_ce1 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln73_reg_408_pp0_iter1_reg == 1'd0))) begin
        min_dist_index_out_ap_vld = 1'b1;
    end else begin
        min_dist_index_out_ap_vld = 1'b0;
    end
end

always @ (*) begin
    if ((((icmp_ln73_reg_408 == 1'd1) & (1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln79_fu_246_p2 == 1'd1)) | ((icmp_ln73_reg_408 == 1'd1) & (1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln79_fu_246_p2 == 1'd0)))) begin
        node_x_coords_address0 = node_x_coords_addr_reg_391;
    end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        node_x_coords_address0 = zext_ln69_cast_fu_189_p1;
    end else begin
        node_x_coords_address0 = 'bx;
    end
end

always @ (*) begin
    if ((((icmp_ln73_reg_408 == 1'd1) & (1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln77_fu_240_p2 == 1'd1)) | ((icmp_ln73_reg_408 == 1'd1) & (1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln77_fu_240_p2 == 1'd0)))) begin
        node_x_coords_address1 = node_x_coords_addr_reg_391;
    end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        node_x_coords_address1 = zext_ln69_cast_fu_189_p1;
    end else begin
        node_x_coords_address1 = 'bx;
    end
end

always @ (*) begin
    if ((((icmp_ln73_reg_408 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln79_fu_246_p2 == 1'd1)) | ((icmp_ln73_reg_408 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln79_fu_246_p2 == 1'd0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        node_x_coords_ce0 = 1'b1;
    end else begin
        node_x_coords_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((icmp_ln73_reg_408 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln77_fu_240_p2 == 1'd1)) | ((icmp_ln73_reg_408 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln77_fu_240_p2 == 1'd0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        node_x_coords_ce1 = 1'b1;
    end else begin
        node_x_coords_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((((icmp_ln73_reg_408 == 1'd1) & (1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln83_fu_258_p2 == 1'd1)) | ((icmp_ln73_reg_408 == 1'd1) & (1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln83_fu_258_p2 == 1'd0)))) begin
        node_y_coords_address0 = node_y_coords_addr_reg_397;
    end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        node_y_coords_address0 = zext_ln69_cast_fu_189_p1;
    end else begin
        node_y_coords_address0 = 'bx;
    end
end

always @ (*) begin
    if ((((icmp_ln73_reg_408 == 1'd1) & (1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln81_fu_252_p2 == 1'd1)) | ((icmp_ln73_reg_408 == 1'd1) & (1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln81_fu_252_p2 == 1'd0)))) begin
        node_y_coords_address1 = node_y_coords_addr_reg_397;
    end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        node_y_coords_address1 = zext_ln69_cast_fu_189_p1;
    end else begin
        node_y_coords_address1 = 'bx;
    end
end

always @ (*) begin
    if ((((icmp_ln73_reg_408 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln83_fu_258_p2 == 1'd1)) | ((icmp_ln73_reg_408 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln83_fu_258_p2 == 1'd0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        node_y_coords_ce0 = 1'b1;
    end else begin
        node_y_coords_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((((icmp_ln73_reg_408 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln81_fu_252_p2 == 1'd1)) | ((icmp_ln73_reg_408 == 1'd1) & (1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (icmp_ln81_fu_252_p2 == 1'd0)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        node_y_coords_ce1 = 1'b1;
    end else begin
        node_y_coords_ce1 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((ap_start_int == 1'b0) & (ap_done_pending_pp0 == 1'b0) & (ap_idle_pp0_1to2 == 1'b1)) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_pp0_stage1 : begin
            if ((1'b0 == ap_block_pp0_stage1_subdone)) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign add_ln73_fu_213_p2 = (ap_sig_allocacmp_j_1 + 31'd1);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_pp0_stage1 = ap_CS_fsm[32'd1];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_01001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_subdone = ~(1'b1 == 1'b1);

assign ap_block_state1_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage1_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state4_pp0_stage1_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state5_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_block_state6_pp0_stage1_iter2 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_loop_exit_ready = ap_condition_exit_pp0_iter0_stage1;

assign ap_phi_reg_pp0_iter0_cond48_reg_160 = 'bx;

assign ap_phi_reg_pp0_iter0_cond68_reg_169 = 'bx;

assign ap_phi_reg_pp0_iter0_cond87_reg_179 = 'bx;

assign ap_phi_reg_pp0_iter0_cond_reg_151 = 'bx;

assign centroid_dist_fu_330_p2 = (mul_ln83_reg_485 + mul_ln79_reg_480);

assign icmp_ln73_fu_223_p2 = (($signed(j_cast_fu_219_p1) < $signed(k)) ? 1'b1 : 1'b0);

assign icmp_ln77_fu_240_p2 = ((node_x_coords_q1 < centroid_x_coords_q1) ? 1'b1 : 1'b0);

assign icmp_ln79_fu_246_p2 = ((node_x_coords_q0 < centroid_x_coords_q0) ? 1'b1 : 1'b0);

assign icmp_ln81_fu_252_p2 = ((node_y_coords_q1 < centroid_y_coords_q1) ? 1'b1 : 1'b0);

assign icmp_ln83_fu_258_p2 = ((node_y_coords_q0 < centroid_y_coords_q0) ? 1'b1 : 1'b0);

assign icmp_ln87_fu_334_p2 = ((centroid_dist_fu_330_p2 < min_dist_fu_52) ? 1'b1 : 1'b0);

assign j_cast_fu_219_p1 = ap_sig_allocacmp_j_1;

assign min_dist_1_fu_347_p3 = ((icmp_ln87_fu_334_p2[0:0] == 1'b1) ? centroid_dist_fu_330_p2 : min_dist_fu_52);

assign min_dist_index_1_fu_340_p3 = ((icmp_ln87_fu_334_p2[0:0] == 1'b1) ? j_cast_reg_403_pp0_iter2_reg : min_dist_index_fu_48);

assign min_dist_index_out = min_dist_index_fu_48;

assign sub_ln78_fu_270_p2 = (centroid_x_coords_q1 - node_x_coords_q1);

assign sub_ln79_fu_264_p2 = (node_x_coords_q1 - centroid_x_coords_q1);

assign sub_ln80_fu_282_p2 = (centroid_x_coords_q0 - node_x_coords_q0);

assign sub_ln81_fu_276_p2 = (node_x_coords_q0 - centroid_x_coords_q0);

assign sub_ln82_fu_294_p2 = (centroid_y_coords_q1 - node_y_coords_q1);

assign sub_ln83_fu_288_p2 = (node_y_coords_q1 - centroid_y_coords_q1);

assign sub_ln84_fu_306_p2 = (centroid_y_coords_q0 - node_y_coords_q0);

assign sub_ln85_fu_300_p2 = (node_y_coords_q0 - centroid_y_coords_q0);

assign trunc_ln87_cast_fu_229_p1 = ap_sig_allocacmp_j_1;

assign zext_ln69_cast_fu_189_p1 = zext_ln69;

always @ (posedge ap_clk) begin
    j_cast_reg_403[31] <= 1'b0;
    j_cast_reg_403_pp0_iter1_reg[31] <= 1'b0;
    j_cast_reg_403_pp0_iter2_reg[31] <= 1'b0;
end

endmodule //kmeans_top_kmeans_Pipeline_VITIS_LOOP_73_3


// Content from kmeans_top_kmeans_Pipeline_1.v
// ==============================================================
// RTL generated by Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2022.2 (64-bit)
// Version: 2022.2
// Copyright (C) Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// 
// ===========================================================

`timescale 1 ns / 1 ps 

module kmeans_top_kmeans_Pipeline_1 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        centroid_x_coords_address0,
        centroid_x_coords_ce0,
        centroid_x_coords_q0,
        centroid_x_coords_prev_address0,
        centroid_x_coords_prev_ce0,
        centroid_x_coords_prev_we0,
        centroid_x_coords_prev_d0,
        p_cast12
);

parameter    ap_ST_fsm_pp0_stage0 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
output  [7:0] centroid_x_coords_address0;
output   centroid_x_coords_ce0;
input  [63:0] centroid_x_coords_q0;
output  [7:0] centroid_x_coords_prev_address0;
output   centroid_x_coords_prev_ce0;
output   centroid_x_coords_prev_we0;
output  [63:0] centroid_x_coords_prev_d0;
input  [31:0] p_cast12;

reg ap_idle;
reg centroid_x_coords_ce0;
reg centroid_x_coords_prev_ce0;
reg centroid_x_coords_prev_we0;

(* fsm_encoding = "none" *) reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_enable_reg_pp0_iter0;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter2;
reg    ap_idle_pp0;
wire    ap_block_state1_pp0_stage0_iter0;
wire    ap_block_state2_pp0_stage0_iter1;
wire    ap_block_state3_pp0_stage0_iter2;
wire    ap_block_pp0_stage0_subdone;
wire   [0:0] exitcond_fu_90_p2;
reg    ap_condition_exit_pp0_iter1_stage0;
wire    ap_loop_exit_ready;
reg    ap_ready_int;
wire  signed [60:0] p_cast12_cast_fu_67_p1;
reg  signed [60:0] p_cast12_cast_reg_107;
wire    ap_block_pp0_stage0_11001;
wire   [63:0] loop_index_cast_fu_85_p1;
reg   [63:0] loop_index_cast_reg_112;
wire    ap_block_pp0_stage0;
reg   [60:0] loop_index_fu_30;
wire   [60:0] empty_fu_79_p2;
wire    ap_loop_init;
reg    ap_done_reg;
wire    ap_continue_int;
reg    ap_done_int;
reg    ap_loop_exit_ready_pp0_iter2_reg;
reg   [0:0] ap_NS_fsm;
wire    ap_enable_pp0;
wire    ap_start_int;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_CS_fsm = 1'd1;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_done_reg = 1'b0;
end

kmeans_top_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(ap_start),
    .ap_ready(ap_ready),
    .ap_done(ap_done),
    .ap_start_int(ap_start_int),
    .ap_loop_init(ap_loop_init),
    .ap_ready_int(ap_ready_int),
    .ap_loop_exit_ready(ap_condition_exit_pp0_iter1_stage0),
    .ap_loop_exit_done(ap_done_int),
    .ap_continue_int(ap_continue_int),
    .ap_done_int(ap_done_int)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue_int == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter2_reg == 1'b1))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b1 == ap_condition_exit_pp0_iter1_stage0)) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_enable_reg_pp0_iter1 <= ap_start_int;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((ap_loop_exit_ready == 1'b0) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
        ap_loop_exit_ready_pp0_iter2_reg <= 1'b0;
    end else if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_loop_exit_ready_pp0_iter2_reg <= ap_loop_exit_ready;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        if ((ap_loop_init == 1'b1)) begin
            loop_index_fu_30 <= 61'd0;
        end else if (((exitcond_fu_90_p2 == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
            loop_index_fu_30 <= empty_fu_79_p2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        loop_index_cast_reg_112[60 : 0] <= loop_index_cast_fu_85_p1[60 : 0];
        p_cast12_cast_reg_107 <= p_cast12_cast_fu_67_p1;
    end
end

always @ (*) begin
    if (((exitcond_fu_90_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_condition_exit_pp0_iter1_stage0 = 1'b1;
    end else begin
        ap_condition_exit_pp0_iter1_stage0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter2_reg == 1'b1))) begin
        ap_done_int = 1'b1;
    end else begin
        ap_done_int = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_idle_pp0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_start_int == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_ready_int = 1'b1;
    end else begin
        ap_ready_int = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        centroid_x_coords_ce0 = 1'b1;
    end else begin
        centroid_x_coords_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        centroid_x_coords_prev_ce0 = 1'b1;
    end else begin
        centroid_x_coords_prev_ce0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        centroid_x_coords_prev_we0 = 1'b1;
    end else begin
        centroid_x_coords_prev_we0 = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_pp0_stage0 : begin
            ap_NS_fsm = ap_ST_fsm_pp0_stage0;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

assign ap_block_state1_pp0_stage0_iter0 = ~(1'b1 == 1'b1);

assign ap_block_state2_pp0_stage0_iter1 = ~(1'b1 == 1'b1);

assign ap_block_state3_pp0_stage0_iter2 = ~(1'b1 == 1'b1);

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_enable_reg_pp0_iter0 = ap_start_int;

assign ap_loop_exit_ready = ap_condition_exit_pp0_iter1_stage0;

assign centroid_x_coords_address0 = loop_index_cast_fu_85_p1;

assign centroid_x_coords_prev_address0 = loop_index_cast_reg_112;

assign centroid_x_coords_prev_d0 = centroid_x_coords_q0;

assign empty_fu_79_p2 = (loop_index_fu_30 + 61'd1);

assign exitcond_fu_90_p2 = ((empty_fu_79_p2 == p_cast12_cast_reg_107) ? 1'b1 : 1'b0);

assign loop_index_cast_fu_85_p1 = loop_index_fu_30;

assign p_cast12_cast_fu_67_p1 = $signed(p_cast12);

always @ (posedge ap_clk) begin
    loop_index_cast_reg_112[63:61] <= 3'b000;
end

endmodule //kmeans_top_kmeans_Pipeline_1


// Content from kmeans_top_centroid_x_coords_RAM_1WNR_AUTO_1R1W.v
// ==============================================================
// Vitis HLS - High-Level Synthesis from C, C++ and OpenCL v2022.2 (64-bit)
// Version: 2022.2
// Copyright 1986-2022 Xilinx, Inc. All Rights Reserved.
// ==============================================================
`timescale 1 ns / 1 ps
module kmeans_top_centroid_x_coords_RAM_1WNR_AUTO_1R1W (
     
    address0, ce0,
    d0, we0, 
    q0, 
     
    address1, ce1,
    
    q1, 
    
    reset, clk);

parameter DataWidth = 64;
parameter AddressWidth = 8;
parameter AddressRange = 256;

input[AddressWidth-1:0] address0;
input ce0;
input[DataWidth-1:0] d0;
input we0; 
output reg[DataWidth-1:0] q0; 

input[AddressWidth-1:0] address1;
input ce1;

output reg[DataWidth-1:0] q1; 

input reset;
input clk;


(* ram_style = "auto"  *)reg [DataWidth-1:0] ram0[0:AddressRange-1];


 


// write to all ram
always @(posedge clk)  
begin 
    if (ce0) begin
        if (we0) 
            ram0[address0] <= d0; 

        q0 <= ram0[address0]; 
    end
end

always @(posedge clk)  
begin 
    if (ce1) begin
        q1 <= ram0[address1];
    end
end


endmodule





// Content from axi_interconnect_wrap_2x1.v
/*

Copyright (c) 2020 Alex Forencich

Permission is hereby granted, free of charge, to any person obtaining a copy
of this software and associated documentation files (the "Software"), to deal
in the Software without restriction, including without limitation the rights
to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
copies of the Software, and to permit persons to whom the Software is
furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in
all copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY
FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
THE SOFTWARE.

*/

// Language: Verilog 2001

/*
 * AXI4 2x1 interconnect (wrapper)
 */
module axi_interconnect_wrap_2x1 #
(
    parameter DATA_WIDTH = 32,
    parameter ADDR_WIDTH = 32,
    parameter STRB_WIDTH = (DATA_WIDTH/8),
    parameter ID_WIDTH = 8,
    parameter AWUSER_ENABLE = 0,
    parameter AWUSER_WIDTH = 1,
    parameter WUSER_ENABLE = 0,
    parameter WUSER_WIDTH = 1,
    parameter BUSER_ENABLE = 0,
    parameter BUSER_WIDTH = 1,
    parameter ARUSER_ENABLE = 0,
    parameter ARUSER_WIDTH = 1,
    parameter RUSER_ENABLE = 0,
    parameter RUSER_WIDTH = 1,
    parameter FORWARD_ID = 0,
    parameter M_REGIONS = 1,
    parameter M00_BASE_ADDR = 0,
    parameter M00_ADDR_WIDTH = {M_REGIONS{32'd24}},
    parameter M00_CONNECT_READ = 2'b11,
    parameter M00_CONNECT_WRITE = 2'b11,
    parameter M00_SECURE = 1'b0
)
(
    input  wire                     clk,
    input  wire                     rst,

    /*
     * AXI slave interface
     */
    input  wire [ID_WIDTH-1:0]      s00_axi_awid,
    input  wire [ADDR_WIDTH-1:0]    s00_axi_awaddr,
    input  wire [7:0]               s00_axi_awlen,
    input  wire [2:0]               s00_axi_awsize,
    input  wire [1:0]               s00_axi_awburst,
    input  wire                     s00_axi_awlock,
    input  wire [3:0]               s00_axi_awcache,
    input  wire [2:0]               s00_axi_awprot,
    input  wire [3:0]               s00_axi_awqos,
    input  wire [AWUSER_WIDTH-1:0]  s00_axi_awuser,
    input  wire                     s00_axi_awvalid,
    output wire                     s00_axi_awready,
    input  wire [DATA_WIDTH-1:0]    s00_axi_wdata,
    input  wire [STRB_WIDTH-1:0]    s00_axi_wstrb,
    input  wire                     s00_axi_wlast,
    input  wire [WUSER_WIDTH-1:0]   s00_axi_wuser,
    input  wire                     s00_axi_wvalid,
    output wire                     s00_axi_wready,
    output wire [ID_WIDTH-1:0]      s00_axi_bid,
    output wire [1:0]               s00_axi_bresp,
    output wire [BUSER_WIDTH-1:0]   s00_axi_buser,
    output wire                     s00_axi_bvalid,
    input  wire                     s00_axi_bready,
    input  wire [ID_WIDTH-1:0]      s00_axi_arid,
    input  wire [ADDR_WIDTH-1:0]    s00_axi_araddr,
    input  wire [7:0]               s00_axi_arlen,
    input  wire [2:0]               s00_axi_arsize,
    input  wire [1:0]               s00_axi_arburst,
    input  wire                     s00_axi_arlock,
    input  wire [3:0]               s00_axi_arcache,
    input  wire [2:0]               s00_axi_arprot,
    input  wire [3:0]               s00_axi_arqos,
    input  wire [ARUSER_WIDTH-1:0]  s00_axi_aruser,
    input  wire                     s00_axi_arvalid,
    output wire                     s00_axi_arready,
    output wire [ID_WIDTH-1:0]      s00_axi_rid,
    output wire [DATA_WIDTH-1:0]    s00_axi_rdata,
    output wire [1:0]               s00_axi_rresp,
    output wire                     s00_axi_rlast,
    output wire [RUSER_WIDTH-1:0]   s00_axi_ruser,
    output wire                     s00_axi_rvalid,
    input  wire                     s00_axi_rready,

    input  wire [ID_WIDTH-1:0]      s01_axi_awid,
    input  wire [ADDR_WIDTH-1:0]    s01_axi_awaddr,
    input  wire [7:0]               s01_axi_awlen,
    input  wire [2:0]               s01_axi_awsize,
    input  wire [1:0]               s01_axi_awburst,
    input  wire                     s01_axi_awlock,
    input  wire [3:0]               s01_axi_awcache,
    input  wire [2:0]               s01_axi_awprot,
    input  wire [3:0]               s01_axi_awqos,
    input  wire [AWUSER_WIDTH-1:0]  s01_axi_awuser,
    input  wire                     s01_axi_awvalid,
    output wire                     s01_axi_awready,
    input  wire [DATA_WIDTH-1:0]    s01_axi_wdata,
    input  wire [STRB_WIDTH-1:0]    s01_axi_wstrb,
    input  wire                     s01_axi_wlast,
    input  wire [WUSER_WIDTH-1:0]   s01_axi_wuser,
    input  wire                     s01_axi_wvalid,
    output wire                     s01_axi_wready,
    output wire [ID_WIDTH-1:0]      s01_axi_bid,
    output wire [1:0]               s01_axi_bresp,
    output wire [BUSER_WIDTH-1:0]   s01_axi_buser,
    output wire                     s01_axi_bvalid,
    input  wire                     s01_axi_bready,
    input  wire [ID_WIDTH-1:0]      s01_axi_arid,
    input  wire [ADDR_WIDTH-1:0]    s01_axi_araddr,
    input  wire [7:0]               s01_axi_arlen,
    input  wire [2:0]               s01_axi_arsize,
    input  wire [1:0]               s01_axi_arburst,
    input  wire                     s01_axi_arlock,
    input  wire [3:0]               s01_axi_arcache,
    input  wire [2:0]               s01_axi_arprot,
    input  wire [3:0]               s01_axi_arqos,
    input  wire [ARUSER_WIDTH-1:0]  s01_axi_aruser,
    input  wire                     s01_axi_arvalid,
    output wire                     s01_axi_arready,
    output wire [ID_WIDTH-1:0]      s01_axi_rid,
    output wire [DATA_WIDTH-1:0]    s01_axi_rdata,
    output wire [1:0]               s01_axi_rresp,
    output wire                     s01_axi_rlast,
    output wire [RUSER_WIDTH-1:0]   s01_axi_ruser,
    output wire                     s01_axi_rvalid,
    input  wire                     s01_axi_rready,

    /*
     * AXI master interface
     */
    output wire [ID_WIDTH-1:0]      m00_axi_awid,
    output wire [ADDR_WIDTH-1:0]    m00_axi_awaddr,
    output wire [7:0]               m00_axi_awlen,
    output wire [2:0]               m00_axi_awsize,
    output wire [1:0]               m00_axi_awburst,
    output wire                     m00_axi_awlock,
    output wire [3:0]               m00_axi_awcache,
    output wire [2:0]               m00_axi_awprot,
    output wire [3:0]               m00_axi_awqos,
    output wire [3:0]               m00_axi_awregion,
    output wire [AWUSER_WIDTH-1:0]  m00_axi_awuser,
    output wire                     m00_axi_awvalid,
    input  wire                     m00_axi_awready,
    output wire [DATA_WIDTH-1:0]    m00_axi_wdata,
    output wire [STRB_WIDTH-1:0]    m00_axi_wstrb,
    output wire                     m00_axi_wlast,
    output wire [WUSER_WIDTH-1:0]   m00_axi_wuser,
    output wire                     m00_axi_wvalid,
    input  wire                     m00_axi_wready,
    input  wire [ID_WIDTH-1:0]      m00_axi_bid,
    input  wire [1:0]               m00_axi_bresp,
    input  wire [BUSER_WIDTH-1:0]   m00_axi_buser,
    input  wire                     m00_axi_bvalid,
    output wire                     m00_axi_bready,
    output wire [ID_WIDTH-1:0]      m00_axi_arid,
    output wire [ADDR_WIDTH-1:0]    m00_axi_araddr,
    output wire [7:0]               m00_axi_arlen,
    output wire [2:0]               m00_axi_arsize,
    output wire [1:0]               m00_axi_arburst,
    output wire                     m00_axi_arlock,
    output wire [3:0]               m00_axi_arcache,
    output wire [2:0]               m00_axi_arprot,
    output wire [3:0]               m00_axi_arqos,
    output wire [3:0]               m00_axi_arregion,
    output wire [ARUSER_WIDTH-1:0]  m00_axi_aruser,
    output wire                     m00_axi_arvalid,
    input  wire                     m00_axi_arready,
    input  wire [ID_WIDTH-1:0]      m00_axi_rid,
    input  wire [DATA_WIDTH-1:0]    m00_axi_rdata,
    input  wire [1:0]               m00_axi_rresp,
    input  wire                     m00_axi_rlast,
    input  wire [RUSER_WIDTH-1:0]   m00_axi_ruser,
    input  wire                     m00_axi_rvalid,
    output wire                     m00_axi_rready
);

localparam S_COUNT = 2;
localparam M_COUNT = 1;

// parameter sizing helpers
function [ADDR_WIDTH*M_REGIONS-1:0] w_a_r(input [ADDR_WIDTH*M_REGIONS-1:0] val);
    w_a_r = val;
endfunction

function [32*M_REGIONS-1:0] w_32_r(input [32*M_REGIONS-1:0] val);
    w_32_r = val;
endfunction

function [S_COUNT-1:0] w_s(input [S_COUNT-1:0] val);
    w_s = val;
endfunction

function w_1(input val);
    w_1 = val;
endfunction

axi_interconnect #(
    .S_COUNT(S_COUNT),
    .M_COUNT(M_COUNT),
    .DATA_WIDTH(DATA_WIDTH),
    .ADDR_WIDTH(ADDR_WIDTH),
    .STRB_WIDTH(STRB_WIDTH),
    .ID_WIDTH(ID_WIDTH),
    .AWUSER_ENABLE(AWUSER_ENABLE),
    .AWUSER_WIDTH(AWUSER_WIDTH),
    .WUSER_ENABLE(WUSER_ENABLE),
    .WUSER_WIDTH(WUSER_WIDTH),
    .BUSER_ENABLE(BUSER_ENABLE),
    .BUSER_WIDTH(BUSER_WIDTH),
    .ARUSER_ENABLE(ARUSER_ENABLE),
    .ARUSER_WIDTH(ARUSER_WIDTH),
    .RUSER_ENABLE(RUSER_ENABLE),
    .RUSER_WIDTH(RUSER_WIDTH),
    .FORWARD_ID(FORWARD_ID),
    .M_REGIONS(M_REGIONS),
    .M_BASE_ADDR({ w_a_r(M00_BASE_ADDR) }),
    .M_ADDR_WIDTH({ w_32_r(M00_ADDR_WIDTH) }),
    .M_CONNECT_READ({ w_s(M00_CONNECT_READ) }),
    .M_CONNECT_WRITE({ w_s(M00_CONNECT_WRITE) }),
    .M_SECURE({ w_1(M00_SECURE) })
)
axi_interconnect_inst (
    .clk(clk),
    .rst(rst),
    .s_axi_awid({ s01_axi_awid, s00_axi_awid }),
    .s_axi_awaddr({ s01_axi_awaddr, s00_axi_awaddr }),
    .s_axi_awlen({ s01_axi_awlen, s00_axi_awlen }),
    .s_axi_awsize({ s01_axi_awsize, s00_axi_awsize }),
    .s_axi_awburst({ s01_axi_awburst, s00_axi_awburst }),
    .s_axi_awlock({ s01_axi_awlock, s00_axi_awlock }),
    .s_axi_awcache({ s01_axi_awcache, s00_axi_awcache }),
    .s_axi_awprot({ s01_axi_awprot, s00_axi_awprot }),
    .s_axi_awqos({ s01_axi_awqos, s00_axi_awqos }),
    .s_axi_awuser({ s01_axi_awuser, s00_axi_awuser }),
    .s_axi_awvalid({ s01_axi_awvalid, s00_axi_awvalid }),
    .s_axi_awready({ s01_axi_awready, s00_axi_awready }),
    .s_axi_wdata({ s01_axi_wdata, s00_axi_wdata }),
    .s_axi_wstrb({ s01_axi_wstrb, s00_axi_wstrb }),
    .s_axi_wlast({ s01_axi_wlast, s00_axi_wlast }),
    .s_axi_wuser({ s01_axi_wuser, s00_axi_wuser }),
    .s_axi_wvalid({ s01_axi_wvalid, s00_axi_wvalid }),
    .s_axi_wready({ s01_axi_wready, s00_axi_wready }),
    .s_axi_bid({ s01_axi_bid, s00_axi_bid }),
    .s_axi_bresp({ s01_axi_bresp, s00_axi_bresp }),
    .s_axi_buser({ s01_axi_buser, s00_axi_buser }),
    .s_axi_bvalid({ s01_axi_bvalid, s00_axi_bvalid }),
    .s_axi_bready({ s01_axi_bready, s00_axi_bready }),
    .s_axi_arid({ s01_axi_arid, s00_axi_arid }),
    .s_axi_araddr({ s01_axi_araddr, s00_axi_araddr }),
    .s_axi_arlen({ s01_axi_arlen, s00_axi_arlen }),
    .s_axi_arsize({ s01_axi_arsize, s00_axi_arsize }),
    .s_axi_arburst({ s01_axi_arburst, s00_axi_arburst }),
    .s_axi_arlock({ s01_axi_arlock, s00_axi_arlock }),
    .s_axi_arcache({ s01_axi_arcache, s00_axi_arcache }),
    .s_axi_arprot({ s01_axi_arprot, s00_axi_arprot }),
    .s_axi_arqos({ s01_axi_arqos, s00_axi_arqos }),
    .s_axi_aruser({ s01_axi_aruser, s00_axi_aruser }),
    .s_axi_arvalid({ s01_axi_arvalid, s00_axi_arvalid }),
    .s_axi_arready({ s01_axi_arready, s00_axi_arready }),
    .s_axi_rid({ s01_axi_rid, s00_axi_rid }),
    .s_axi_rdata({ s01_axi_rdata, s00_axi_rdata }),
    .s_axi_rresp({ s01_axi_rresp, s00_axi_rresp }),
    .s_axi_rlast({ s01_axi_rlast, s00_axi_rlast }),
    .s_axi_ruser({ s01_axi_ruser, s00_axi_ruser }),
    .s_axi_rvalid({ s01_axi_rvalid, s00_axi_rvalid }),
    .s_axi_rready({ s01_axi_rready, s00_axi_rready }),
    .m_axi_awid({ m00_axi_awid }),
    .m_axi_awaddr({ m00_axi_awaddr }),
    .m_axi_awlen({ m00_axi_awlen }),
    .m_axi_awsize({ m00_axi_awsize }),
    .m_axi_awburst({ m00_axi_awburst }),
    .m_axi_awlock({ m00_axi_awlock }),
    .m_axi_awcache({ m00_axi_awcache }),
    .m_axi_awprot({ m00_axi_awprot }),
    .m_axi_awqos({ m00_axi_awqos }),
    .m_axi_awregion({ m00_axi_awregion }),
    .m_axi_awuser({ m00_axi_awuser }),
    .m_axi_awvalid({ m00_axi_awvalid }),
    .m_axi_awready({ m00_axi_awready }),
    .m_axi_wdata({ m00_axi_wdata }),
    .m_axi_wstrb({ m00_axi_wstrb }),
    .m_axi_wlast({ m00_axi_wlast }),
    .m_axi_wuser({ m00_axi_wuser }),
    .m_axi_wvalid({ m00_axi_wvalid }),
    .m_axi_wready({ m00_axi_wready }),
    .m_axi_bid({ m00_axi_bid }),
    .m_axi_bresp({ m00_axi_bresp }),
    .m_axi_buser({ m00_axi_buser }),
    .m_axi_bvalid({ m00_axi_bvalid }),
    .m_axi_bready({ m00_axi_bready }),
    .m_axi_arid({ m00_axi_arid }),
    .m_axi_araddr({ m00_axi_araddr }),
    .m_axi_arlen({ m00_axi_arlen }),
    .m_axi_arsize({ m00_axi_arsize }),
    .m_axi_arburst({ m00_axi_arburst }),
    .m_axi_arlock({ m00_axi_arlock }),
    .m_axi_arcache({ m00_axi_arcache }),
    .m_axi_arprot({ m00_axi_arprot }),
    .m_axi_arqos({ m00_axi_arqos }),
    .m_axi_arregion({ m00_axi_arregion }),
    .m_axi_aruser({ m00_axi_aruser }),
    .m_axi_arvalid({ m00_axi_arvalid }),
    .m_axi_arready({ m00_axi_arready }),
    .m_axi_rid({ m00_axi_rid }),
    .m_axi_rdata({ m00_axi_rdata }),
    .m_axi_rresp({ m00_axi_rresp }),
    .m_axi_rlast({ m00_axi_rlast }),
    .m_axi_ruser({ m00_axi_ruser }),
    .m_axi_rvalid({ m00_axi_rvalid }),
    .m_axi_rready({ m00_axi_rready })
);

endmodule

`resetall


// Content from arbiter.v
/*

Copyright (c) 2014-2021 Alex Forencich

Permission is hereby granted, free of charge, to any person obtaining a copy
of this software and associated documentation files (the "Software"), to deal
in the Software without restriction, including without limitation the rights
to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
copies of the Software, and to permit persons to whom the Software is
furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in
all copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY
FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
THE SOFTWARE.

*/

// Language: Verilog 2001


/*
 * Arbiter module
 */
module arbiter #
(
    parameter PORTS = 4,
    // select round robin arbitration
    parameter ARB_TYPE_ROUND_ROBIN = 0,
    // blocking arbiter enable
    parameter ARB_BLOCK = 0,
    // block on acknowledge assert when nonzero, request deassert when 0
    parameter ARB_BLOCK_ACK = 1,
    // LSB priority selection
    parameter ARB_LSB_HIGH_PRIORITY = 0
)
(
    input  wire                     clk,
    input  wire                     rst,

    input  wire [PORTS-1:0]         request,
    input  wire [PORTS-1:0]         acknowledge,

    output wire [PORTS-1:0]         grant,
    output wire                     grant_valid,
    output wire [$clog2(PORTS)-1:0] grant_encoded
);

reg [PORTS-1:0] grant_reg = 0, grant_next;
reg grant_valid_reg = 0, grant_valid_next;
reg [$clog2(PORTS)-1:0] grant_encoded_reg = 0, grant_encoded_next;

assign grant_valid = grant_valid_reg;
assign grant = grant_reg;
assign grant_encoded = grant_encoded_reg;

wire request_valid;
wire [$clog2(PORTS)-1:0] request_index;
wire [PORTS-1:0] request_mask;

priority_encoder #(
    .WIDTH(PORTS),
    .LSB_HIGH_PRIORITY(ARB_LSB_HIGH_PRIORITY)
)
priority_encoder_inst (
    .input_unencoded(request),
    .output_valid(request_valid),
    .output_encoded(request_index),
    .output_unencoded(request_mask)
);

reg [PORTS-1:0] mask_reg = 0, mask_next;

wire masked_request_valid;
wire [$clog2(PORTS)-1:0] masked_request_index;
wire [PORTS-1:0] masked_request_mask;

priority_encoder #(
    .WIDTH(PORTS),
    .LSB_HIGH_PRIORITY(ARB_LSB_HIGH_PRIORITY)
)
priority_encoder_masked (
    .input_unencoded(request & mask_reg),
    .output_valid(masked_request_valid),
    .output_encoded(masked_request_index),
    .output_unencoded(masked_request_mask)
);

always @* begin
    grant_next = 0;
    grant_valid_next = 0;
    grant_encoded_next = 0;
    mask_next = mask_reg;

    if (ARB_BLOCK && !ARB_BLOCK_ACK && grant_reg & request) begin
        // granted request still asserted; hold it
        grant_valid_next = grant_valid_reg;
        grant_next = grant_reg;
        grant_encoded_next = grant_encoded_reg;
    end else if (ARB_BLOCK && ARB_BLOCK_ACK && grant_valid && !(grant_reg & acknowledge)) begin
        // granted request not yet acknowledged; hold it
        grant_valid_next = grant_valid_reg;
        grant_next = grant_reg;
        grant_encoded_next = grant_encoded_reg;
    end else if (request_valid) begin
        if (ARB_TYPE_ROUND_ROBIN) begin
            if (masked_request_valid) begin
                grant_valid_next = 1;
                grant_next = masked_request_mask;
                grant_encoded_next = masked_request_index;
                if (ARB_LSB_HIGH_PRIORITY) begin
                    mask_next = {PORTS{1'b1}} << (masked_request_index + 1);
                end else begin
                    mask_next = {PORTS{1'b1}} >> (PORTS - masked_request_index);
                end
            end else begin
                grant_valid_next = 1;
                grant_next = request_mask;
                grant_encoded_next = request_index;
                if (ARB_LSB_HIGH_PRIORITY) begin
                    mask_next = {PORTS{1'b1}} << (request_index + 1);
                end else begin
                    mask_next = {PORTS{1'b1}} >> (PORTS - request_index);
                end
            end
        end else begin
            grant_valid_next = 1;
            grant_next = request_mask;
            grant_encoded_next = request_index;
        end
    end
end

always @(posedge clk) begin
    if (rst) begin
        grant_reg <= 0;
        grant_valid_reg <= 0;
        grant_encoded_reg <= 0;
        mask_reg <= 0;
    end else begin
        grant_reg <= grant_next;
        grant_valid_reg <= grant_valid_next;
        grant_encoded_reg <= grant_encoded_next;
        mask_reg <= mask_next;
    end
end

endmodule

`resetall


