/*
 * This header file provides definitions for ch_intrinsic_modified.v
 * located at: 
 *      vtr_flow/benchmarks/hdl_include/ch_intrinsic_modified.v
*/
`define MEMORY_CONTROLLER_ADDR_SIZE 32
`define MEMORY_CONTROLLER_DATA_SIZE 32