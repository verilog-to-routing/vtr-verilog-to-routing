module simple_op(in,out);
    input  in;
    output out;

    assign out = in;
endmodule