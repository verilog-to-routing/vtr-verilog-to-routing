`define UNARY_OP(out,a) buf(out, a);
`include "wire_test.v"