/*
 * Wide range test
*/

`define WIDTH 3
`define operator nor
`include "../.generic/range_any_width_binary_test.v"