`define BINARY_OP(out,a,b) and(out, a, b);
`include "wire_test.v"