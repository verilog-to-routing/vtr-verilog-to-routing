/*
 * Wide range test
*/

`define WIDTH 3
`define operator notif0
`include "../.generic/replicate_any_width_binary_test.v"