module simple_op(a,b);
input signed [3:0] a;
output unsigned [5:0] b;

assign b = a;

endmodule