`define BINARY_OP(out,a,b) notif0(out, a, b);
`include "../.generic/wire_test.v"