/*
 * Integer range test
*/

`define WIDTH 32
`define operator buf
`include "../.generic/replicate_any_width_unary_test.v"