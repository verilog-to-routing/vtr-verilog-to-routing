
 module ex4LS16_fir(clk, In_X, Out_Y); 

 input clk;
 input [11:0] In_X; 
 output [28 :0] Out_Y; 

 reg [11:0] x0 ;

 wire [14:0] x1 ;
 wire [17:0] x6 ;
 wire [24:0] x59 ;
 wire [24:0] x117 ;
 wire [24:0] y96 ;
 wire [24:0] y153 ;
 wire [22:0] x74 ;
 wire [22:0] x113 ;
 wire [22:0] y86 ;
 wire [22:0] y163 ;
 wire [25:0] x76 ;
 wire [25:0] x76_0_1 ;
 wire [26:0] y122 ;
 wire [25:0] x76_1_1 ;
 wire [26:0] y127 ;
 wire [17:0] x102 ;
 wire [17:0] x102_0_1 ;
 wire [20:0] y41 ;
 wire [17:0] x102_1_1 ;
 wire [18:0] y52 ;
 wire [17:0] x102_2_1 ;
 wire [18:0] y197 ;
 wire [17:0] x102_3_1 ;
 wire [20:0] y208 ;
 wire [17:0] x6_4_1 ;
 wire [17:0] x6_4_2 ;
 wire [17:0] y3 ;
 wire [17:0] x6_5_1 ;
 wire [17:0] x6_5_2 ;
 wire [17:0] y246 ;
 wire [19:0] x10 ;
 wire [21:0] x45 ;
 wire [21:0] x45_0_1 ;
 wire [22:0] y115 ;
 wire [21:0] x45_1_1 ;
 wire [22:0] y134 ;
 wire [19:0] x105 ;
 wire [19:0] x105_0_1 ;
 wire [19:0] y56 ;
 wire [19:0] x105_1_1 ;
 wire [19:0] y193 ;
 wire [19:0] x10_2_1 ;
 wire [19:0] x10_2_2 ;
 wire [19:0] y27 ;
 wire [19:0] x10_3_1 ;
 wire [19:0] x10_3_2 ;
 wire [19:0] y222 ;
 wire [19:0] x11 ;
 wire [24:0] x70 ;
 wire [24:0] x70_0_1 ;
 wire [24:0] y100 ;
 wire [24:0] x70_1_1 ;
 wire [24:0] y149 ;
 wire [19:0] x111 ;
 wire [19:0] x111_0_1 ;
 wire [21:0] y81 ;
 wire [19:0] x111_1_1 ;
 wire [21:0] y168 ;
 wire [19:0] x11_2_1 ;
 wire [19:0] x11_2_2 ;
 wire [21:0] y71 ;
 wire [19:0] x11_3_1 ;
 wire [19:0] x11_3_2 ;
 wire [21:0] y178 ;
 wire [20:0] x12 ;
 wire [20:0] x12_0_1 ;
 wire [20:0] x12_0_2 ;
 wire [20:0] y64 ;
 wire [20:0] x12_1_1 ;
 wire [20:0] x12_1_2 ;
 wire [21:0] y69 ;
 wire [20:0] x12_2_1 ;
 wire [20:0] x12_2_2 ;
 wire [24:0] y112 ;
 wire [20:0] x12_3_1 ;
 wire [20:0] x12_3_2 ;
 wire [24:0] y137 ;
 wire [20:0] x12_4_1 ;
 wire [20:0] x12_4_2 ;
 wire [21:0] y180 ;
 wire [20:0] x12_5_1 ;
 wire [20:0] x12_5_2 ;
 wire [20:0] y185 ;
 wire [18:0] x14 ;
 wire [22:0] x64 ;
 wire [22:0] x64_0_1 ;
 wire [24:0] y110 ;
 wire [22:0] x64_1_1 ;
 wire [24:0] y139 ;
 wire [18:0] x96 ;
 wire [18:0] x96_0_1 ;
 wire [18:0] y17 ;
 wire [18:0] x96_1_1 ;
 wire [18:0] y232 ;
 wire [16:0] x15 ;
 wire [16:0] x15_0_1 ;
 wire [16:0] x15_0_2 ;
 wire [16:0] y26 ;
 wire [16:0] x15_1_1 ;
 wire [16:0] x15_1_2 ;
 wire [16:0] y34 ;
 wire [16:0] x15_2_1 ;
 wire [16:0] x15_2_2 ;
 wire [16:0] y215 ;
 wire [16:0] x15_3_1 ;
 wire [16:0] x15_3_2 ;
 wire [16:0] y223 ;
 wire [21:0] x16 ;
 wire [21:0] x118 ;
 wire [21:0] x118_0_1 ;
 wire [21:0] y105 ;
 wire [21:0] x118_1_1 ;
 wire [21:0] y144 ;
 wire [21:0] x16_1_1 ;
 wire [21:0] x16_1_2 ;
 wire [21:0] y65 ;
 wire [21:0] x16_2_1 ;
 wire [21:0] x16_2_2 ;
 wire [21:0] y184 ;
 wire [20:0] x20 ;
 wire [20:0] x20_0_1 ;
 wire [20:0] x20_0_2 ;
 wire [21:0] y63 ;
 wire [20:0] x20_1_1 ;
 wire [20:0] x20_1_2 ;
 wire [20:0] y95 ;
 wire [20:0] x20_2_1 ;
 wire [20:0] x20_2_2 ;
 wire [20:0] y154 ;
 wire [20:0] x20_3_1 ;
 wire [20:0] x20_3_2 ;
 wire [21:0] y186 ;
 wire [20:0] x21 ;
 wire [20:0] x120 ;
 wire [20:0] x120_0_1 ;
 wire [22:0] y109 ;
 wire [20:0] x120_1_1 ;
 wire [22:0] y140 ;
 wire [20:0] x21_1_1 ;
 wire [20:0] x21_1_2 ;
 wire [20:0] y45 ;
 wire [20:0] x21_2_1 ;
 wire [20:0] x21_2_2 ;
 wire [20:0] y204 ;
 wire [21:0] x22 ;
 wire [21:0] x112 ;
 wire [21:0] x112_0_1 ;
 wire [22:0] y82 ;
 wire [21:0] x112_1_1 ;
 wire [22:0] y167 ;
 wire [21:0] x22_1_1 ;
 wire [21:0] x22_1_2 ;
 wire [21:0] y61 ;
 wire [21:0] x22_2_1 ;
 wire [21:0] x22_2_2 ;
 wire [21:0] y188 ;
 wire [17:0] x27 ;
 wire [17:0] x27_0_1 ;
 wire [17:0] x27_0_2 ;
 wire [17:0] y21 ;
 wire [17:0] x27_1_1 ;
 wire [17:0] x27_1_2 ;
 wire [17:0] y228 ;
 wire [19:0] x28 ;
 wire [19:0] x100 ;
 wire [19:0] x100_0_1 ;
 wire [19:0] y29 ;
 wire [19:0] x100_1_1 ;
 wire [19:0] y220 ;
 wire [18:0] x29 ;
 wire [18:0] x29_0_1 ;
 wire [18:0] x29_0_2 ;
 wire [18:0] y35 ;
 wire [18:0] x29_1_1 ;
 wire [18:0] x29_1_2 ;
 wire [18:0] y214 ;
 wire [20:0] x30 ;
 wire [20:0] x30_0_1 ;
 wire [20:0] x30_0_2 ;
 wire [20:0] y43 ;
 wire [20:0] x30_1_1 ;
 wire [20:0] x30_1_2 ;
 wire [20:0] y206 ;
 wire [17:0] x31 ;
 wire [17:0] x31_0_1 ;
 wire [17:0] x31_0_2 ;
 wire [18:0] y60 ;
 wire [17:0] x31_1_1 ;
 wire [17:0] x31_1_2 ;
 wire [18:0] y189 ;
 wire [19:0] x32 ;
 wire [19:0] x32_0_1 ;
 wire [19:0] x32_0_2 ;
 wire [20:0] y76 ;
 wire [19:0] x32_1_1 ;
 wire [19:0] x32_1_2 ;
 wire [20:0] y173 ;
 wire [23:0] x33 ;
 wire [24:0] x71 ;
 wire [24:0] x71_0_1 ;
 wire [26:0] y118 ;
 wire [24:0] x71_1_1 ;
 wire [26:0] y131 ;
 wire [20:0] x34 ;
 wire [20:0] x34_0_1 ;
 wire [20:0] x34_0_2 ;
 wire [22:0] y104 ;
 wire [20:0] x34_1_1 ;
 wire [20:0] x34_1_2 ;
 wire [22:0] y145 ;
 wire [19:0] x46 ;
 wire [19:0] x46_0_1 ;
 wire [19:0] x46_0_2 ;
 wire [19:0] y101 ;
 wire [19:0] x46_1_1 ;
 wire [19:0] x46_1_2 ;
 wire [19:0] y148 ;
 wire [21:0] x47 ;
 wire [21:0] x47_0_1 ;
 wire [21:0] x47_0_2 ;
 wire [21:0] y85 ;
 wire [21:0] x47_1_1 ;
 wire [21:0] x47_1_2 ;
 wire [21:0] y164 ;
 wire [25:0] x48 ;
 wire [25:0] x48_0_1 ;
 wire [25:0] x48_0_2 ;
 wire [26:0] y123 ;
 wire [25:0] x48_1_1 ;
 wire [25:0] x48_1_2 ;
 wire [26:0] y126 ;
 wire [20:0] x49 ;
 wire [20:0] x49_0_1 ;
 wire [20:0] x49_0_2 ;
 wire [20:0] y62 ;
 wire [20:0] x49_1_1 ;
 wire [20:0] x49_1_2 ;
 wire [20:0] y187 ;
 wire [21:0] x50 ;
 wire [21:0] x50_0_1 ;
 wire [21:0] x50_0_2 ;
 wire [21:0] y67 ;
 wire [21:0] x50_1_1 ;
 wire [21:0] x50_1_2 ;
 wire [21:0] y182 ;
 wire [22:0] x51 ;
 wire [22:0] x51_0_1 ;
 wire [22:0] x51_0_2 ;
 wire [22:0] y84 ;
 wire [22:0] x51_1_1 ;
 wire [22:0] x51_1_2 ;
 wire [22:0] y165 ;
 wire [23:0] x52 ;
 wire [23:0] x52_0_1 ;
 wire [23:0] x52_0_2 ;
 wire [23:0] y98 ;
 wire [23:0] x52_1_1 ;
 wire [23:0] x52_1_2 ;
 wire [23:0] y151 ;
 wire [23:0] x53 ;
 wire [23:0] x119 ;
 wire [23:0] x119_0_1 ;
 wire [23:0] y106 ;
 wire [23:0] x119_1_1 ;
 wire [23:0] y143 ;
 wire [24:0] x54 ;
 wire [24:0] x54_0_1 ;
 wire [24:0] x54_0_2 ;
 wire [24:0] y116 ;
 wire [24:0] x54_1_1 ;
 wire [24:0] x54_1_2 ;
 wire [24:0] y133 ;
 wire [21:0] x55 ;
 wire [21:0] x109 ;
 wire [21:0] x109_0_1 ;
 wire [21:0] y74 ;
 wire [21:0] x109_1_1 ;
 wire [21:0] y175 ;
 wire [20:0] x56 ;
 wire [20:0] x110 ;
 wire [20:0] x110_0_1 ;
 wire [21:0] y75 ;
 wire [20:0] x110_1_1 ;
 wire [21:0] y174 ;
 wire [21:0] x57 ;
 wire [21:0] x57_0_1 ;
 wire [21:0] x57_0_2 ;
 wire [21:0] y87 ;
 wire [21:0] x57_1_1 ;
 wire [21:0] x57_1_2 ;
 wire [21:0] y162 ;
 wire [21:0] x58 ;
 wire [21:0] x58_0_1 ;
 wire [21:0] x58_0_2 ;
 wire [21:0] y83 ;
 wire [21:0] x58_1_1 ;
 wire [21:0] x58_1_2 ;
 wire [21:0] y166 ;
 wire [23:0] x60 ;
 wire [23:0] x60_0_1 ;
 wire [24:0] y117 ;
 wire [23:0] x60_1_1 ;
 wire [24:0] y132 ;
 wire [22:0] x61 ;
 wire [22:0] x61_0_1 ;
 wire [22:0] x61_0_2 ;
 wire [23:0] y113 ;
 wire [22:0] x61_1_1 ;
 wire [22:0] x61_1_2 ;
 wire [23:0] y136 ;
 wire [20:0] x62 ;
 wire [20:0] x62_0_1 ;
 wire [20:0] x62_0_2 ;
 wire [20:0] y47 ;
 wire [20:0] x62_1_1 ;
 wire [20:0] x62_1_2 ;
 wire [20:0] y202 ;
 wire [20:0] x63 ;
 wire [20:0] x63_0_1 ;
 wire [20:0] x63_0_2 ;
 wire [20:0] y55 ;
 wire [20:0] x63_1_1 ;
 wire [20:0] x63_1_2 ;
 wire [20:0] y194 ;
 wire [20:0] x65 ;
 wire [20:0] x65_0_1 ;
 wire [20:0] x65_0_2 ;
 wire [20:0] y53 ;
 wire [20:0] x65_1_1 ;
 wire [20:0] x65_1_2 ;
 wire [20:0] y196 ;
 wire [24:0] x66 ;
 wire [24:0] x121 ;
 wire [24:0] x121_0_1 ;
 wire [25:0] y121 ;
 wire [24:0] x121_1_1 ;
 wire [25:0] y128 ;
 wire [14:0] x92 ;
 wire [14:0] x92_0_1 ;
 wire [14:0] x92_0_2 ;
 wire [16:0] y5 ;
 wire [14:0] x92_1_1 ;
 wire [14:0] x92_1_2 ;
 wire [16:0] y14 ;
 wire [14:0] x92_2_1 ;
 wire [14:0] x92_2_2 ;
 wire [15:0] y48 ;
 wire [14:0] x92_3_1 ;
 wire [14:0] x92_3_2 ;
 wire [20:0] y72 ;
 wire [14:0] x92_4_1 ;
 wire [14:0] x92_4_2 ;
 wire [20:0] y177 ;
 wire [14:0] x92_5_1 ;
 wire [14:0] x92_5_2 ;
 wire [15:0] y201 ;
 wire [14:0] x92_6_1 ;
 wire [14:0] x92_6_2 ;
 wire [16:0] y235 ;
 wire [14:0] x92_7_1 ;
 wire [14:0] x92_7_2 ;
 wire [16:0] y244 ;
 wire [14:0] x1_42_1 ;
 wire [14:0] x1_42_2 ;
 wire [14:0] x1_42_3 ;
 wire [14:0] y4 ;
 wire [14:0] x1_43_1 ;
 wire [14:0] x1_43_2 ;
 wire [14:0] x1_43_3 ;
 wire [16:0] y12 ;
 wire [14:0] x1_44_1 ;
 wire [14:0] x1_44_2 ;
 wire [14:0] x1_44_3 ;
 wire [15:0] y44 ;
 wire [14:0] x1_45_1 ;
 wire [14:0] x1_45_2 ;
 wire [14:0] x1_45_3 ;
 wire [15:0] y205 ;
 wire [14:0] x1_46_1 ;
 wire [14:0] x1_46_2 ;
 wire [14:0] x1_46_3 ;
 wire [16:0] y237 ;
 wire [14:0] x1_47_1 ;
 wire [14:0] x1_47_2 ;
 wire [14:0] x1_47_3 ;
 wire [14:0] y245 ;
 wire [14:0] x2 ;
 wire [17:0] x7 ;
 wire [19:0] x77 ;
 wire [19:0] x77_0_1 ;
 wire [20:0] y73 ;
 wire [21:0] x80 ;
 wire [21:0] x114 ;
 wire [21:0] y90 ;
 wire [19:0] x81 ;
 wire [19:0] x115 ;
 wire [19:0] y91 ;
 wire [20:0] x82 ;
 wire [20:0] x82_0_1 ;
 wire [22:0] y102 ;
 wire [20:0] x85 ;
 wire [20:0] x85_0_1 ;
 wire [22:0] y147 ;
 wire [19:0] x86 ;
 wire [19:0] x122 ;
 wire [19:0] y158 ;
 wire [21:0] x87 ;
 wire [21:0] x123 ;
 wire [21:0] y159 ;
 wire [19:0] x90 ;
 wire [19:0] x90_0_1 ;
 wire [20:0] y176 ;
 wire [17:0] x95 ;
 wire [17:0] x95_0_1 ;
 wire [17:0] y15 ;
 wire [17:0] x95_1_1 ;
 wire [17:0] y28 ;
 wire [17:0] x95_2_1 ;
 wire [20:0] y70 ;
 wire [17:0] x95_3_1 ;
 wire [20:0] y179 ;
 wire [17:0] x95_4_1 ;
 wire [17:0] y221 ;
 wire [17:0] x95_5_1 ;
 wire [17:0] y234 ;
 wire [17:0] x7_10_1 ;
 wire [17:0] x7_10_2 ;
 wire [20:0] y89 ;
 wire [17:0] x7_11_1 ;
 wire [17:0] x7_11_2 ;
 wire [20:0] y160 ;
 wire [17:0] x9 ;
 wire [21:0] x78 ;
 wire [21:0] x78_0_1 ;
 wire [21:0] y77 ;
 wire [21:0] x79 ;
 wire [21:0] x79_0_1 ;
 wire [21:0] y79 ;
 wire [23:0] x83 ;
 wire [23:0] x83_0_1 ;
 wire [24:0] y120 ;
 wire [23:0] x84 ;
 wire [23:0] x84_0_1 ;
 wire [24:0] y129 ;
 wire [21:0] x88 ;
 wire [21:0] x88_0_1 ;
 wire [21:0] y170 ;
 wire [21:0] x89 ;
 wire [21:0] x89_0_1 ;
 wire [21:0] y172 ;
 wire [17:0] x9_7_1 ;
 wire [17:0] x9_7_2 ;
 wire [17:0] y19 ;
 wire [17:0] x9_8_1 ;
 wire [17:0] x9_8_2 ;
 wire [18:0] y31 ;
 wire [17:0] x9_9_1 ;
 wire [17:0] x9_9_2 ;
 wire [18:0] y218 ;
 wire [17:0] x9_10_1 ;
 wire [17:0] x9_10_2 ;
 wire [17:0] y230 ;
 wire [17:0] x17 ;
 wire [24:0] x75 ;
 wire [24:0] x75_0_1 ;
 wire [24:0] y119 ;
 wire [24:0] x75_1_1 ;
 wire [24:0] y130 ;
 wire [17:0] x17_1_1 ;
 wire [17:0] x17_1_2 ;
 wire [17:0] y25 ;
 wire [17:0] x17_2_1 ;
 wire [17:0] x17_2_2 ;
 wire [17:0] y224 ;
 wire [19:0] x18 ;
 wire [19:0] x18_0_1 ;
 wire [19:0] x18_0_2 ;
 wire [19:0] y49 ;
 wire [19:0] x18_1_1 ;
 wire [19:0] x18_1_2 ;
 wire [19:0] y93 ;
 wire [19:0] x18_2_1 ;
 wire [19:0] x18_2_2 ;
 wire [19:0] y156 ;
 wire [19:0] x18_3_1 ;
 wire [19:0] x18_3_2 ;
 wire [19:0] y200 ;
 wire [18:0] x35 ;
 wire [18:0] x35_0_1 ;
 wire [18:0] x35_0_2 ;
 wire [18:0] y33 ;
 wire [18:0] x35_1_1 ;
 wire [18:0] x35_1_2 ;
 wire [18:0] y216 ;
 wire [19:0] x36 ;
 wire [19:0] x101 ;
 wire [19:0] x101_0_1 ;
 wire [19:0] y39 ;
 wire [19:0] x101_1_1 ;
 wire [19:0] y210 ;
 wire [19:0] x37 ;
 wire [19:0] x103 ;
 wire [19:0] x103_0_1 ;
 wire [19:0] y51 ;
 wire [19:0] x103_1_1 ;
 wire [19:0] y198 ;
 wire [19:0] x38 ;
 wire [19:0] x38_0_1 ;
 wire [19:0] x38_0_2 ;
 wire [21:0] y80 ;
 wire [19:0] x38_1_1 ;
 wire [19:0] x38_1_2 ;
 wire [21:0] y169 ;
 wire [23:0] x39 ;
 wire [23:0] x39_0_1 ;
 wire [23:0] x39_0_2 ;
 wire [23:0] y108 ;
 wire [23:0] x39_1_1 ;
 wire [23:0] x39_1_2 ;
 wire [23:0] y141 ;
 wire [19:0] x67 ;
 wire [19:0] x107 ;
 wire [19:0] x107_0_1 ;
 wire [20:0] y59 ;
 wire [19:0] x107_1_1 ;
 wire [20:0] y190 ;
 wire [22:0] x68 ;
 wire [22:0] x116 ;
 wire [22:0] x116_0_1 ;
 wire [22:0] y94 ;
 wire [22:0] x116_1_1 ;
 wire [22:0] y155 ;
 wire [21:0] x69 ;
 wire [21:0] x69_0_1 ;
 wire [21:0] x69_0_2 ;
 wire [21:0] y78 ;
 wire [21:0] x69_1_1 ;
 wire [21:0] x69_1_2 ;
 wire [21:0] y171 ;
 wire [14:0] x99 ;
 wire [14:0] x99_0_1 ;
 wire [14:0] x99_0_2 ;
 wire [16:0] y24 ;
 wire [14:0] x99_1_1 ;
 wire [14:0] x99_1_2 ;
 wire [16:0] y32 ;
 wire [14:0] x99_2_1 ;
 wire [14:0] x99_2_2 ;
 wire [15:0] y99 ;
 wire [14:0] x99_3_1 ;
 wire [14:0] x99_3_2 ;
 wire [15:0] y150 ;
 wire [14:0] x99_4_1 ;
 wire [14:0] x99_4_2 ;
 wire [16:0] y217 ;
 wire [14:0] x99_5_1 ;
 wire [14:0] x99_5_2 ;
 wire [16:0] y225 ;
 wire [14:0] x2_21_1 ;
 wire [14:0] x2_21_2 ;
 wire [14:0] x2_21_3 ;
 wire [14:0] y0 ;
 wire [14:0] x2_22_1 ;
 wire [14:0] x2_22_2 ;
 wire [14:0] x2_22_3 ;
 wire [14:0] y6 ;
 wire [14:0] x2_23_1 ;
 wire [14:0] x2_23_2 ;
 wire [14:0] x2_23_3 ;
 wire [16:0] y30 ;
 wire [14:0] x2_24_1 ;
 wire [14:0] x2_24_2 ;
 wire [14:0] x2_24_3 ;
 wire [19:0] y57 ;
 wire [14:0] x2_25_1 ;
 wire [14:0] x2_25_2 ;
 wire [14:0] x2_25_3 ;
 wire [19:0] y192 ;
 wire [14:0] x2_26_1 ;
 wire [14:0] x2_26_2 ;
 wire [14:0] x2_26_3 ;
 wire [16:0] y219 ;
 wire [14:0] x2_27_1 ;
 wire [14:0] x2_27_2 ;
 wire [14:0] x2_27_3 ;
 wire [14:0] y243 ;
 wire [14:0] x2_28_1 ;
 wire [14:0] x2_28_2 ;
 wire [14:0] x2_28_3 ;
 wire [14:0] y249 ;
 wire [15:0] x3 ;
 wire [19:0] x19 ;
 wire [19:0] x19_0_1 ;
 wire [19:0] x19_0_2 ;
 wire [19:0] y37 ;
 wire [19:0] x19_1_1 ;
 wire [19:0] x19_1_2 ;
 wire [21:0] y107 ;
 wire [19:0] x19_2_1 ;
 wire [19:0] x19_2_2 ;
 wire [21:0] y142 ;
 wire [19:0] x19_3_1 ;
 wire [19:0] x19_3_2 ;
 wire [19:0] y212 ;
 wire [18:0] x40 ;
 wire [18:0] x40_0_1 ;
 wire [18:0] x40_0_2 ;
 wire [18:0] y97 ;
 wire [18:0] x40_1_1 ;
 wire [18:0] x40_1_2 ;
 wire [18:0] y152 ;
 wire [22:0] x72 ;
 wire [22:0] x72_0_1 ;
 wire [22:0] x72_0_2 ;
 wire [22:0] y92 ;
 wire [22:0] x72_1_1 ;
 wire [22:0] x72_1_2 ;
 wire [22:0] y157 ;
 wire [22:0] x73 ;
 wire [22:0] x73_0_1 ;
 wire [22:0] x73_0_2 ;
 wire [22:0] y111 ;
 wire [22:0] x73_1_1 ;
 wire [22:0] x73_1_2 ;
 wire [22:0] y138 ;
 wire [15:0] x98 ;
 wire [15:0] x98_0_1 ;
 wire [15:0] x98_0_2 ;
 wire [16:0] y20 ;
 wire [15:0] x98_1_1 ;
 wire [15:0] x98_1_2 ;
 wire [16:0] y36 ;
 wire [15:0] x98_2_1 ;
 wire [15:0] x98_2_2 ;
 wire [16:0] y213 ;
 wire [15:0] x98_3_1 ;
 wire [15:0] x98_3_2 ;
 wire [16:0] y229 ;
 wire [15:0] x3_14_1 ;
 wire [15:0] x3_14_2 ;
 wire [15:0] x3_14_3 ;
 wire [15:0] y10 ;
 wire [15:0] x3_15_1 ;
 wire [15:0] x3_15_2 ;
 wire [15:0] x3_15_3 ;
 wire [16:0] y13 ;
 wire [15:0] x3_16_1 ;
 wire [15:0] x3_16_2 ;
 wire [15:0] x3_16_3 ;
 wire [16:0] y22 ;
 wire [15:0] x3_17_1 ;
 wire [15:0] x3_17_2 ;
 wire [15:0] x3_17_3 ;
 wire [15:0] y42 ;
 wire [15:0] x3_18_1 ;
 wire [15:0] x3_18_2 ;
 wire [15:0] x3_18_3 ;
 wire [19:0] y68 ;
 wire [15:0] x3_19_1 ;
 wire [15:0] x3_19_2 ;
 wire [15:0] x3_19_3 ;
 wire [19:0] y181 ;
 wire [15:0] x3_20_1 ;
 wire [15:0] x3_20_2 ;
 wire [15:0] x3_20_3 ;
 wire [15:0] y207 ;
 wire [15:0] x3_21_1 ;
 wire [15:0] x3_21_2 ;
 wire [15:0] x3_21_3 ;
 wire [16:0] y227 ;
 wire [15:0] x3_22_1 ;
 wire [15:0] x3_22_2 ;
 wire [15:0] x3_22_3 ;
 wire [16:0] y236 ;
 wire [15:0] x3_23_1 ;
 wire [15:0] x3_23_2 ;
 wire [15:0] x3_23_3 ;
 wire [15:0] y239 ;
 wire [15:0] x4 ;
 wire [19:0] x41 ;
 wire [19:0] x106 ;
 wire [19:0] x106_0_1 ;
 wire [19:0] y58 ;
 wire [19:0] x106_1_1 ;
 wire [19:0] y191 ;
 wire [20:0] x42 ;
 wire [20:0] x42_0_1 ;
 wire [20:0] x42_0_2 ;
 wire [20:0] y103 ;
 wire [20:0] x42_1_1 ;
 wire [20:0] x42_1_2 ;
 wire [20:0] y146 ;
 wire [15:0] x93 ;
 wire [15:0] x93_0_1 ;
 wire [15:0] x93_0_2 ;
 wire [16:0] y7 ;
 wire [15:0] x93_1_1 ;
 wire [15:0] x93_1_2 ;
 wire [16:0] y40 ;
 wire [15:0] x93_2_1 ;
 wire [15:0] x93_2_2 ;
 wire [16:0] y50 ;
 wire [15:0] x93_3_1 ;
 wire [15:0] x93_3_2 ;
 wire [16:0] y199 ;
 wire [15:0] x93_4_1 ;
 wire [15:0] x93_4_2 ;
 wire [16:0] y209 ;
 wire [15:0] x93_5_1 ;
 wire [15:0] x93_5_2 ;
 wire [16:0] y242 ;
 wire [15:0] x4_10_1 ;
 wire [15:0] x4_10_2 ;
 wire [15:0] x4_10_3 ;
 wire [15:0] y1 ;
 wire [15:0] x4_11_1 ;
 wire [15:0] x4_11_2 ;
 wire [15:0] x4_11_3 ;
 wire [16:0] y9 ;
 wire [15:0] x4_12_1 ;
 wire [15:0] x4_12_2 ;
 wire [15:0] x4_12_3 ;
 wire [16:0] y240 ;
 wire [15:0] x4_13_1 ;
 wire [15:0] x4_13_2 ;
 wire [15:0] x4_13_3 ;
 wire [15:0] y248 ;
 wire [16:0] x5 ;
 wire [21:0] x43 ;
 wire [21:0] x43_0_1 ;
 wire [21:0] x43_0_2 ;
 wire [22:0] y88 ;
 wire [21:0] x43_1_1 ;
 wire [21:0] x43_1_2 ;
 wire [22:0] y161 ;
 wire [24:0] x44 ;
 wire [24:0] x44_0_1 ;
 wire [24:0] x44_0_2 ;
 wire [24:0] y114 ;
 wire [24:0] x44_1_1 ;
 wire [24:0] x44_1_2 ;
 wire [24:0] y135 ;
 wire [16:0] x97 ;
 wire [16:0] x97_0_1 ;
 wire [16:0] x97_0_2 ;
 wire [16:0] y18 ;
 wire [16:0] x97_1_1 ;
 wire [16:0] x97_1_2 ;
 wire [16:0] y38 ;
 wire [16:0] x97_2_1 ;
 wire [16:0] x97_2_2 ;
 wire [16:0] y211 ;
 wire [16:0] x97_3_1 ;
 wire [16:0] x97_3_2 ;
 wire [16:0] y231 ;
 wire [16:0] x5_5_1 ;
 wire [16:0] x5_5_2 ;
 wire [16:0] x5_5_3 ;
 wire [16:0] y16 ;
 wire [16:0] x5_6_1 ;
 wire [16:0] x5_6_2 ;
 wire [16:0] x5_6_3 ;
 wire [16:0] y233 ;
 wire [16:0] x8 ;
 wire [16:0] x94 ;
 wire [16:0] x94_0_1 ;
 wire [16:0] x94_0_2 ;
 wire [16:0] y11 ;
 wire [16:0] x94_1_1 ;
 wire [16:0] x94_1_2 ;
 wire [17:0] y23 ;
 wire [16:0] x94_2_1 ;
 wire [16:0] x94_2_2 ;
 wire [17:0] y226 ;
 wire [16:0] x94_3_1 ;
 wire [16:0] x94_3_2 ;
 wire [16:0] y238 ;
 wire [19:0] x13 ;
 wire [17:0] x23 ;
 wire [17:0] x108 ;
 wire [17:0] x108_0_1 ;
 wire [17:0] x108_0_2 ;
 wire [19:0] y66 ;
 wire [17:0] x108_1_1 ;
 wire [17:0] x108_1_2 ;
 wire [19:0] y183 ;
 wire [17:0] x24 ;
 wire [17:0] x104 ;
 wire [17:0] x104_0_1 ;
 wire [17:0] x104_0_2 ;
 wire [17:0] y54 ;
 wire [17:0] x104_1_1 ;
 wire [17:0] x104_1_2 ;
 wire [17:0] y195 ;
 wire [19:0] x25 ;
 wire [23:0] x26 ;
 wire [11:0] x77_50_1 ;
 wire [11:0] x77_50_2 ;
 wire [11:0] x78_51_1 ;
 wire [11:0] x78_51_2 ;
 wire [11:0] x79_52_1 ;
 wire [11:0] x79_52_2 ;
 wire [11:0] x80_53_1 ;
 wire [11:0] x80_53_2 ;
 wire [11:0] x81_54_1 ;
 wire [11:0] x81_54_2 ;
 wire [11:0] x82_55_1 ;
 wire [11:0] x82_55_2 ;
 wire [11:0] x83_56_1 ;
 wire [11:0] x83_56_2 ;
 wire [11:0] x84_57_1 ;
 wire [11:0] x84_57_2 ;
 wire [11:0] x85_58_1 ;
 wire [11:0] x85_58_2 ;
 wire [11:0] x86_59_1 ;
 wire [11:0] x86_59_2 ;
 wire [11:0] x87_60_1 ;
 wire [11:0] x87_60_2 ;
 wire [11:0] x88_61_1 ;
 wire [11:0] x88_61_2 ;
 wire [11:0] x89_62_1 ;
 wire [11:0] x89_62_2 ;
 wire [11:0] x90_63_1 ;
 wire [11:0] x90_63_2 ;
 wire [11:0] x91 ;
 wire [11:0] x91_0_1 ;
 wire [11:0] x91_0_2 ;
 wire [11:0] x91_0_3 ;
 wire [12:0] y2 ;
 wire [11:0] x91_1_1 ;
 wire [11:0] x91_1_2 ;
 wire [11:0] x91_1_3 ;
 wire [14:0] y8 ;
 wire [11:0] x91_2_1 ;
 wire [11:0] x91_2_2 ;
 wire [11:0] x91_2_3 ;
 wire [11:0] y46 ;
 wire [11:0] x91_3_1 ;
 wire [11:0] x91_3_2 ;
 wire [11:0] x91_3_3 ;
 wire [11:0] y203 ;
 wire [11:0] x91_4_1 ;
 wire [11:0] x91_4_2 ;
 wire [11:0] x91_4_3 ;
 wire [14:0] y241 ;
 wire [11:0] x91_5_1 ;
 wire [11:0] x91_5_2 ;
 wire [11:0] x91_5_3 ;
 wire [12:0] y247 ;
 wire [11:0] x0_65_1 ;
 wire [11:0] x0_65_2 ;
 wire [11:0] x0_65_3 ;
 wire [11:0] x0_65_4 ;
 wire [26:0] y124 ;
 wire [11:0] x0_66_1 ;
 wire [11:0] x0_66_2 ;
 wire [11:0] x0_66_3 ;
 wire [11:0] x0_66_4 ;
 wire [26:0] y125 ;
 wire [14:0] x124 ;
 wire [16:0] x125 ;
 wire [16:0] x125_1 ;
 wire [17:0] x126 ;
 wire [17:0] x126_1 ;
 wire [18:0] x127 ;
 wire [18:0] x127_1 ;
 wire [19:0] x128 ;
 wire [19:0] x128_1 ;
 wire [20:0] x129 ;
 wire [20:0] x129_1 ;
 wire [21:0] x130 ;
 wire [21:0] x130_1 ;
 wire [22:0] x131 ;
 wire [22:0] x131_1 ;
 wire [23:0] x132 ;
 wire [23:0] x132_1 ;
 wire [24:0] x133 ;
 wire [24:0] x133_1 ;
 wire [25:0] x134 ;
 wire [25:0] x134_1 ;
 wire [26:0] x135 ;
 wire [26:0] x135_1 ;
 wire [27:0] x136 ;
 wire [27:0] x136_1 ;
 wire [28:0] x137 ;
 wire [28:0] x137_1 ;
 wire [28:0] x138 ;
 wire [28:0] x138_1 ;
 wire [28:0] x139 ;
 wire [28:0] x139_1 ;
 wire [28:0] x140 ;
 wire [28:0] x140_1 ;
 wire [28:0] x141 ;
 wire [28:0] x141_1 ;
 wire [28:0] x142 ;
 wire [28:0] x142_1 ;
 wire [28:0] x143 ;
 wire [28:0] x143_1 ;
 wire [28:0] x144 ;
 wire [28:0] x144_1 ;
 wire [28:0] x145 ;
 wire [28:0] x145_1 ;
 wire [28:0] x146 ;
 wire [28:0] x146_1 ;
 wire [28:0] x147 ;
 wire [28:0] x147_1 ;
 wire [28:0] x148 ;
 wire [28:0] x148_1 ;
 wire [28:0] x149 ;
 wire [28:0] x149_1 ;
 wire [28:0] x150 ;
 wire [28:0] x150_1 ;
 wire [28:0] x151 ;
 wire [28:0] x151_1 ;
 wire [28:0] x152 ;
 wire [28:0] x152_1 ;
 wire [28:0] x153 ;
 wire [28:0] x153_1 ;
 wire [28:0] x154 ;
 wire [28:0] x154_1 ;
 wire [28:0] x155 ;
 wire [28:0] x155_1 ;
 wire [28:0] x156 ;
 wire [28:0] x156_1 ;
 wire [28:0] x157 ;
 wire [28:0] x157_1 ;
 wire [28:0] x158 ;
 wire [28:0] x158_1 ;
 wire [28:0] x159 ;
 wire [28:0] x159_1 ;
 wire [28:0] x160 ;
 wire [28:0] x160_1 ;
 wire [28:0] x161 ;
 wire [28:0] x161_1 ;
 wire [28:0] x162 ;
 wire [28:0] x162_1 ;
 wire [28:0] x163 ;
 wire [28:0] x163_1 ;
 wire [28:0] x164 ;
 wire [28:0] x164_1 ;
 wire [28:0] x165 ;
 wire [28:0] x165_1 ;
 wire [28:0] x166 ;
 wire [28:0] x166_1 ;
 wire [28:0] x167 ;
 wire [28:0] x167_1 ;
 wire [28:0] x168 ;
 wire [28:0] x168_1 ;
 wire [28:0] x169 ;
 wire [28:0] x169_1 ;
 wire [28:0] x170 ;
 wire [28:0] x170_1 ;
 wire [28:0] x171 ;
 wire [28:0] x171_1 ;
 wire [28:0] x172 ;
 wire [28:0] x172_1 ;
 wire [28:0] x173 ;
 wire [28:0] x173_1 ;
 wire [28:0] x174 ;
 wire [28:0] x174_1 ;
 wire [28:0] x175 ;
 wire [28:0] x175_1 ;
 wire [28:0] x176 ;
 wire [28:0] x176_1 ;
 wire [28:0] x177 ;
 wire [28:0] x177_1 ;
 wire [28:0] x178 ;
 wire [28:0] x178_1 ;
 wire [28:0] x179 ;
 wire [28:0] x179_1 ;
 wire [28:0] x180 ;
 wire [28:0] x180_1 ;
 wire [28:0] x181 ;
 wire [28:0] x181_1 ;
 wire [28:0] x182 ;
 wire [28:0] x182_1 ;
 wire [28:0] x183 ;
 wire [28:0] x183_1 ;
 wire [28:0] x184 ;
 wire [28:0] x184_1 ;
 wire [28:0] x185 ;
 wire [28:0] x185_1 ;
 wire [28:0] x186 ;
 wire [28:0] x186_1 ;
 wire [28:0] x187 ;
 wire [28:0] x187_1 ;
 wire [28:0] x188 ;
 wire [28:0] x188_1 ;
 wire [28:0] x189 ;
 wire [28:0] x189_1 ;
 wire [28:0] x190 ;
 wire [28:0] x190_1 ;
 wire [28:0] x191 ;
 wire [28:0] x191_1 ;
 wire [28:0] x192 ;
 wire [28:0] x192_1 ;
 wire [28:0] x193 ;
 wire [28:0] x193_1 ;
 wire [28:0] x194 ;
 wire [28:0] x194_1 ;
 wire [28:0] x195 ;
 wire [28:0] x195_1 ;
 wire [28:0] x196 ;
 wire [28:0] x196_1 ;
 wire [28:0] x197 ;
 wire [28:0] x197_1 ;
 wire [28:0] x198 ;
 wire [28:0] x198_1 ;
 wire [28:0] x199 ;
 wire [28:0] x199_1 ;
 wire [28:0] x200 ;
 wire [28:0] x200_1 ;
 wire [28:0] x201 ;
 wire [28:0] x201_1 ;
 wire [28:0] x202 ;
 wire [28:0] x202_1 ;
 wire [28:0] x203 ;
 wire [28:0] x203_1 ;
 wire [28:0] x204 ;
 wire [28:0] x204_1 ;
 wire [28:0] x205 ;
 wire [28:0] x205_1 ;
 wire [28:0] x206 ;
 wire [28:0] x206_1 ;
 wire [28:0] x207 ;
 wire [28:0] x207_1 ;
 wire [28:0] x208 ;
 wire [28:0] x208_1 ;
 wire [28:0] x209 ;
 wire [28:0] x209_1 ;
 wire [28:0] x210 ;
 wire [28:0] x210_1 ;
 wire [28:0] x211 ;
 wire [28:0] x211_1 ;
 wire [28:0] x212 ;
 wire [28:0] x212_1 ;
 wire [28:0] x213 ;
 wire [28:0] x213_1 ;
 wire [28:0] x214 ;
 wire [28:0] x214_1 ;
 wire [28:0] x215 ;
 wire [28:0] x215_1 ;
 wire [28:0] x216 ;
 wire [28:0] x216_1 ;
 wire [28:0] x217 ;
 wire [28:0] x217_1 ;
 wire [28:0] x218 ;
 wire [28:0] x218_1 ;
 wire [28:0] x219 ;
 wire [28:0] x219_1 ;
 wire [28:0] x220 ;
 wire [28:0] x220_1 ;
 wire [28:0] x221 ;
 wire [28:0] x221_1 ;
 wire [28:0] x222 ;
 wire [28:0] x222_1 ;
 wire [28:0] x223 ;
 wire [28:0] x223_1 ;
 wire [28:0] x224 ;
 wire [28:0] x224_1 ;
 wire [28:0] x225 ;
 wire [28:0] x225_1 ;
 wire [28:0] x226 ;
 wire [28:0] x226_1 ;
 wire [28:0] x227 ;
 wire [28:0] x227_1 ;
 wire [28:0] x228 ;
 wire [28:0] x228_1 ;
 wire [28:0] x229 ;
 wire [28:0] x229_1 ;
 wire [28:0] x230 ;
 wire [28:0] x230_1 ;
 wire [28:0] x231 ;
 wire [28:0] x231_1 ;
 wire [28:0] x232 ;
 wire [28:0] x232_1 ;
 wire [28:0] x233 ;
 wire [28:0] x233_1 ;
 wire [28:0] x234 ;
 wire [28:0] x234_1 ;
 wire [28:0] x235 ;
 wire [28:0] x235_1 ;
 wire [28:0] x236 ;
 wire [28:0] x236_1 ;
 wire [28:0] x237 ;
 wire [28:0] x237_1 ;
 wire [28:0] x238 ;
 wire [28:0] x238_1 ;
 wire [28:0] x239 ;
 wire [28:0] x239_1 ;
 wire [28:0] x240 ;
 wire [28:0] x240_1 ;
 wire [28:0] x241 ;
 wire [28:0] x241_1 ;
 wire [28:0] x242 ;
 wire [28:0] x242_1 ;
 wire [28:0] x243 ;
 wire [28:0] x243_1 ;
 wire [28:0] x244 ;
 wire [28:0] x244_1 ;
 wire [28:0] x245 ;
 wire [28:0] x245_1 ;
 wire [28:0] x246 ;
 wire [28:0] x246_1 ;
 wire [28:0] x247 ;
 wire [28:0] x247_1 ;
 wire [28:0] x248 ;
 wire [28:0] x248_1 ;
 wire [28:0] x249 ;
 wire [28:0] x249_1 ;
 wire [28:0] x250 ;
 wire [28:0] x250_1 ;
 wire [28:0] x251 ;
 wire [28:0] x251_1 ;
 wire [28:0] x252 ;
 wire [28:0] x252_1 ;
 wire [28:0] x253 ;
 wire [28:0] x253_1 ;
 wire [28:0] x254 ;
 wire [28:0] x254_1 ;
 wire [28:0] x255 ;
 wire [28:0] x255_1 ;
 wire [28:0] x256 ;
 wire [28:0] x256_1 ;
 wire [28:0] x257 ;
 wire [28:0] x257_1 ;
 wire [28:0] x258 ;
 wire [28:0] x258_1 ;
 wire [28:0] x259 ;
 wire [28:0] x259_1 ;
 wire [28:0] x260 ;
 wire [28:0] x260_1 ;
 wire [28:0] x261 ;
 wire [28:0] x261_1 ;
 wire [28:0] x262 ;
 wire [28:0] x262_1 ;
 wire [28:0] x263 ;
 wire [28:0] x263_1 ;
 wire [28:0] x264 ;
 wire [28:0] x264_1 ;
 wire [28:0] x265 ;
 wire [28:0] x265_1 ;
 wire [28:0] x266 ;
 wire [28:0] x266_1 ;
 wire [28:0] x267 ;
 wire [28:0] x267_1 ;
 wire [28:0] x268 ;
 wire [28:0] x268_1 ;
 wire [28:0] x269 ;
 wire [28:0] x269_1 ;
 wire [28:0] x270 ;
 wire [28:0] x270_1 ;
 wire [28:0] x271 ;
 wire [28:0] x271_1 ;
 wire [28:0] x272 ;
 wire [28:0] x272_1 ;
 wire [28:0] x273 ;
 wire [28:0] x273_1 ;
 wire [28:0] x274 ;
 wire [28:0] x274_1 ;
 wire [28:0] x275 ;
 wire [28:0] x275_1 ;
 wire [28:0] x276 ;
 wire [28:0] x276_1 ;
 wire [28:0] x277 ;
 wire [28:0] x277_1 ;
 wire [28:0] x278 ;
 wire [28:0] x278_1 ;
 wire [28:0] x279 ;
 wire [28:0] x279_1 ;
 wire [28:0] x280 ;
 wire [28:0] x280_1 ;
 wire [28:0] x281 ;
 wire [28:0] x281_1 ;
 wire [28:0] x282 ;
 wire [28:0] x282_1 ;
 wire [28:0] x283 ;
 wire [28:0] x283_1 ;
 wire [28:0] x284 ;
 wire [28:0] x284_1 ;
 wire [28:0] x285 ;
 wire [28:0] x285_1 ;
 wire [28:0] x286 ;
 wire [28:0] x286_1 ;
 wire [28:0] x287 ;
 wire [28:0] x287_1 ;
 wire [28:0] x288 ;
 wire [28:0] x288_1 ;
 wire [28:0] x289 ;
 wire [28:0] x289_1 ;
 wire [28:0] x290 ;
 wire [28:0] x290_1 ;
 wire [28:0] x291 ;
 wire [28:0] x291_1 ;
 wire [28:0] x292 ;
 wire [28:0] x292_1 ;
 wire [28:0] x293 ;
 wire [28:0] x293_1 ;
 wire [28:0] x294 ;
 wire [28:0] x294_1 ;
 wire [28:0] x295 ;
 wire [28:0] x295_1 ;
 wire [28:0] x296 ;
 wire [28:0] x296_1 ;
 wire [28:0] x297 ;
 wire [28:0] x297_1 ;
 wire [28:0] x298 ;
 wire [28:0] x298_1 ;
 wire [28:0] x299 ;
 wire [28:0] x299_1 ;
 wire [28:0] x300 ;
 wire [28:0] x300_1 ;
 wire [28:0] x301 ;
 wire [28:0] x301_1 ;
 wire [28:0] x302 ;
 wire [28:0] x302_1 ;
 wire [28:0] x303 ;
 wire [28:0] x303_1 ;
 wire [28:0] x304 ;
 wire [28:0] x304_1 ;
 wire [28:0] x305 ;
 wire [28:0] x305_1 ;
 wire [28:0] x306 ;
 wire [28:0] x306_1 ;
 wire [28:0] x307 ;
 wire [28:0] x307_1 ;
 wire [28:0] x308 ;
 wire [28:0] x308_1 ;
 wire [28:0] x309 ;
 wire [28:0] x309_1 ;
 wire [28:0] x310 ;
 wire [28:0] x310_1 ;
 wire [28:0] x311 ;
 wire [28:0] x311_1 ;
 wire [28:0] x312 ;
 wire [28:0] x312_1 ;
 wire [28:0] x313 ;
 wire [28:0] x313_1 ;
 wire [28:0] x314 ;
 wire [28:0] x314_1 ;
 wire [28:0] x315 ;
 wire [28:0] x315_1 ;
 wire [28:0] x316 ;
 wire [28:0] x316_1 ;
 wire [28:0] x317 ;
 wire [28:0] x317_1 ;
 wire [28:0] x318 ;
 wire [28:0] x318_1 ;
 wire [28:0] x319 ;
 wire [28:0] x319_1 ;
 wire [28:0] x320 ;
 wire [28:0] x320_1 ;
 wire [28:0] x321 ;
 wire [28:0] x321_1 ;
 wire [28:0] x322 ;
 wire [28:0] x322_1 ;
 wire [28:0] x323 ;
 wire [28:0] x323_1 ;
 wire [28:0] x324 ;
 wire [28:0] x324_1 ;
 wire [28:0] x325 ;
 wire [28:0] x325_1 ;
 wire [28:0] x326 ;
 wire [28:0] x326_1 ;
 wire [28:0] x327 ;
 wire [28:0] x327_1 ;
 wire [28:0] x328 ;
 wire [28:0] x328_1 ;
 wire [28:0] x329 ;
 wire [28:0] x329_1 ;
 wire [28:0] x330 ;
 wire [28:0] x330_1 ;
 wire [28:0] x331 ;
 wire [28:0] x331_1 ;
 wire [28:0] x332 ;
 wire [28:0] x332_1 ;
 wire [28:0] x333 ;
 wire [28:0] x333_1 ;
 wire [28:0] x334 ;
 wire [28:0] x334_1 ;
 wire [28:0] x335 ;
 wire [28:0] x335_1 ;
 wire [28:0] x336 ;
 wire [28:0] x336_1 ;
 wire [28:0] x337 ;
 wire [28:0] x337_1 ;
 wire [28:0] x338 ;
 wire [28:0] x338_1 ;
 wire [28:0] x339 ;
 wire [28:0] x339_1 ;
 wire [28:0] x340 ;
 wire [28:0] x340_1 ;
 wire [28:0] x341 ;
 wire [28:0] x341_1 ;
 wire [28:0] x342 ;
 wire [28:0] x342_1 ;
 wire [28:0] x343 ;
 wire [28:0] x343_1 ;
 wire [28:0] x344 ;
 wire [28:0] x344_1 ;
 wire [28:0] x345 ;
 wire [28:0] x345_1 ;
 wire [28:0] x346 ;
 wire [28:0] x346_1 ;
 wire [28:0] x347 ;
 wire [28:0] x347_1 ;
 wire [28:0] x348 ;
 wire [28:0] x348_1 ;
 wire [28:0] x349 ;
 wire [28:0] x349_1 ;
 wire [28:0] x350 ;
 wire [28:0] x350_1 ;
 wire [28:0] x351 ;
 wire [28:0] x351_1 ;
 wire [28:0] x352 ;
 wire [28:0] x352_1 ;
 wire [28:0] x353 ;
 wire [28:0] x353_1 ;
 wire [28:0] x354 ;
 wire [28:0] x354_1 ;
 wire [28:0] x355 ;
 wire [28:0] x355_1 ;
 wire [28:0] x356 ;
 wire [28:0] x356_1 ;
 wire [28:0] x357 ;
 wire [28:0] x357_1 ;
 wire [28:0] x358 ;
 wire [28:0] x358_1 ;
 wire [28:0] x359 ;
 wire [28:0] x359_1 ;
 wire [28:0] x360 ;
 wire [28:0] x360_1 ;
 wire [28:0] x361 ;
 wire [28:0] x361_1 ;
 wire [28:0] x362 ;
 wire [28:0] x362_1 ;
 wire [28:0] x363 ;
 wire [28:0] x363_1 ;
 wire [28:0] x364 ;
 wire [28:0] x364_1 ;
 wire [28:0] x365 ;
 wire [28:0] x365_1 ;
 wire [28:0] x366 ;
 wire [28:0] x366_1 ;
 wire [28:0] x367 ;
 wire [28:0] x367_1 ;
 wire [28:0] x368 ;
 wire [28:0] x368_1 ;
 wire [28:0] x369 ;
 wire [28:0] x369_1 ;
 wire [28:0] x370 ;
 wire [28:0] x370_1 ;
 wire [28:0] x371 ;
 wire [28:0] x371_1 ;
 wire [28:0] x372 ;
 wire [28:0] x372_1 ;
 wire [28:0] Out_Y_wire ;
 reg [28:0] Out_Y;


 always @(posedge clk) 
 begin
 x0 <= In_X; 
 end 


 always @(posedge clk) 
 begin
 Out_Y = Out_Y_wire;
 end


 Subtractor14Bit Sub0(clk, {x0[11],x0[11], x0[11: 0] },  { x0[11: 0], 2'b0 },x1); 


 Adder17Bit Adder0(clk,  {x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] },  { x1[14: 0], 2'b0 },x6); 


 Adder24Bit Adder1(clk,  {x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0] },  { x6[17: 0], 6'b0 },x59); 

 Negator25Bit Neg0(clk, x59, x117 );
 Register25Bit Reg0 (clk,x117, y96 );
 Register25Bit Reg1 (clk,x117, y153 );
 Negator18Bit Neg1(clk, x6, x102 );
 Register18Bit Reg2 (clk,x102, x102_0_1 );
 Register21Bit Reg3 (clk, {x102_0_1, 3'b0}, y41 );
 Register18Bit Reg4 (clk,x102, x102_1_1 );
 Register19Bit Reg5 (clk, {x102_1_1, 1'b0}, y52 );
 Register18Bit Reg6 (clk,x102, x102_2_1 );
 Register19Bit Reg7 (clk, {x102_2_1, 1'b0}, y197 );
 Register18Bit Reg8 (clk,x102, x102_3_1 );
 Register21Bit Reg9 (clk, {x102_3_1, 3'b0}, y208 );
 Register18Bit Reg10 (clk,x6, x6_4_1 );
 Register18Bit Reg11 (clk,x6_4_1, x6_4_2 );
 Register18Bit Reg12 (clk,x6_4_2, y3 );
 Register18Bit Reg13 (clk,x6, x6_5_1 );
 Register18Bit Reg14 (clk,x6_5_1, x6_5_2 );
 Register18Bit Reg15 (clk,x6_5_2, y246 );

 Adder18Bit Adder2(clk,  {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] },  { x1[14: 0], 3'b0 },x14); 


 Subtractor22Bit Sub1(clk, { x1[14: 0], 7'b0 }, {x14[18],x14[18],x14[18], x14[18: 0] }, x64); 

 Register23Bit Reg16 (clk,x64, x64_0_1 );
 Register25Bit Reg17 (clk, {x64_0_1, 2'b0}, y110 );
 Register23Bit Reg18 (clk,x64, x64_1_1 );
 Register25Bit Reg19 (clk, {x64_1_1, 2'b0}, y139 );
 Negator19Bit Neg2(clk, x14, x96 );
 Register19Bit Reg20 (clk,x96, x96_0_1 );
 Register19Bit Reg21 (clk,x96_0_1, y17 );
 Register19Bit Reg22 (clk,x96, x96_1_1 );
 Register19Bit Reg23 (clk,x96_1_1, y232 );

 Subtractor16Bit Sub2(clk, { x0[11: 0], 4'b0 }, {x1[14], x1[14: 0] }, x15); 

 Register17Bit Reg24 (clk,x15, x15_0_1 );
 Register17Bit Reg25 (clk,x15_0_1, x15_0_2 );
 Register17Bit Reg26 (clk,x15_0_2, y26 );
 Register17Bit Reg27 (clk,x15, x15_1_1 );
 Register17Bit Reg28 (clk,x15_1_1, x15_1_2 );
 Register17Bit Reg29 (clk,x15_1_2, y34 );
 Register17Bit Reg30 (clk,x15, x15_2_1 );
 Register17Bit Reg31 (clk,x15_2_1, x15_2_2 );
 Register17Bit Reg32 (clk,x15_2_2, y215 );
 Register17Bit Reg33 (clk,x15, x15_3_1 );
 Register17Bit Reg34 (clk,x15_3_1, x15_3_2 );
 Register17Bit Reg35 (clk,x15_3_2, y223 );

 Subtractor21Bit Sub3(clk, {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] },  { x1[14: 0], 6'b0 },x16); 

 Negator22Bit Neg3(clk, x16, x118 );
 Register22Bit Reg36 (clk,x118, x118_0_1 );
 Register22Bit Reg37 (clk,x118_0_1, y105 );
 Register22Bit Reg38 (clk,x118, x118_1_1 );
 Register22Bit Reg39 (clk,x118_1_1, y144 );
 Register22Bit Reg40 (clk,x16, x16_1_1 );
 Register22Bit Reg41 (clk,x16_1_1, x16_1_2 );
 Register22Bit Reg42 (clk,x16_1_2, y65 );
 Register22Bit Reg43 (clk,x16, x16_2_1 );
 Register22Bit Reg44 (clk,x16_2_1, x16_2_2 );
 Register22Bit Reg45 (clk,x16_2_2, y184 );

 Subtractor20Bit Sub4(clk, { x1[14: 0], 5'b0 }, {x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0] }, x20); 

 Register21Bit Reg46 (clk,x20, x20_0_1 );
 Register21Bit Reg47 (clk,x20_0_1, x20_0_2 );
 Register22Bit Reg48 (clk, {x20_0_2, 1'b0}, y63 );
 Register21Bit Reg49 (clk,x20, x20_1_1 );
 Register21Bit Reg50 (clk,x20_1_1, x20_1_2 );
 Register21Bit Reg51 (clk,x20_1_2, y95 );
 Register21Bit Reg52 (clk,x20, x20_2_1 );
 Register21Bit Reg53 (clk,x20_2_1, x20_2_2 );
 Register21Bit Reg54 (clk,x20_2_2, y154 );
 Register21Bit Reg55 (clk,x20, x20_3_1 );
 Register21Bit Reg56 (clk,x20_3_1, x20_3_2 );
 Register22Bit Reg57 (clk, {x20_3_2, 1'b0}, y186 );

 Adder17Bit Adder3(clk,  { x0[11: 0], 5'b0 }, {x1[14],x1[14], x1[14: 0]  }, x27); 

 Register18Bit Reg58 (clk,x27, x27_0_1 );
 Register18Bit Reg59 (clk,x27_0_1, x27_0_2 );
 Register18Bit Reg60 (clk,x27_0_2, y21 );
 Register18Bit Reg61 (clk,x27, x27_1_1 );
 Register18Bit Reg62 (clk,x27_1_1, x27_1_2 );
 Register18Bit Reg63 (clk,x27_1_2, y228 );

 Adder19Bit Adder4(clk,  {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] },  { x1[14: 0], 4'b0 },x28); 

 Negator20Bit Neg4(clk, x28, x100 );
 Register20Bit Reg64 (clk,x100, x100_0_1 );
 Register20Bit Reg65 (clk,x100_0_1, y29 );
 Register20Bit Reg66 (clk,x100, x100_1_1 );
 Register20Bit Reg67 (clk,x100_1_1, y220 );

 Subtractor18Bit Sub5(clk, {x1[14],x1[14],x1[14], x1[14: 0] },  { x0[11: 0], 6'b0 },x29); 

 Register19Bit Reg68 (clk,x29, x29_0_1 );
 Register19Bit Reg69 (clk,x29_0_1, x29_0_2 );
 Register19Bit Reg70 (clk,x29_0_2, y35 );
 Register19Bit Reg71 (clk,x29, x29_1_1 );
 Register19Bit Reg72 (clk,x29_1_1, x29_1_2 );
 Register19Bit Reg73 (clk,x29_1_2, y214 );

 Subtractor20Bit Sub6(clk, { x1[14: 0], 5'b0 }, {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] }, x30); 

 Register21Bit Reg74 (clk,x30, x30_0_1 );
 Register21Bit Reg75 (clk,x30_0_1, x30_0_2 );
 Register21Bit Reg76 (clk,x30_0_2, y43 );
 Register21Bit Reg77 (clk,x30, x30_1_1 );
 Register21Bit Reg78 (clk,x30_1_1, x30_1_2 );
 Register21Bit Reg79 (clk,x30_1_2, y206 );

 Subtractor17Bit Sub7(clk, { x0[11: 0], 5'b0 }, {x1[14],x1[14], x1[14: 0] }, x31); 

 Register18Bit Reg80 (clk,x31, x31_0_1 );
 Register18Bit Reg81 (clk,x31_0_1, x31_0_2 );
 Register19Bit Reg82 (clk, {x31_0_2, 1'b0}, y60 );
 Register18Bit Reg83 (clk,x31, x31_1_1 );
 Register18Bit Reg84 (clk,x31_1_1, x31_1_2 );
 Register19Bit Reg85 (clk, {x31_1_2, 1'b0}, y189 );

 Adder19Bit Adder5(clk,  { x0[11: 0], 7'b0 }, {x1[14],x1[14],x1[14],x1[14], x1[14: 0]  }, x32); 

 Register20Bit Reg86 (clk,x32, x32_0_1 );
 Register20Bit Reg87 (clk,x32_0_1, x32_0_2 );
 Register21Bit Reg88 (clk, {x32_0_2, 1'b0}, y76 );
 Register20Bit Reg89 (clk,x32, x32_1_1 );
 Register20Bit Reg90 (clk,x32_1_1, x32_1_2 );
 Register21Bit Reg91 (clk, {x32_1_2, 1'b0}, y173 );

 Subtractor23Bit Sub8(clk, { x1[14: 0], 8'b0 }, {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] }, x33); 


 Subtractor20Bit Sub9(clk, { x0[11: 0], 8'b0 }, {x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0] }, x34); 

 Register21Bit Reg92 (clk,x34, x34_0_1 );
 Register21Bit Reg93 (clk,x34_0_1, x34_0_2 );
 Register23Bit Reg94 (clk, {x34_0_2, 2'b0}, y104 );
 Register21Bit Reg95 (clk,x34, x34_1_1 );
 Register21Bit Reg96 (clk,x34_1_1, x34_1_2 );
 Register23Bit Reg97 (clk, {x34_1_2, 2'b0}, y145 );

 Subtractor19Bit Sub10(clk, { x1[14: 0], 4'b0 }, {x1[14],x1[14],x1[14],x1[14], x1[14: 0] }, x46); 

 Register20Bit Reg98 (clk,x46, x46_0_1 );
 Register20Bit Reg99 (clk,x46_0_1, x46_0_2 );
 Register20Bit Reg100 (clk,x46_0_2, y101 );
 Register20Bit Reg101 (clk,x46, x46_1_1 );
 Register20Bit Reg102 (clk,x46_1_1, x46_1_2 );
 Register20Bit Reg103 (clk,x46_1_2, y148 );
 Negator15Bit Neg5(clk, x1, x92 );
 Register15Bit Reg104 (clk,x92, x92_0_1 );
 Register15Bit Reg105 (clk,x92_0_1, x92_0_2 );
 Register17Bit Reg106 (clk, {x92_0_2, 2'b0}, y5 );
 Register15Bit Reg107 (clk,x92, x92_1_1 );
 Register15Bit Reg108 (clk,x92_1_1, x92_1_2 );
 Register17Bit Reg109 (clk, {x92_1_2, 2'b0}, y14 );
 Register15Bit Reg110 (clk,x92, x92_2_1 );
 Register15Bit Reg111 (clk,x92_2_1, x92_2_2 );
 Register16Bit Reg112 (clk, {x92_2_2, 1'b0}, y48 );
 Register15Bit Reg113 (clk,x92, x92_3_1 );
 Register15Bit Reg114 (clk,x92_3_1, x92_3_2 );
 Register21Bit Reg115 (clk, {x92_3_2, 6'b0}, y72 );
 Register15Bit Reg116 (clk,x92, x92_4_1 );
 Register15Bit Reg117 (clk,x92_4_1, x92_4_2 );
 Register21Bit Reg118 (clk, {x92_4_2, 6'b0}, y177 );
 Register15Bit Reg119 (clk,x92, x92_5_1 );
 Register15Bit Reg120 (clk,x92_5_1, x92_5_2 );
 Register16Bit Reg121 (clk, {x92_5_2, 1'b0}, y201 );
 Register15Bit Reg122 (clk,x92, x92_6_1 );
 Register15Bit Reg123 (clk,x92_6_1, x92_6_2 );
 Register17Bit Reg124 (clk, {x92_6_2, 2'b0}, y235 );
 Register15Bit Reg125 (clk,x92, x92_7_1 );
 Register15Bit Reg126 (clk,x92_7_1, x92_7_2 );
 Register17Bit Reg127 (clk, {x92_7_2, 2'b0}, y244 );
 Register15Bit Reg128 (clk,x1, x1_42_1 );
 Register15Bit Reg129 (clk,x1_42_1, x1_42_2 );
 Register15Bit Reg130 (clk,x1_42_2, x1_42_3 );
 Register15Bit Reg131 (clk,x1_42_3, y4 );
 Register15Bit Reg132 (clk,x1, x1_43_1 );
 Register15Bit Reg133 (clk,x1_43_1, x1_43_2 );
 Register15Bit Reg134 (clk,x1_43_2, x1_43_3 );
 Register17Bit Reg135 (clk, {x1_43_3, 2'b0}, y12 );
 Register15Bit Reg136 (clk,x1, x1_44_1 );
 Register15Bit Reg137 (clk,x1_44_1, x1_44_2 );
 Register15Bit Reg138 (clk,x1_44_2, x1_44_3 );
 Register16Bit Reg139 (clk, {x1_44_3, 1'b0}, y44 );
 Register15Bit Reg140 (clk,x1, x1_45_1 );
 Register15Bit Reg141 (clk,x1_45_1, x1_45_2 );
 Register15Bit Reg142 (clk,x1_45_2, x1_45_3 );
 Register16Bit Reg143 (clk, {x1_45_3, 1'b0}, y205 );
 Register15Bit Reg144 (clk,x1, x1_46_1 );
 Register15Bit Reg145 (clk,x1_46_1, x1_46_2 );
 Register15Bit Reg146 (clk,x1_46_2, x1_46_3 );
 Register17Bit Reg147 (clk, {x1_46_3, 2'b0}, y237 );
 Register15Bit Reg148 (clk,x1, x1_47_1 );
 Register15Bit Reg149 (clk,x1_47_1, x1_47_2 );
 Register15Bit Reg150 (clk,x1_47_2, x1_47_3 );
 Register15Bit Reg151 (clk,x1_47_3, y245 );

 Adder14Bit Adder6(clk,  {x0[11],x0[11], x0[11: 0] },  { x0[11: 0], 2'b0 },x2); 


 Adder17Bit Adder7(clk,  {x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] },  { x2[14: 0], 2'b0 },x7); 


 Subtractor23Bit Sub11(clk, { x1[14: 0], 8'b0 }, {x7[17],x7[17],x7[17],x7[17],x7[17], x7[17: 0] }, x60); 

 Register24Bit Reg152 (clk,x60, x60_0_1 );
 Register25Bit Reg153 (clk, {x60_0_1, 1'b0}, y117 );
 Register24Bit Reg154 (clk,x60, x60_1_1 );
 Register25Bit Reg155 (clk, {x60_1_1, 1'b0}, y132 );
 Negator18Bit Neg6(clk, x7, x95 );
 Register18Bit Reg156 (clk,x95, x95_0_1 );
 Register18Bit Reg157 (clk,x95_0_1, y15 );
 Register18Bit Reg158 (clk,x95, x95_1_1 );
 Register18Bit Reg159 (clk,x95_1_1, y28 );
 Register18Bit Reg160 (clk,x95, x95_2_1 );
 Register21Bit Reg161 (clk, {x95_2_1, 3'b0}, y70 );
 Register18Bit Reg162 (clk,x95, x95_3_1 );
 Register21Bit Reg163 (clk, {x95_3_1, 3'b0}, y179 );
 Register18Bit Reg164 (clk,x95, x95_4_1 );
 Register18Bit Reg165 (clk,x95_4_1, y221 );
 Register18Bit Reg166 (clk,x95, x95_5_1 );
 Register18Bit Reg167 (clk,x95_5_1, y234 );
 Register18Bit Reg168 (clk,x7, x7_10_1 );
 Register18Bit Reg169 (clk,x7_10_1, x7_10_2 );
 Register21Bit Reg170 (clk, {x7_10_2, 3'b0}, y89 );
 Register18Bit Reg171 (clk,x7, x7_11_1 );
 Register18Bit Reg172 (clk,x7_11_1, x7_11_2 );
 Register21Bit Reg173 (clk, {x7_11_2, 3'b0}, y160 );

 Subtractor17Bit Sub12(clk, {x2[14],x2[14], x2[14: 0] },  { x0[11: 0], 5'b0 },x9); 


 Adder25Bit Adder8(clk,  {x6[17],x6[17],x6[17],x6[17],x6[17],x6[17],x6[17], x6[17: 0] },  { x9[17: 0], 7'b0 },x76); 

 Register26Bit Reg174 (clk,x76, x76_0_1 );
 Register27Bit Reg175 (clk, {x76_0_1, 1'b0}, y122 );
 Register26Bit Reg176 (clk,x76, x76_1_1 );
 Register27Bit Reg177 (clk, {x76_1_1, 1'b0}, y127 );
 Register18Bit Reg178 (clk,x9, x9_7_1 );
 Register18Bit Reg179 (clk,x9_7_1, x9_7_2 );
 Register18Bit Reg180 (clk,x9_7_2, y19 );
 Register18Bit Reg181 (clk,x9, x9_8_1 );
 Register18Bit Reg182 (clk,x9_8_1, x9_8_2 );
 Register19Bit Reg183 (clk, {x9_8_2, 1'b0}, y31 );
 Register18Bit Reg184 (clk,x9, x9_9_1 );
 Register18Bit Reg185 (clk,x9_9_1, x9_9_2 );
 Register19Bit Reg186 (clk, {x9_9_2, 1'b0}, y218 );
 Register18Bit Reg187 (clk,x9, x9_10_1 );
 Register18Bit Reg188 (clk,x9_10_1, x9_10_2 );
 Register18Bit Reg189 (clk,x9_10_2, y230 );

 Adder19Bit Adder9(clk,  { x1[14: 0], 4'b0 }, {x2[14],x2[14],x2[14],x2[14], x2[14: 0]  }, x10); 


 Subtractor21Bit Sub13(clk, { x0[11: 0], 9'b0 }, {x10[19], x10[19: 0] }, x45); 

 Register22Bit Reg190 (clk,x45, x45_0_1 );
 Register23Bit Reg191 (clk, {x45_0_1, 1'b0}, y115 );
 Register22Bit Reg192 (clk,x45, x45_1_1 );
 Register23Bit Reg193 (clk, {x45_1_1, 1'b0}, y134 );
 Negator20Bit Neg7(clk, x10, x105 );
 Register20Bit Reg194 (clk,x105, x105_0_1 );
 Register20Bit Reg195 (clk,x105_0_1, y56 );
 Register20Bit Reg196 (clk,x105, x105_1_1 );
 Register20Bit Reg197 (clk,x105_1_1, y193 );
 Register20Bit Reg198 (clk,x10, x10_2_1 );
 Register20Bit Reg199 (clk,x10_2_1, x10_2_2 );
 Register20Bit Reg200 (clk,x10_2_2, y27 );
 Register20Bit Reg201 (clk,x10, x10_3_1 );
 Register20Bit Reg202 (clk,x10_3_1, x10_3_2 );
 Register20Bit Reg203 (clk,x10_3_2, y222 );

 Subtractor19Bit Sub14(clk, { x1[14: 0], 4'b0 }, {x2[14],x2[14],x2[14],x2[14], x2[14: 0] }, x11); 


 Subtractor24Bit Sub15(clk, {x2[14],x2[14],x2[14],x2[14],x2[14],x2[14],x2[14],x2[14],x2[14], x2[14: 0] },  { x11[19: 0], 4'b0 },x70); 

 Register25Bit Reg204 (clk,x70, x70_0_1 );
 Register25Bit Reg205 (clk,x70_0_1, y100 );
 Register25Bit Reg206 (clk,x70, x70_1_1 );
 Register25Bit Reg207 (clk,x70_1_1, y149 );
 Negator20Bit Neg8(clk, x11, x111 );
 Register20Bit Reg208 (clk,x111, x111_0_1 );
 Register22Bit Reg209 (clk, {x111_0_1, 2'b0}, y81 );
 Register20Bit Reg210 (clk,x111, x111_1_1 );
 Register22Bit Reg211 (clk, {x111_1_1, 2'b0}, y168 );
 Register20Bit Reg212 (clk,x11, x11_2_1 );
 Register20Bit Reg213 (clk,x11_2_1, x11_2_2 );
 Register22Bit Reg214 (clk, {x11_2_2, 2'b0}, y71 );
 Register20Bit Reg215 (clk,x11, x11_3_1 );
 Register20Bit Reg216 (clk,x11_3_1, x11_3_2 );
 Register22Bit Reg217 (clk, {x11_3_2, 2'b0}, y178 );

 Adder17Bit Adder10(clk,  { x0[11: 0], 5'b0 }, {x2[14],x2[14], x2[14: 0]  }, x17); 

 Register18Bit Reg218 (clk,x17, x17_1_1 );
 Register18Bit Reg219 (clk,x17_1_1, x17_1_2 );
 Register18Bit Reg220 (clk,x17_1_2, y25 );
 Register18Bit Reg221 (clk,x17, x17_2_1 );
 Register18Bit Reg222 (clk,x17_2_1, x17_2_2 );
 Register18Bit Reg223 (clk,x17_2_2, y224 );

 Subtractor19Bit Sub16(clk, { x0[11: 0], 7'b0 }, {x2[14],x2[14],x2[14],x2[14], x2[14: 0] }, x18); 

 Register20Bit Reg224 (clk,x18, x18_0_1 );
 Register20Bit Reg225 (clk,x18_0_1, x18_0_2 );
 Register20Bit Reg226 (clk,x18_0_2, y49 );
 Register20Bit Reg227 (clk,x18, x18_1_1 );
 Register20Bit Reg228 (clk,x18_1_1, x18_1_2 );
 Register20Bit Reg229 (clk,x18_1_2, y93 );
 Register20Bit Reg230 (clk,x18, x18_2_1 );
 Register20Bit Reg231 (clk,x18_2_1, x18_2_2 );
 Register20Bit Reg232 (clk,x18_2_2, y156 );
 Register20Bit Reg233 (clk,x18, x18_3_1 );
 Register20Bit Reg234 (clk,x18_3_1, x18_3_2 );
 Register20Bit Reg235 (clk,x18_3_2, y200 );

 Subtractor18Bit Sub17(clk, { x0[11: 0], 6'b0 }, {x2[14],x2[14],x2[14], x2[14: 0] }, x35); 

 Register19Bit Reg236 (clk,x35, x35_0_1 );
 Register19Bit Reg237 (clk,x35_0_1, x35_0_2 );
 Register19Bit Reg238 (clk,x35_0_2, y33 );
 Register19Bit Reg239 (clk,x35, x35_1_1 );
 Register19Bit Reg240 (clk,x35_1_1, x35_1_2 );
 Register19Bit Reg241 (clk,x35_1_2, y216 );

 Adder19Bit Adder11(clk,  {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] },  { x2[14: 0], 4'b0 },x36); 

 Negator20Bit Neg9(clk, x36, x101 );
 Register20Bit Reg242 (clk,x101, x101_0_1 );
 Register20Bit Reg243 (clk,x101_0_1, y39 );
 Register20Bit Reg244 (clk,x101, x101_1_1 );
 Register20Bit Reg245 (clk,x101_1_1, y210 );

 Adder19Bit Adder12(clk,  { x0[11: 0], 7'b0 }, {x2[14],x2[14],x2[14],x2[14], x2[14: 0]  }, x37); 

 Negator20Bit Neg10(clk, x37, x103 );
 Register20Bit Reg246 (clk,x103, x103_0_1 );
 Register20Bit Reg247 (clk,x103_0_1, y51 );
 Register20Bit Reg248 (clk,x103, x103_1_1 );
 Register20Bit Reg249 (clk,x103_1_1, y198 );

 Subtractor19Bit Sub18(clk, { x2[14: 0], 4'b0 }, {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] }, x38); 

 Register20Bit Reg250 (clk,x38, x38_0_1 );
 Register20Bit Reg251 (clk,x38_0_1, x38_0_2 );
 Register22Bit Reg252 (clk, {x38_0_2, 2'b0}, y80 );
 Register20Bit Reg253 (clk,x38, x38_1_1 );
 Register20Bit Reg254 (clk,x38_1_1, x38_1_2 );
 Register22Bit Reg255 (clk, {x38_1_2, 2'b0}, y169 );

 Adder23Bit Adder13(clk,  {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] },  { x2[14: 0], 8'b0 },x39); 

 Register24Bit Reg256 (clk,x39, x39_0_1 );
 Register24Bit Reg257 (clk,x39_0_1, x39_0_2 );
 Register24Bit Reg258 (clk,x39_0_2, y108 );
 Register24Bit Reg259 (clk,x39, x39_1_1 );
 Register24Bit Reg260 (clk,x39_1_1, x39_1_2 );
 Register24Bit Reg261 (clk,x39_1_2, y141 );

 Subtractor21Bit Sub19(clk, {x2[14],x2[14],x2[14],x2[14],x2[14],x2[14], x2[14: 0] },  { x1[14: 0], 6'b0 },x47); 

 Register22Bit Reg262 (clk,x47, x47_0_1 );
 Register22Bit Reg263 (clk,x47_0_1, x47_0_2 );
 Register22Bit Reg264 (clk,x47_0_2, y85 );
 Register22Bit Reg265 (clk,x47, x47_1_1 );
 Register22Bit Reg266 (clk,x47_1_1, x47_1_2 );
 Register22Bit Reg267 (clk,x47_1_2, y164 );

 Adder25Bit Adder14(clk,  {x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0] },  { x2[14: 0], 10'b0 },x48); 

 Register26Bit Reg268 (clk,x48, x48_0_1 );
 Register26Bit Reg269 (clk,x48_0_1, x48_0_2 );
 Register27Bit Reg270 (clk, {x48_0_2, 1'b0}, y123 );
 Register26Bit Reg271 (clk,x48, x48_1_1 );
 Register26Bit Reg272 (clk,x48_1_1, x48_1_2 );
 Register27Bit Reg273 (clk, {x48_1_2, 1'b0}, y126 );

 Adder19Bit Adder15(clk,  {x2[14],x2[14],x2[14],x2[14], x2[14: 0] },  { x2[14: 0], 4'b0 },x67); 

 Negator20Bit Neg11(clk, x67, x107 );
 Register20Bit Reg274 (clk,x107, x107_0_1 );
 Register21Bit Reg275 (clk, {x107_0_1, 1'b0}, y59 );
 Register20Bit Reg276 (clk,x107, x107_1_1 );
 Register21Bit Reg277 (clk, {x107_1_1, 1'b0}, y190 );

 Adder22Bit Adder16(clk,  {x2[14],x2[14],x2[14],x2[14],x2[14],x2[14],x2[14], x2[14: 0] },  { x2[14: 0], 7'b0 },x68); 

 Negator23Bit Neg12(clk, x68, x116 );
 Register23Bit Reg278 (clk,x116, x116_0_1 );
 Register23Bit Reg279 (clk,x116_0_1, y94 );
 Register23Bit Reg280 (clk,x116, x116_1_1 );
 Register23Bit Reg281 (clk,x116_1_1, y155 );

 Adder24Bit Adder17(clk,  {x2[14],x2[14],x2[14],x2[14],x2[14],x2[14], x2[14: 0], 3'b0 }, { x33[23: 0]  }, x71); 

 Register25Bit Reg282 (clk,x71, x71_0_1 );
 Register27Bit Reg283 (clk, {x71_0_1, 2'b0}, y118 );
 Register25Bit Reg284 (clk,x71, x71_1_1 );
 Register27Bit Reg285 (clk, {x71_1_1, 2'b0}, y131 );
 Negator15Bit Neg13(clk, x2, x99 );
 Register15Bit Reg286 (clk,x99, x99_0_1 );
 Register15Bit Reg287 (clk,x99_0_1, x99_0_2 );
 Register17Bit Reg288 (clk, {x99_0_2, 2'b0}, y24 );
 Register15Bit Reg289 (clk,x99, x99_1_1 );
 Register15Bit Reg290 (clk,x99_1_1, x99_1_2 );
 Register17Bit Reg291 (clk, {x99_1_2, 2'b0}, y32 );
 Register15Bit Reg292 (clk,x99, x99_2_1 );
 Register15Bit Reg293 (clk,x99_2_1, x99_2_2 );
 Register16Bit Reg294 (clk, {x99_2_2, 1'b0}, y99 );
 Register15Bit Reg295 (clk,x99, x99_3_1 );
 Register15Bit Reg296 (clk,x99_3_1, x99_3_2 );
 Register16Bit Reg297 (clk, {x99_3_2, 1'b0}, y150 );
 Register15Bit Reg298 (clk,x99, x99_4_1 );
 Register15Bit Reg299 (clk,x99_4_1, x99_4_2 );
 Register17Bit Reg300 (clk, {x99_4_2, 2'b0}, y217 );
 Register15Bit Reg301 (clk,x99, x99_5_1 );
 Register15Bit Reg302 (clk,x99_5_1, x99_5_2 );
 Register17Bit Reg303 (clk, {x99_5_2, 2'b0}, y225 );
 Register15Bit Reg304 (clk,x2, x2_21_1 );
 Register15Bit Reg305 (clk,x2_21_1, x2_21_2 );
 Register15Bit Reg306 (clk,x2_21_2, x2_21_3 );
 Register15Bit Reg307 (clk,x2_21_3, y0 );
 Register15Bit Reg308 (clk,x2, x2_22_1 );
 Register15Bit Reg309 (clk,x2_22_1, x2_22_2 );
 Register15Bit Reg310 (clk,x2_22_2, x2_22_3 );
 Register15Bit Reg311 (clk,x2_22_3, y6 );
 Register15Bit Reg312 (clk,x2, x2_23_1 );
 Register15Bit Reg313 (clk,x2_23_1, x2_23_2 );
 Register15Bit Reg314 (clk,x2_23_2, x2_23_3 );
 Register17Bit Reg315 (clk, {x2_23_3, 2'b0}, y30 );
 Register15Bit Reg316 (clk,x2, x2_24_1 );
 Register15Bit Reg317 (clk,x2_24_1, x2_24_2 );
 Register15Bit Reg318 (clk,x2_24_2, x2_24_3 );
 Register20Bit Reg319 (clk, {x2_24_3, 5'b0}, y57 );
 Register15Bit Reg320 (clk,x2, x2_25_1 );
 Register15Bit Reg321 (clk,x2_25_1, x2_25_2 );
 Register15Bit Reg322 (clk,x2_25_2, x2_25_3 );
 Register20Bit Reg323 (clk, {x2_25_3, 5'b0}, y192 );
 Register15Bit Reg324 (clk,x2, x2_26_1 );
 Register15Bit Reg325 (clk,x2_26_1, x2_26_2 );
 Register15Bit Reg326 (clk,x2_26_2, x2_26_3 );
 Register17Bit Reg327 (clk, {x2_26_3, 2'b0}, y219 );
 Register15Bit Reg328 (clk,x2, x2_27_1 );
 Register15Bit Reg329 (clk,x2_27_1, x2_27_2 );
 Register15Bit Reg330 (clk,x2_27_2, x2_27_3 );
 Register15Bit Reg331 (clk,x2_27_3, y243 );
 Register15Bit Reg332 (clk,x2, x2_28_1 );
 Register15Bit Reg333 (clk,x2_28_1, x2_28_2 );
 Register15Bit Reg334 (clk,x2_28_2, x2_28_3 );
 Register15Bit Reg335 (clk,x2_28_3, y249 );

 Adder15Bit Adder18(clk,  {x0[11],x0[11],x0[11], x0[11: 0] },  { x0[11: 0], 3'b0 },x3); 


 Adder19Bit Adder19(clk,  {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] },  { x3[15: 0], 3'b0 },x19); 

 Register20Bit Reg336 (clk,x19, x19_0_1 );
 Register20Bit Reg337 (clk,x19_0_1, x19_0_2 );
 Register20Bit Reg338 (clk,x19_0_2, y37 );
 Register20Bit Reg339 (clk,x19, x19_1_1 );
 Register20Bit Reg340 (clk,x19_1_1, x19_1_2 );
 Register22Bit Reg341 (clk, {x19_1_2, 2'b0}, y107 );
 Register20Bit Reg342 (clk,x19, x19_2_1 );
 Register20Bit Reg343 (clk,x19_2_1, x19_2_2 );
 Register22Bit Reg344 (clk, {x19_2_2, 2'b0}, y142 );
 Register20Bit Reg345 (clk,x19, x19_3_1 );
 Register20Bit Reg346 (clk,x19_3_1, x19_3_2 );
 Register20Bit Reg347 (clk,x19_3_2, y212 );

 Subtractor20Bit Sub20(clk, {x3[15],x3[15],x3[15],x3[15], x3[15: 0] },  { x1[14: 0], 5'b0 },x21); 

 Negator21Bit Neg14(clk, x21, x120 );
 Register21Bit Reg348 (clk,x120, x120_0_1 );
 Register23Bit Reg349 (clk, {x120_0_1, 2'b0}, y109 );
 Register21Bit Reg350 (clk,x120, x120_1_1 );
 Register23Bit Reg351 (clk, {x120_1_1, 2'b0}, y140 );
 Register21Bit Reg352 (clk,x21, x21_1_1 );
 Register21Bit Reg353 (clk,x21_1_1, x21_1_2 );
 Register21Bit Reg354 (clk,x21_1_2, y45 );
 Register21Bit Reg355 (clk,x21, x21_2_1 );
 Register21Bit Reg356 (clk,x21_2_1, x21_2_2 );
 Register21Bit Reg357 (clk,x21_2_2, y204 );

 Subtractor18Bit Sub21(clk, { x0[11: 0], 6'b0 }, {x3[15],x3[15], x3[15: 0] }, x40); 

 Register19Bit Reg358 (clk,x40, x40_0_1 );
 Register19Bit Reg359 (clk,x40_0_1, x40_0_2 );
 Register19Bit Reg360 (clk,x40_0_2, y97 );
 Register19Bit Reg361 (clk,x40, x40_1_1 );
 Register19Bit Reg362 (clk,x40_1_1, x40_1_2 );
 Register19Bit Reg363 (clk,x40_1_2, y152 );

 Adder20Bit Adder20(clk,  { x1[14: 0], 5'b0 }, {x3[15],x3[15],x3[15],x3[15], x3[15: 0]  }, x49); 

 Register21Bit Reg364 (clk,x49, x49_0_1 );
 Register21Bit Reg365 (clk,x49_0_1, x49_0_2 );
 Register21Bit Reg366 (clk,x49_0_2, y62 );
 Register21Bit Reg367 (clk,x49, x49_1_1 );
 Register21Bit Reg368 (clk,x49_1_1, x49_1_2 );
 Register21Bit Reg369 (clk,x49_1_2, y187 );

 Subtractor21Bit Sub22(clk, { x1[14: 0], 6'b0 }, {x3[15],x3[15],x3[15],x3[15],x3[15], x3[15: 0] }, x50); 

 Register22Bit Reg370 (clk,x50, x50_0_1 );
 Register22Bit Reg371 (clk,x50_0_1, x50_0_2 );
 Register22Bit Reg372 (clk,x50_0_2, y67 );
 Register22Bit Reg373 (clk,x50, x50_1_1 );
 Register22Bit Reg374 (clk,x50_1_1, x50_1_2 );
 Register22Bit Reg375 (clk,x50_1_2, y182 );

 Subtractor22Bit Sub23(clk, {x3[15],x3[15],x3[15],x3[15],x3[15],x3[15], x3[15: 0] },  { x1[14: 0], 7'b0 },x51); 

 Register23Bit Reg376 (clk,x51, x51_0_1 );
 Register23Bit Reg377 (clk,x51_0_1, x51_0_2 );
 Register23Bit Reg378 (clk,x51_0_2, y84 );
 Register23Bit Reg379 (clk,x51, x51_1_1 );
 Register23Bit Reg380 (clk,x51_1_1, x51_1_2 );
 Register23Bit Reg381 (clk,x51_1_2, y165 );

 Subtractor23Bit Sub24(clk, { x1[14: 0], 8'b0 }, {x3[15],x3[15],x3[15],x3[15],x3[15],x3[15],x3[15], x3[15: 0] }, x52); 

 Register24Bit Reg382 (clk,x52, x52_0_1 );
 Register24Bit Reg383 (clk,x52_0_1, x52_0_2 );
 Register24Bit Reg384 (clk,x52_0_2, y98 );
 Register24Bit Reg385 (clk,x52, x52_1_1 );
 Register24Bit Reg386 (clk,x52_1_1, x52_1_2 );
 Register24Bit Reg387 (clk,x52_1_2, y151 );

 Adder23Bit Adder21(clk,  {x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0] },  { x3[15: 0], 7'b0 },x53); 

 Negator24Bit Neg15(clk, x53, x119 );
 Register24Bit Reg388 (clk,x119, x119_0_1 );
 Register24Bit Reg389 (clk,x119_0_1, y106 );
 Register24Bit Reg390 (clk,x119, x119_1_1 );
 Register24Bit Reg391 (clk,x119_1_1, y143 );

 Subtractor24Bit Sub25(clk, { x3[15: 0], 8'b0 }, {x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0] }, x54); 

 Register25Bit Reg392 (clk,x54, x54_0_1 );
 Register25Bit Reg393 (clk,x54_0_1, x54_0_2 );
 Register25Bit Reg394 (clk,x54_0_2, y116 );
 Register25Bit Reg395 (clk,x54, x54_1_1 );
 Register25Bit Reg396 (clk,x54_1_1, x54_1_2 );
 Register25Bit Reg397 (clk,x54_1_2, y133 );

 Subtractor21Bit Sub26(clk, {x2[14],x2[14],x2[14],x2[14],x2[14],x2[14], x2[14: 0] },  { x3[15: 0], 5'b0 },x69); 

 Register22Bit Reg398 (clk,x69, x69_0_1 );
 Register22Bit Reg399 (clk,x69_0_1, x69_0_2 );
 Register22Bit Reg400 (clk,x69_0_2, y78 );
 Register22Bit Reg401 (clk,x69, x69_1_1 );
 Register22Bit Reg402 (clk,x69_1_1, x69_1_2 );
 Register22Bit Reg403 (clk,x69_1_2, y171 );

 Adder22Bit Adder22(clk,  {x3[15],x3[15],x3[15],x3[15],x3[15],x3[15], x3[15: 0] },  { x3[15: 0], 6'b0 },x72); 

 Register23Bit Reg404 (clk,x72, x72_0_1 );
 Register23Bit Reg405 (clk,x72_0_1, x72_0_2 );
 Register23Bit Reg406 (clk,x72_0_2, y92 );
 Register23Bit Reg407 (clk,x72, x72_1_1 );
 Register23Bit Reg408 (clk,x72_1_1, x72_1_2 );
 Register23Bit Reg409 (clk,x72_1_2, y157 );
 Negator16Bit Neg16(clk, x3, x98 );
 Register16Bit Reg410 (clk,x98, x98_0_1 );
 Register16Bit Reg411 (clk,x98_0_1, x98_0_2 );
 Register17Bit Reg412 (clk, {x98_0_2, 1'b0}, y20 );
 Register16Bit Reg413 (clk,x98, x98_1_1 );
 Register16Bit Reg414 (clk,x98_1_1, x98_1_2 );
 Register17Bit Reg415 (clk, {x98_1_2, 1'b0}, y36 );
 Register16Bit Reg416 (clk,x98, x98_2_1 );
 Register16Bit Reg417 (clk,x98_2_1, x98_2_2 );
 Register17Bit Reg418 (clk, {x98_2_2, 1'b0}, y213 );
 Register16Bit Reg419 (clk,x98, x98_3_1 );
 Register16Bit Reg420 (clk,x98_3_1, x98_3_2 );
 Register17Bit Reg421 (clk, {x98_3_2, 1'b0}, y229 );
 Register16Bit Reg422 (clk,x3, x3_14_1 );
 Register16Bit Reg423 (clk,x3_14_1, x3_14_2 );
 Register16Bit Reg424 (clk,x3_14_2, x3_14_3 );
 Register16Bit Reg425 (clk,x3_14_3, y10 );
 Register16Bit Reg426 (clk,x3, x3_15_1 );
 Register16Bit Reg427 (clk,x3_15_1, x3_15_2 );
 Register16Bit Reg428 (clk,x3_15_2, x3_15_3 );
 Register17Bit Reg429 (clk, {x3_15_3, 1'b0}, y13 );
 Register16Bit Reg430 (clk,x3, x3_16_1 );
 Register16Bit Reg431 (clk,x3_16_1, x3_16_2 );
 Register16Bit Reg432 (clk,x3_16_2, x3_16_3 );
 Register17Bit Reg433 (clk, {x3_16_3, 1'b0}, y22 );
 Register16Bit Reg434 (clk,x3, x3_17_1 );
 Register16Bit Reg435 (clk,x3_17_1, x3_17_2 );
 Register16Bit Reg436 (clk,x3_17_2, x3_17_3 );
 Register16Bit Reg437 (clk,x3_17_3, y42 );
 Register16Bit Reg438 (clk,x3, x3_18_1 );
 Register16Bit Reg439 (clk,x3_18_1, x3_18_2 );
 Register16Bit Reg440 (clk,x3_18_2, x3_18_3 );
 Register20Bit Reg441 (clk, {x3_18_3, 4'b0}, y68 );
 Register16Bit Reg442 (clk,x3, x3_19_1 );
 Register16Bit Reg443 (clk,x3_19_1, x3_19_2 );
 Register16Bit Reg444 (clk,x3_19_2, x3_19_3 );
 Register20Bit Reg445 (clk, {x3_19_3, 4'b0}, y181 );
 Register16Bit Reg446 (clk,x3, x3_20_1 );
 Register16Bit Reg447 (clk,x3_20_1, x3_20_2 );
 Register16Bit Reg448 (clk,x3_20_2, x3_20_3 );
 Register16Bit Reg449 (clk,x3_20_3, y207 );
 Register16Bit Reg450 (clk,x3, x3_21_1 );
 Register16Bit Reg451 (clk,x3_21_1, x3_21_2 );
 Register16Bit Reg452 (clk,x3_21_2, x3_21_3 );
 Register17Bit Reg453 (clk, {x3_21_3, 1'b0}, y227 );
 Register16Bit Reg454 (clk,x3, x3_22_1 );
 Register16Bit Reg455 (clk,x3_22_1, x3_22_2 );
 Register16Bit Reg456 (clk,x3_22_2, x3_22_3 );
 Register17Bit Reg457 (clk, {x3_22_3, 1'b0}, y236 );
 Register16Bit Reg458 (clk,x3, x3_23_1 );
 Register16Bit Reg459 (clk,x3_23_1, x3_23_2 );
 Register16Bit Reg460 (clk,x3_23_2, x3_23_3 );
 Register16Bit Reg461 (clk,x3_23_3, y239 );

 Subtractor15Bit Sub27(clk, { x0[11: 0], 3'b0 }, {x0[11],x0[11],x0[11], x0[11: 0] }, x4); 


 Subtractor20Bit Sub28(clk, {x4[15],x4[15],x4[15],x4[15], x4[15: 0] },  { x1[14: 0], 5'b0 },x12); 

 Register21Bit Reg462 (clk,x12, x12_0_1 );
 Register21Bit Reg463 (clk,x12_0_1, x12_0_2 );
 Register21Bit Reg464 (clk,x12_0_2, y64 );
 Register21Bit Reg465 (clk,x12, x12_1_1 );
 Register21Bit Reg466 (clk,x12_1_1, x12_1_2 );
 Register22Bit Reg467 (clk, {x12_1_2, 1'b0}, y69 );
 Register21Bit Reg468 (clk,x12, x12_2_1 );
 Register21Bit Reg469 (clk,x12_2_1, x12_2_2 );
 Register25Bit Reg470 (clk, {x12_2_2, 4'b0}, y112 );
 Register21Bit Reg471 (clk,x12, x12_3_1 );
 Register21Bit Reg472 (clk,x12_3_1, x12_3_2 );
 Register25Bit Reg473 (clk, {x12_3_2, 4'b0}, y137 );
 Register21Bit Reg474 (clk,x12, x12_4_1 );
 Register21Bit Reg475 (clk,x12_4_1, x12_4_2 );
 Register22Bit Reg476 (clk, {x12_4_2, 1'b0}, y180 );
 Register21Bit Reg477 (clk,x12, x12_5_1 );
 Register21Bit Reg478 (clk,x12_5_1, x12_5_2 );
 Register21Bit Reg479 (clk,x12_5_2, y185 );

 Adder19Bit Adder23(clk,  {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] },  { x4[15: 0], 3'b0 },x41); 

 Negator20Bit Neg17(clk, x41, x106 );
 Register20Bit Reg480 (clk,x106, x106_0_1 );
 Register20Bit Reg481 (clk,x106_0_1, y58 );
 Register20Bit Reg482 (clk,x106, x106_1_1 );
 Register20Bit Reg483 (clk,x106_1_1, y191 );

 Subtractor20Bit Sub29(clk, { x4[15: 0], 4'b0 }, {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] }, x42); 

 Register21Bit Reg484 (clk,x42, x42_0_1 );
 Register21Bit Reg485 (clk,x42_0_1, x42_0_2 );
 Register21Bit Reg486 (clk,x42_0_2, y103 );
 Register21Bit Reg487 (clk,x42, x42_1_1 );
 Register21Bit Reg488 (clk,x42_1_1, x42_1_2 );
 Register21Bit Reg489 (clk,x42_1_2, y146 );

 Adder21Bit Adder24(clk,  {x1[14],x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0] },  { x4[15: 0], 5'b0 },x55); 

 Negator22Bit Neg18(clk, x55, x109 );
 Register22Bit Reg490 (clk,x109, x109_0_1 );
 Register22Bit Reg491 (clk,x109_0_1, y74 );
 Register22Bit Reg492 (clk,x109, x109_1_1 );
 Register22Bit Reg493 (clk,x109_1_1, y175 );

 Adder20Bit Adder25(clk,  {x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0] },  { x4[15: 0], 4'b0 },x56); 

 Negator21Bit Neg19(clk, x56, x110 );
 Register21Bit Reg494 (clk,x110, x110_0_1 );
 Register22Bit Reg495 (clk, {x110_0_1, 1'b0}, y75 );
 Register21Bit Reg496 (clk,x110, x110_1_1 );
 Register22Bit Reg497 (clk, {x110_1_1, 1'b0}, y174 );

 Adder21Bit Adder26(clk,  { x1[14: 0], 6'b0 }, {x4[15],x4[15],x4[15],x4[15],x4[15], x4[15: 0]  }, x57); 

 Register22Bit Reg498 (clk,x57, x57_0_1 );
 Register22Bit Reg499 (clk,x57_0_1, x57_0_2 );
 Register22Bit Reg500 (clk,x57_0_2, y87 );
 Register22Bit Reg501 (clk,x57, x57_1_1 );
 Register22Bit Reg502 (clk,x57_1_1, x57_1_2 );
 Register22Bit Reg503 (clk,x57_1_2, y162 );

 Adder22Bit Adder27(clk,  { x3[15: 0], 6'b0 }, {x4[15],x4[15],x4[15],x4[15],x4[15],x4[15], x4[15: 0]  }, x73); 

 Register23Bit Reg504 (clk,x73, x73_0_1 );
 Register23Bit Reg505 (clk,x73_0_1, x73_0_2 );
 Register23Bit Reg506 (clk,x73_0_2, y111 );
 Register23Bit Reg507 (clk,x73, x73_1_1 );
 Register23Bit Reg508 (clk,x73_1_1, x73_1_2 );
 Register23Bit Reg509 (clk,x73_1_2, y138 );

 Adder22Bit Adder28(clk,  { x4[15: 0], 6'b0 }, {x6[17],x6[17],x6[17],x6[17], x6[17: 0]  }, x74); 

 Negator23Bit Neg20(clk, x74, x113 );
 Register23Bit Reg510 (clk,x113, y86 );
 Register23Bit Reg511 (clk,x113, y163 );

 Adder24Bit Adder29(clk,  {x4[15],x4[15],x4[15],x4[15],x4[15],x4[15],x4[15],x4[15], x4[15: 0] },  { x17[17: 0], 6'b0 },x75); 

 Register25Bit Reg512 (clk,x75, x75_0_1 );
 Register25Bit Reg513 (clk,x75_0_1, y119 );
 Register25Bit Reg514 (clk,x75, x75_1_1 );
 Register25Bit Reg515 (clk,x75_1_1, y130 );
 Negator16Bit Neg21(clk, x4, x93 );
 Register16Bit Reg516 (clk,x93, x93_0_1 );
 Register16Bit Reg517 (clk,x93_0_1, x93_0_2 );
 Register17Bit Reg518 (clk, {x93_0_2, 1'b0}, y7 );
 Register16Bit Reg519 (clk,x93, x93_1_1 );
 Register16Bit Reg520 (clk,x93_1_1, x93_1_2 );
 Register17Bit Reg521 (clk, {x93_1_2, 1'b0}, y40 );
 Register16Bit Reg522 (clk,x93, x93_2_1 );
 Register16Bit Reg523 (clk,x93_2_1, x93_2_2 );
 Register17Bit Reg524 (clk, {x93_2_2, 1'b0}, y50 );
 Register16Bit Reg525 (clk,x93, x93_3_1 );
 Register16Bit Reg526 (clk,x93_3_1, x93_3_2 );
 Register17Bit Reg527 (clk, {x93_3_2, 1'b0}, y199 );
 Register16Bit Reg528 (clk,x93, x93_4_1 );
 Register16Bit Reg529 (clk,x93_4_1, x93_4_2 );
 Register17Bit Reg530 (clk, {x93_4_2, 1'b0}, y209 );
 Register16Bit Reg531 (clk,x93, x93_5_1 );
 Register16Bit Reg532 (clk,x93_5_1, x93_5_2 );
 Register17Bit Reg533 (clk, {x93_5_2, 1'b0}, y242 );
 Register16Bit Reg534 (clk,x4, x4_10_1 );
 Register16Bit Reg535 (clk,x4_10_1, x4_10_2 );
 Register16Bit Reg536 (clk,x4_10_2, x4_10_3 );
 Register16Bit Reg537 (clk,x4_10_3, y1 );
 Register16Bit Reg538 (clk,x4, x4_11_1 );
 Register16Bit Reg539 (clk,x4_11_1, x4_11_2 );
 Register16Bit Reg540 (clk,x4_11_2, x4_11_3 );
 Register17Bit Reg541 (clk, {x4_11_3, 1'b0}, y9 );
 Register16Bit Reg542 (clk,x4, x4_12_1 );
 Register16Bit Reg543 (clk,x4_12_1, x4_12_2 );
 Register16Bit Reg544 (clk,x4_12_2, x4_12_3 );
 Register17Bit Reg545 (clk, {x4_12_3, 1'b0}, y240 );
 Register16Bit Reg546 (clk,x4, x4_13_1 );
 Register16Bit Reg547 (clk,x4_13_1, x4_13_2 );
 Register16Bit Reg548 (clk,x4_13_2, x4_13_3 );
 Register16Bit Reg549 (clk,x4_13_3, y248 );

 Subtractor16Bit Sub30(clk, {x0[11],x0[11],x0[11],x0[11], x0[11: 0] },  { x0[11: 0], 4'b0 },x5); 


 Subtractor21Bit Sub31(clk, {x5[16],x5[16],x5[16],x5[16], x5[16: 0] },  { x1[14: 0], 6'b0 },x22); 

 Negator22Bit Neg22(clk, x22, x112 );
 Register22Bit Reg550 (clk,x112, x112_0_1 );
 Register23Bit Reg551 (clk, {x112_0_1, 1'b0}, y82 );
 Register22Bit Reg552 (clk,x112, x112_1_1 );
 Register23Bit Reg553 (clk, {x112_1_1, 1'b0}, y167 );
 Register22Bit Reg554 (clk,x22, x22_1_1 );
 Register22Bit Reg555 (clk,x22_1_1, x22_1_2 );
 Register22Bit Reg556 (clk,x22_1_2, y61 );
 Register22Bit Reg557 (clk,x22, x22_2_1 );
 Register22Bit Reg558 (clk,x22_2_1, x22_2_2 );
 Register22Bit Reg559 (clk,x22_2_2, y188 );

 Subtractor21Bit Sub32(clk, {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] },  { x5[16: 0], 4'b0 },x43); 

 Register22Bit Reg560 (clk,x43, x43_0_1 );
 Register22Bit Reg561 (clk,x43_0_1, x43_0_2 );
 Register23Bit Reg562 (clk, {x43_0_2, 1'b0}, y88 );
 Register22Bit Reg563 (clk,x43, x43_1_1 );
 Register22Bit Reg564 (clk,x43_1_1, x43_1_2 );
 Register23Bit Reg565 (clk, {x43_1_2, 1'b0}, y161 );

 Subtractor24Bit Sub33(clk, { x5[16: 0], 7'b0 }, {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] }, x44); 

 Register25Bit Reg566 (clk,x44, x44_0_1 );
 Register25Bit Reg567 (clk,x44_0_1, x44_0_2 );
 Register25Bit Reg568 (clk,x44_0_2, y114 );
 Register25Bit Reg569 (clk,x44, x44_1_1 );
 Register25Bit Reg570 (clk,x44_1_1, x44_1_2 );
 Register25Bit Reg571 (clk,x44_1_2, y135 );

 Adder21Bit Adder30(clk,  { x1[14: 0], 6'b0 }, {x5[16],x5[16],x5[16],x5[16], x5[16: 0]  }, x58); 

 Register22Bit Reg572 (clk,x58, x58_0_1 );
 Register22Bit Reg573 (clk,x58_0_1, x58_0_2 );
 Register22Bit Reg574 (clk,x58_0_2, y83 );
 Register22Bit Reg575 (clk,x58, x58_1_1 );
 Register22Bit Reg576 (clk,x58_1_1, x58_1_2 );
 Register22Bit Reg577 (clk,x58_1_2, y166 );
 Negator17Bit Neg23(clk, x5, x97 );
 Register17Bit Reg578 (clk,x97, x97_0_1 );
 Register17Bit Reg579 (clk,x97_0_1, x97_0_2 );
 Register17Bit Reg580 (clk,x97_0_2, y18 );
 Register17Bit Reg581 (clk,x97, x97_1_1 );
 Register17Bit Reg582 (clk,x97_1_1, x97_1_2 );
 Register17Bit Reg583 (clk,x97_1_2, y38 );
 Register17Bit Reg584 (clk,x97, x97_2_1 );
 Register17Bit Reg585 (clk,x97_2_1, x97_2_2 );
 Register17Bit Reg586 (clk,x97_2_2, y211 );
 Register17Bit Reg587 (clk,x97, x97_3_1 );
 Register17Bit Reg588 (clk,x97_3_1, x97_3_2 );
 Register17Bit Reg589 (clk,x97_3_2, y231 );
 Register17Bit Reg590 (clk,x5, x5_5_1 );
 Register17Bit Reg591 (clk,x5_5_1, x5_5_2 );
 Register17Bit Reg592 (clk,x5_5_2, x5_5_3 );
 Register17Bit Reg593 (clk,x5_5_3, y16 );
 Register17Bit Reg594 (clk,x5, x5_6_1 );
 Register17Bit Reg595 (clk,x5_6_1, x5_6_2 );
 Register17Bit Reg596 (clk,x5_6_2, x5_6_3 );
 Register17Bit Reg597 (clk,x5_6_3, y233 );

 Adder16Bit Adder31(clk,  {x0[11],x0[11],x0[11],x0[11], x0[11: 0] },  { x0[11: 0], 4'b0 },x8); 


 Subtractor22Bit Sub34(clk, { x1[14: 0], 7'b0 }, {x8[16],x8[16],x8[16],x8[16],x8[16], x8[16: 0] }, x61); 

 Register23Bit Reg598 (clk,x61, x61_0_1 );
 Register23Bit Reg599 (clk,x61_0_1, x61_0_2 );
 Register24Bit Reg600 (clk, {x61_0_2, 1'b0}, y113 );
 Register23Bit Reg601 (clk,x61, x61_1_1 );
 Register23Bit Reg602 (clk,x61_1_1, x61_1_2 );
 Register24Bit Reg603 (clk, {x61_1_2, 1'b0}, y136 );
 Negator17Bit Neg24(clk, x8, x94 );
 Register17Bit Reg604 (clk,x94, x94_0_1 );
 Register17Bit Reg605 (clk,x94_0_1, x94_0_2 );
 Register17Bit Reg606 (clk,x94_0_2, y11 );
 Register17Bit Reg607 (clk,x94, x94_1_1 );
 Register17Bit Reg608 (clk,x94_1_1, x94_1_2 );
 Register18Bit Reg609 (clk, {x94_1_2, 1'b0}, y23 );
 Register17Bit Reg610 (clk,x94, x94_2_1 );
 Register17Bit Reg611 (clk,x94_2_1, x94_2_2 );
 Register18Bit Reg612 (clk, {x94_2_2, 1'b0}, y226 );
 Register17Bit Reg613 (clk,x94, x94_3_1 );
 Register17Bit Reg614 (clk,x94_3_1, x94_3_2 );
 Register17Bit Reg615 (clk,x94_3_2, y238 );

 Subtractor19Bit Sub35(clk, {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] },  { x0[11: 0], 7'b0 },x13); 


 Subtractor20Bit Sub36(clk, { x13[19: 0] },  {x1[14],x1[14],x1[14], x1[14: 0], 2'b0 },x62); 

 Register21Bit Reg616 (clk,x62, x62_0_1 );
 Register21Bit Reg617 (clk,x62_0_1, x62_0_2 );
 Register21Bit Reg618 (clk,x62_0_2, y47 );
 Register21Bit Reg619 (clk,x62, x62_1_1 );
 Register21Bit Reg620 (clk,x62_1_1, x62_1_2 );
 Register21Bit Reg621 (clk,x62_1_2, y202 );

 Adder20Bit Adder32(clk,  {x1[14],x1[14], x1[14: 0], 3'b0 }, { x13[19: 0]  }, x63); 

 Register21Bit Reg622 (clk,x63, x63_0_1 );
 Register21Bit Reg623 (clk,x63_0_1, x63_0_2 );
 Register21Bit Reg624 (clk,x63_0_2, y55 );
 Register21Bit Reg625 (clk,x63, x63_1_1 );
 Register21Bit Reg626 (clk,x63_1_1, x63_1_2 );
 Register21Bit Reg627 (clk,x63_1_2, y194 );

 Subtractor17Bit Sub37(clk, { x0[11: 0], 5'b0 }, {x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] }, x23); 

 Negator18Bit Neg25(clk, x23, x108 );
 Register18Bit Reg628 (clk,x108, x108_0_1 );
 Register18Bit Reg629 (clk,x108_0_1, x108_0_2 );
 Register20Bit Reg630 (clk, {x108_0_2, 2'b0}, y66 );
 Register18Bit Reg631 (clk,x108, x108_1_1 );
 Register18Bit Reg632 (clk,x108_1_1, x108_1_2 );
 Register20Bit Reg633 (clk, {x108_1_2, 2'b0}, y183 );

 Adder17Bit Adder33(clk,  {x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] },  { x0[11: 0], 5'b0 },x24); 

 Negator18Bit Neg26(clk, x24, x104 );
 Register18Bit Reg634 (clk,x104, x104_0_1 );
 Register18Bit Reg635 (clk,x104_0_1, x104_0_2 );
 Register18Bit Reg636 (clk,x104_0_2, y54 );
 Register18Bit Reg637 (clk,x104, x104_1_1 );
 Register18Bit Reg638 (clk,x104_1_1, x104_1_2 );
 Register18Bit Reg639 (clk,x104_1_2, y195 );

 Adder19Bit Adder34(clk,  {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] },  { x0[11: 0], 7'b0 },x25); 


 Subtractor20Bit Sub38(clk, { x25[19: 0] },  {x1[14],x1[14],x1[14], x1[14: 0], 2'b0 },x65); 

 Register21Bit Reg640 (clk,x65, x65_0_1 );
 Register21Bit Reg641 (clk,x65_0_1, x65_0_2 );
 Register21Bit Reg642 (clk,x65_0_2, y53 );
 Register21Bit Reg643 (clk,x65, x65_1_1 );
 Register21Bit Reg644 (clk,x65_1_1, x65_1_2 );
 Register21Bit Reg645 (clk,x65_1_2, y196 );

 Subtractor23Bit Sub39(clk, { x0[11: 0], 11'b0 }, {x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11],x0[11], x0[11: 0] }, x26); 


 Adder24Bit Adder35(clk,  {x1[14],x1[14],x1[14],x1[14],x1[14],x1[14],x1[14], x1[14: 0], 2'b0 }, { x26[23: 0]  }, x66); 

 Negator25Bit Neg27(clk, x66, x121 );
 Register25Bit Reg646 (clk,x121, x121_0_1 );
 Register26Bit Reg647 (clk, {x121_0_1, 1'b0}, y121 );
 Register25Bit Reg648 (clk,x121, x121_1_1 );
 Register26Bit Reg649 (clk, {x121_1_1, 1'b0}, y128 );
 Register12Bit Reg650 (clk,x0, x77_50_1 );
 Register12Bit Reg651 (clk,x77_50_1, x77_50_2 );

 Subtractor19Bit Sub40(clk, { x77_50_2[11: 0], 7'b0 }, {x7[17], x7[17: 0] }, x77); 

 Register20Bit Reg652 (clk,x77, x77_0_1 );
 Register21Bit Reg653 (clk, {x77_0_1, 1'b0}, y73 );
 Register12Bit Reg654 (clk,x0, x78_51_1 );
 Register12Bit Reg655 (clk,x78_51_1, x78_51_2 );

 Subtractor21Bit Sub41(clk, {x78_51_2[11],x78_51_2[11],x78_51_2[11],x78_51_2[11],x78_51_2[11],x78_51_2[11],x78_51_2[11],x78_51_2[11],x78_51_2[11], x78_51_2[11: 0] },  { x9[17: 0], 3'b0 },x78); 

 Register22Bit Reg656 (clk,x78, x78_0_1 );
 Register22Bit Reg657 (clk,x78_0_1, y77 );
 Register12Bit Reg658 (clk,x0, x79_52_1 );
 Register12Bit Reg659 (clk,x79_52_1, x79_52_2 );

 Subtractor21Bit Sub42(clk, { x9[17: 0], 3'b0 }, {x79_52_2[11],x79_52_2[11],x79_52_2[11],x79_52_2[11],x79_52_2[11],x79_52_2[11],x79_52_2[11],x79_52_2[11],x79_52_2[11], x79_52_2[11: 0] }, x79); 

 Register22Bit Reg660 (clk,x79, x79_0_1 );
 Register22Bit Reg661 (clk,x79_0_1, y79 );
 Register12Bit Reg662 (clk,x0, x80_53_1 );
 Register12Bit Reg663 (clk,x80_53_1, x80_53_2 );

 Adder21Bit Adder36(clk,  { x80_53_2[11: 0], 9'b0 }, {x7[17],x7[17],x7[17], x7[17: 0]  }, x80); 

 Negator22Bit Neg28(clk, x80, x114 );
 Register22Bit Reg664 (clk,x114, y90 );
 Register12Bit Reg665 (clk,x0, x81_54_1 );
 Register12Bit Reg666 (clk,x81_54_1, x81_54_2 );

 Adder19Bit Adder37(clk,  { x81_54_2[11: 0], 7'b0 }, {x7[17], x7[17: 0]  }, x81); 

 Negator20Bit Neg29(clk, x81, x115 );
 Register20Bit Reg667 (clk,x115, y91 );
 Register12Bit Reg668 (clk,x0, x82_55_1 );
 Register12Bit Reg669 (clk,x82_55_1, x82_55_2 );

 Subtractor20Bit Sub43(clk, {x7[17],x7[17], x7[17: 0] },  { x82_55_2[11: 0], 8'b0 },x82); 

 Register21Bit Reg670 (clk,x82, x82_0_1 );
 Register23Bit Reg671 (clk, {x82_0_1, 2'b0}, y102 );
 Register12Bit Reg672 (clk,x0, x83_56_1 );
 Register12Bit Reg673 (clk,x83_56_1, x83_56_2 );

 Adder23Bit Adder38(clk,  { x83_56_2[11: 0], 11'b0 }, {x9[17],x9[17],x9[17],x9[17],x9[17], x9[17: 0]  }, x83); 

 Register24Bit Reg674 (clk,x83, x83_0_1 );
 Register25Bit Reg675 (clk, {x83_0_1, 1'b0}, y120 );
 Register12Bit Reg676 (clk,x0, x84_57_1 );
 Register12Bit Reg677 (clk,x84_57_1, x84_57_2 );

 Adder23Bit Adder39(clk,  { x84_57_2[11: 0], 11'b0 }, {x9[17],x9[17],x9[17],x9[17],x9[17], x9[17: 0]  }, x84); 

 Register24Bit Reg678 (clk,x84, x84_0_1 );
 Register25Bit Reg679 (clk, {x84_0_1, 1'b0}, y129 );
 Register12Bit Reg680 (clk,x0, x85_58_1 );
 Register12Bit Reg681 (clk,x85_58_1, x85_58_2 );

 Subtractor20Bit Sub44(clk, {x7[17],x7[17], x7[17: 0] },  { x85_58_2[11: 0], 8'b0 },x85); 

 Register21Bit Reg682 (clk,x85, x85_0_1 );
 Register23Bit Reg683 (clk, {x85_0_1, 2'b0}, y147 );
 Register12Bit Reg684 (clk,x0, x86_59_1 );
 Register12Bit Reg685 (clk,x86_59_1, x86_59_2 );

 Adder19Bit Adder40(clk,  { x86_59_2[11: 0], 7'b0 }, {x7[17], x7[17: 0]  }, x86); 

 Negator20Bit Neg30(clk, x86, x122 );
 Register20Bit Reg686 (clk,x122, y158 );
 Register12Bit Reg687 (clk,x0, x87_60_1 );
 Register12Bit Reg688 (clk,x87_60_1, x87_60_2 );

 Adder21Bit Adder41(clk,  { x87_60_2[11: 0], 9'b0 }, {x7[17],x7[17],x7[17], x7[17: 0]  }, x87); 

 Negator22Bit Neg31(clk, x87, x123 );
 Register22Bit Reg689 (clk,x123, y159 );
 Register12Bit Reg690 (clk,x0, x88_61_1 );
 Register12Bit Reg691 (clk,x88_61_1, x88_61_2 );

 Subtractor21Bit Sub45(clk, { x9[17: 0], 3'b0 }, {x88_61_2[11],x88_61_2[11],x88_61_2[11],x88_61_2[11],x88_61_2[11],x88_61_2[11],x88_61_2[11],x88_61_2[11],x88_61_2[11], x88_61_2[11: 0] }, x88); 

 Register22Bit Reg692 (clk,x88, x88_0_1 );
 Register22Bit Reg693 (clk,x88_0_1, y170 );
 Register12Bit Reg694 (clk,x0, x89_62_1 );
 Register12Bit Reg695 (clk,x89_62_1, x89_62_2 );

 Subtractor21Bit Sub46(clk, {x89_62_2[11],x89_62_2[11],x89_62_2[11],x89_62_2[11],x89_62_2[11],x89_62_2[11],x89_62_2[11],x89_62_2[11],x89_62_2[11], x89_62_2[11: 0] },  { x9[17: 0], 3'b0 },x89); 

 Register22Bit Reg696 (clk,x89, x89_0_1 );
 Register22Bit Reg697 (clk,x89_0_1, y172 );
 Register12Bit Reg698 (clk,x0, x90_63_1 );
 Register12Bit Reg699 (clk,x90_63_1, x90_63_2 );

 Subtractor19Bit Sub47(clk, { x90_63_2[11: 0], 7'b0 }, {x7[17], x7[17: 0] }, x90); 

 Register20Bit Reg700 (clk,x90, x90_0_1 );
 Register21Bit Reg701 (clk, {x90_0_1, 1'b0}, y176 );
 Negator12Bit Neg32(clk, x0, x91 );
 Register12Bit Reg702 (clk,x91, x91_0_1 );
 Register12Bit Reg703 (clk,x91_0_1, x91_0_2 );
 Register12Bit Reg704 (clk,x91_0_2, x91_0_3 );
 Register13Bit Reg705 (clk, {x91_0_3, 1'b0}, y2 );
 Register12Bit Reg706 (clk,x91, x91_1_1 );
 Register12Bit Reg707 (clk,x91_1_1, x91_1_2 );
 Register12Bit Reg708 (clk,x91_1_2, x91_1_3 );
 Register15Bit Reg709 (clk, {x91_1_3, 3'b0}, y8 );
 Register12Bit Reg710 (clk,x91, x91_2_1 );
 Register12Bit Reg711 (clk,x91_2_1, x91_2_2 );
 Register12Bit Reg712 (clk,x91_2_2, x91_2_3 );
 Register12Bit Reg713 (clk,x91_2_3, y46 );
 Register12Bit Reg714 (clk,x91, x91_3_1 );
 Register12Bit Reg715 (clk,x91_3_1, x91_3_2 );
 Register12Bit Reg716 (clk,x91_3_2, x91_3_3 );
 Register12Bit Reg717 (clk,x91_3_3, y203 );
 Register12Bit Reg718 (clk,x91, x91_4_1 );
 Register12Bit Reg719 (clk,x91_4_1, x91_4_2 );
 Register12Bit Reg720 (clk,x91_4_2, x91_4_3 );
 Register15Bit Reg721 (clk, {x91_4_3, 3'b0}, y241 );
 Register12Bit Reg722 (clk,x91, x91_5_1 );
 Register12Bit Reg723 (clk,x91_5_1, x91_5_2 );
 Register12Bit Reg724 (clk,x91_5_2, x91_5_3 );
 Register13Bit Reg725 (clk, {x91_5_3, 1'b0}, y247 );
 Register12Bit Reg726 (clk,x0, x0_65_1 );
 Register12Bit Reg727 (clk,x0_65_1, x0_65_2 );
 Register12Bit Reg728 (clk,x0_65_2, x0_65_3 );
 Register12Bit Reg729 (clk,x0_65_3, x0_65_4 );
 Register27Bit Reg730 (clk, {x0_65_4, 15'b0}, y124 );
 Register12Bit Reg731 (clk,x0, x0_66_1 );
 Register12Bit Reg732 (clk,x0_66_1, x0_66_2 );
 Register12Bit Reg733 (clk,x0_66_2, x0_66_3 );
 Register12Bit Reg734 (clk,x0_66_3, x0_66_4 );
 Register27Bit Reg735 (clk, {x0_66_4, 15'b0}, y125 );
 Register15Bit Reg736 (clk,y0, x124 );

 Adder16Bit Adder42(clk,  {x124[14], x124[14: 0] },  { y1[15: 0]  }, x125); 

 Register17Bit Reg737 (clk,x125, x125_1 );

 Adder17Bit Adder43(clk,  { x125_1[16: 0] },  {y2[12],y2[12],y2[12],y2[12], y2[12: 0]  }, x126); 

 Register18Bit Reg738 (clk,x126, x126_1 );

 Adder18Bit Adder44(clk,  { x126_1[17: 0] },  { y3[17: 0]  }, x127); 

 Register19Bit Reg739 (clk,x127, x127_1 );

 Adder19Bit Adder45(clk,  { x127_1[18: 0] },  {y4[14],y4[14],y4[14],y4[14], y4[14: 0]  }, x128); 

 Register20Bit Reg740 (clk,x128, x128_1 );

 Adder20Bit Adder46(clk,  { x128_1[19: 0] },  {y5[16],y5[16],y5[16], y5[16: 0]  }, x129); 

 Register21Bit Reg741 (clk,x129, x129_1 );

 Adder21Bit Adder47(clk,  { x129_1[20: 0] },  {y6[14],y6[14],y6[14],y6[14],y6[14],y6[14], y6[14: 0]  }, x130); 

 Register22Bit Reg742 (clk,x130, x130_1 );

 Adder22Bit Adder48(clk,  { x130_1[21: 0] },  {y7[16],y7[16],y7[16],y7[16],y7[16], y7[16: 0]  }, x131); 

 Register23Bit Reg743 (clk,x131, x131_1 );

 Adder23Bit Adder49(clk,  { x131_1[22: 0] },  {y8[14],y8[14],y8[14],y8[14],y8[14],y8[14],y8[14],y8[14], y8[14: 0]  }, x132); 

 Register24Bit Reg744 (clk,x132, x132_1 );

 Adder24Bit Adder50(clk,  { x132_1[23: 0] },  {y9[16],y9[16],y9[16],y9[16],y9[16],y9[16],y9[16], y9[16: 0]  }, x133); 

 Register25Bit Reg745 (clk,x133, x133_1 );

 Adder25Bit Adder51(clk,  { x133_1[24: 0] },  {y10[15],y10[15],y10[15],y10[15],y10[15],y10[15],y10[15],y10[15],y10[15], y10[15: 0]  }, x134); 

 Register26Bit Reg746 (clk,x134, x134_1 );

 Adder26Bit Adder52(clk,  { x134_1[25: 0] },  {y11[16],y11[16],y11[16],y11[16],y11[16],y11[16],y11[16],y11[16],y11[16], y11[16: 0]  }, x135); 

 Register27Bit Reg747 (clk,x135, x135_1 );

 Adder27Bit Adder53(clk,  { x135_1[26: 0] },  {y12[16],y12[16],y12[16],y12[16],y12[16],y12[16],y12[16],y12[16],y12[16],y12[16], y12[16: 0]  }, x136); 

 Register28Bit Reg748 (clk,x136, x136_1 );

 Adder28Bit Adder54(clk,  { x136_1[27: 0] },  {y13[16],y13[16],y13[16],y13[16],y13[16],y13[16],y13[16],y13[16],y13[16],y13[16],y13[16], y13[16: 0]  }, x137); 

 Register29Bit Reg749 (clk,x137, x137_1 );

 Adder29Bit Adder55(clk,  { x137_1[28: 0] },  {y14[16],y14[16],y14[16],y14[16],y14[16],y14[16],y14[16],y14[16],y14[16],y14[16],y14[16],y14[16], y14[16: 0]  }, x138); 

 Register29Bit Reg750 (clk,x138, x138_1 );

 Adder29Bit Adder56(clk,  { x138_1[28: 0] },  {y15[17],y15[17],y15[17],y15[17],y15[17],y15[17],y15[17],y15[17],y15[17],y15[17],y15[17], y15[17: 0]  }, x139); 

 Register29Bit Reg751 (clk,x139, x139_1 );

 Adder29Bit Adder57(clk,  { x139_1[28: 0] },  {y16[16],y16[16],y16[16],y16[16],y16[16],y16[16],y16[16],y16[16],y16[16],y16[16],y16[16],y16[16], y16[16: 0]  }, x140); 

 Register29Bit Reg752 (clk,x140, x140_1 );

 Adder29Bit Adder58(clk,  { x140_1[28: 0] },  {y17[18],y17[18],y17[18],y17[18],y17[18],y17[18],y17[18],y17[18],y17[18],y17[18], y17[18: 0]  }, x141); 

 Register29Bit Reg753 (clk,x141, x141_1 );

 Adder29Bit Adder59(clk,  { x141_1[28: 0] },  {y18[16],y18[16],y18[16],y18[16],y18[16],y18[16],y18[16],y18[16],y18[16],y18[16],y18[16],y18[16], y18[16: 0]  }, x142); 

 Register29Bit Reg754 (clk,x142, x142_1 );

 Adder29Bit Adder60(clk,  { x142_1[28: 0] },  {y19[17],y19[17],y19[17],y19[17],y19[17],y19[17],y19[17],y19[17],y19[17],y19[17],y19[17], y19[17: 0]  }, x143); 

 Register29Bit Reg755 (clk,x143, x143_1 );

 Adder29Bit Adder61(clk,  { x143_1[28: 0] },  {y20[16],y20[16],y20[16],y20[16],y20[16],y20[16],y20[16],y20[16],y20[16],y20[16],y20[16],y20[16], y20[16: 0]  }, x144); 

 Register29Bit Reg756 (clk,x144, x144_1 );

 Adder29Bit Adder62(clk,  { x144_1[28: 0] },  {y21[17],y21[17],y21[17],y21[17],y21[17],y21[17],y21[17],y21[17],y21[17],y21[17],y21[17], y21[17: 0]  }, x145); 

 Register29Bit Reg757 (clk,x145, x145_1 );

 Adder29Bit Adder63(clk,  { x145_1[28: 0] },  {y22[16],y22[16],y22[16],y22[16],y22[16],y22[16],y22[16],y22[16],y22[16],y22[16],y22[16],y22[16], y22[16: 0]  }, x146); 

 Register29Bit Reg758 (clk,x146, x146_1 );

 Adder29Bit Adder64(clk,  { x146_1[28: 0] },  {y23[17],y23[17],y23[17],y23[17],y23[17],y23[17],y23[17],y23[17],y23[17],y23[17],y23[17], y23[17: 0]  }, x147); 

 Register29Bit Reg759 (clk,x147, x147_1 );

 Adder29Bit Adder65(clk,  { x147_1[28: 0] },  {y24[16],y24[16],y24[16],y24[16],y24[16],y24[16],y24[16],y24[16],y24[16],y24[16],y24[16],y24[16], y24[16: 0]  }, x148); 

 Register29Bit Reg760 (clk,x148, x148_1 );

 Adder29Bit Adder66(clk,  { x148_1[28: 0] },  {y25[17],y25[17],y25[17],y25[17],y25[17],y25[17],y25[17],y25[17],y25[17],y25[17],y25[17], y25[17: 0]  }, x149); 

 Register29Bit Reg761 (clk,x149, x149_1 );

 Adder29Bit Adder67(clk,  { x149_1[28: 0] },  {y26[16],y26[16],y26[16],y26[16],y26[16],y26[16],y26[16],y26[16],y26[16],y26[16],y26[16],y26[16], y26[16: 0]  }, x150); 

 Register29Bit Reg762 (clk,x150, x150_1 );

 Adder29Bit Adder68(clk,  { x150_1[28: 0] },  {y27[19],y27[19],y27[19],y27[19],y27[19],y27[19],y27[19],y27[19],y27[19], y27[19: 0]  }, x151); 

 Register29Bit Reg763 (clk,x151, x151_1 );

 Adder29Bit Adder69(clk,  { x151_1[28: 0] },  {y28[17],y28[17],y28[17],y28[17],y28[17],y28[17],y28[17],y28[17],y28[17],y28[17],y28[17], y28[17: 0]  }, x152); 

 Register29Bit Reg764 (clk,x152, x152_1 );

 Adder29Bit Adder70(clk,  { x152_1[28: 0] },  {y29[19],y29[19],y29[19],y29[19],y29[19],y29[19],y29[19],y29[19],y29[19], y29[19: 0]  }, x153); 

 Register29Bit Reg765 (clk,x153, x153_1 );

 Adder29Bit Adder71(clk,  { x153_1[28: 0] },  {y30[16],y30[16],y30[16],y30[16],y30[16],y30[16],y30[16],y30[16],y30[16],y30[16],y30[16],y30[16], y30[16: 0]  }, x154); 

 Register29Bit Reg766 (clk,x154, x154_1 );

 Adder29Bit Adder72(clk,  { x154_1[28: 0] },  {y31[18],y31[18],y31[18],y31[18],y31[18],y31[18],y31[18],y31[18],y31[18],y31[18], y31[18: 0]  }, x155); 

 Register29Bit Reg767 (clk,x155, x155_1 );

 Adder29Bit Adder73(clk,  { x155_1[28: 0] },  {y32[16],y32[16],y32[16],y32[16],y32[16],y32[16],y32[16],y32[16],y32[16],y32[16],y32[16],y32[16], y32[16: 0]  }, x156); 

 Register29Bit Reg768 (clk,x156, x156_1 );

 Adder29Bit Adder74(clk,  { x156_1[28: 0] },  {y33[18],y33[18],y33[18],y33[18],y33[18],y33[18],y33[18],y33[18],y33[18],y33[18], y33[18: 0]  }, x157); 

 Register29Bit Reg769 (clk,x157, x157_1 );

 Adder29Bit Adder75(clk,  { x157_1[28: 0] },  {y34[16],y34[16],y34[16],y34[16],y34[16],y34[16],y34[16],y34[16],y34[16],y34[16],y34[16],y34[16], y34[16: 0]  }, x158); 

 Register29Bit Reg770 (clk,x158, x158_1 );

 Adder29Bit Adder76(clk,  { x158_1[28: 0] },  {y35[18],y35[18],y35[18],y35[18],y35[18],y35[18],y35[18],y35[18],y35[18],y35[18], y35[18: 0]  }, x159); 

 Register29Bit Reg771 (clk,x159, x159_1 );

 Adder29Bit Adder77(clk,  { x159_1[28: 0] },  {y36[16],y36[16],y36[16],y36[16],y36[16],y36[16],y36[16],y36[16],y36[16],y36[16],y36[16],y36[16], y36[16: 0]  }, x160); 

 Register29Bit Reg772 (clk,x160, x160_1 );

 Adder29Bit Adder78(clk,  { x160_1[28: 0] },  {y37[19],y37[19],y37[19],y37[19],y37[19],y37[19],y37[19],y37[19],y37[19], y37[19: 0]  }, x161); 

 Register29Bit Reg773 (clk,x161, x161_1 );

 Adder29Bit Adder79(clk,  { x161_1[28: 0] },  {y38[16],y38[16],y38[16],y38[16],y38[16],y38[16],y38[16],y38[16],y38[16],y38[16],y38[16],y38[16], y38[16: 0]  }, x162); 

 Register29Bit Reg774 (clk,x162, x162_1 );

 Adder29Bit Adder80(clk,  { x162_1[28: 0] },  {y39[19],y39[19],y39[19],y39[19],y39[19],y39[19],y39[19],y39[19],y39[19], y39[19: 0]  }, x163); 

 Register29Bit Reg775 (clk,x163, x163_1 );

 Adder29Bit Adder81(clk,  { x163_1[28: 0] },  {y40[16],y40[16],y40[16],y40[16],y40[16],y40[16],y40[16],y40[16],y40[16],y40[16],y40[16],y40[16], y40[16: 0]  }, x164); 

 Register29Bit Reg776 (clk,x164, x164_1 );

 Adder29Bit Adder82(clk,  { x164_1[28: 0] },  {y41[20],y41[20],y41[20],y41[20],y41[20],y41[20],y41[20],y41[20], y41[20: 0]  }, x165); 

 Register29Bit Reg777 (clk,x165, x165_1 );

 Adder29Bit Adder83(clk,  { x165_1[28: 0] },  {y42[15],y42[15],y42[15],y42[15],y42[15],y42[15],y42[15],y42[15],y42[15],y42[15],y42[15],y42[15],y42[15], y42[15: 0]  }, x166); 

 Register29Bit Reg778 (clk,x166, x166_1 );

 Adder29Bit Adder84(clk,  { x166_1[28: 0] },  {y43[20],y43[20],y43[20],y43[20],y43[20],y43[20],y43[20],y43[20], y43[20: 0]  }, x167); 

 Register29Bit Reg779 (clk,x167, x167_1 );

 Adder29Bit Adder85(clk,  { x167_1[28: 0] },  {y44[15],y44[15],y44[15],y44[15],y44[15],y44[15],y44[15],y44[15],y44[15],y44[15],y44[15],y44[15],y44[15], y44[15: 0]  }, x168); 

 Register29Bit Reg780 (clk,x168, x168_1 );

 Adder29Bit Adder86(clk,  { x168_1[28: 0] },  {y45[20],y45[20],y45[20],y45[20],y45[20],y45[20],y45[20],y45[20], y45[20: 0]  }, x169); 

 Register29Bit Reg781 (clk,x169, x169_1 );

 Adder29Bit Adder87(clk,  { x169_1[28: 0] },  {y46[11],y46[11],y46[11],y46[11],y46[11],y46[11],y46[11],y46[11],y46[11],y46[11],y46[11],y46[11],y46[11],y46[11],y46[11],y46[11],y46[11], y46[11: 0]  }, x170); 

 Register29Bit Reg782 (clk,x170, x170_1 );

 Adder29Bit Adder88(clk,  { x170_1[28: 0] },  {y47[20],y47[20],y47[20],y47[20],y47[20],y47[20],y47[20],y47[20], y47[20: 0]  }, x171); 

 Register29Bit Reg783 (clk,x171, x171_1 );

 Adder29Bit Adder89(clk,  { x171_1[28: 0] },  {y48[15],y48[15],y48[15],y48[15],y48[15],y48[15],y48[15],y48[15],y48[15],y48[15],y48[15],y48[15],y48[15], y48[15: 0]  }, x172); 

 Register29Bit Reg784 (clk,x172, x172_1 );

 Adder29Bit Adder90(clk,  { x172_1[28: 0] },  {y49[19],y49[19],y49[19],y49[19],y49[19],y49[19],y49[19],y49[19],y49[19], y49[19: 0]  }, x173); 

 Register29Bit Reg785 (clk,x173, x173_1 );

 Adder29Bit Adder91(clk,  { x173_1[28: 0] },  {y50[16],y50[16],y50[16],y50[16],y50[16],y50[16],y50[16],y50[16],y50[16],y50[16],y50[16],y50[16], y50[16: 0]  }, x174); 

 Register29Bit Reg786 (clk,x174, x174_1 );

 Adder29Bit Adder92(clk,  { x174_1[28: 0] },  {y51[19],y51[19],y51[19],y51[19],y51[19],y51[19],y51[19],y51[19],y51[19], y51[19: 0]  }, x175); 

 Register29Bit Reg787 (clk,x175, x175_1 );

 Adder29Bit Adder93(clk,  { x175_1[28: 0] },  {y52[18],y52[18],y52[18],y52[18],y52[18],y52[18],y52[18],y52[18],y52[18],y52[18], y52[18: 0]  }, x176); 

 Register29Bit Reg788 (clk,x176, x176_1 );

 Adder29Bit Adder94(clk,  { x176_1[28: 0] },  {y53[20],y53[20],y53[20],y53[20],y53[20],y53[20],y53[20],y53[20], y53[20: 0]  }, x177); 

 Register29Bit Reg789 (clk,x177, x177_1 );

 Adder29Bit Adder95(clk,  { x177_1[28: 0] },  {y54[17],y54[17],y54[17],y54[17],y54[17],y54[17],y54[17],y54[17],y54[17],y54[17],y54[17], y54[17: 0]  }, x178); 

 Register29Bit Reg790 (clk,x178, x178_1 );

 Adder29Bit Adder96(clk,  { x178_1[28: 0] },  {y55[20],y55[20],y55[20],y55[20],y55[20],y55[20],y55[20],y55[20], y55[20: 0]  }, x179); 

 Register29Bit Reg791 (clk,x179, x179_1 );

 Adder29Bit Adder97(clk,  { x179_1[28: 0] },  {y56[19],y56[19],y56[19],y56[19],y56[19],y56[19],y56[19],y56[19],y56[19], y56[19: 0]  }, x180); 

 Register29Bit Reg792 (clk,x180, x180_1 );

 Adder29Bit Adder98(clk,  { x180_1[28: 0] },  {y57[19],y57[19],y57[19],y57[19],y57[19],y57[19],y57[19],y57[19],y57[19], y57[19: 0]  }, x181); 

 Register29Bit Reg793 (clk,x181, x181_1 );

 Adder29Bit Adder99(clk,  { x181_1[28: 0] },  {y58[19],y58[19],y58[19],y58[19],y58[19],y58[19],y58[19],y58[19],y58[19], y58[19: 0]  }, x182); 

 Register29Bit Reg794 (clk,x182, x182_1 );

 Adder29Bit Adder100(clk,  { x182_1[28: 0] },  {y59[20],y59[20],y59[20],y59[20],y59[20],y59[20],y59[20],y59[20], y59[20: 0]  }, x183); 

 Register29Bit Reg795 (clk,x183, x183_1 );

 Adder29Bit Adder101(clk,  { x183_1[28: 0] },  {y60[18],y60[18],y60[18],y60[18],y60[18],y60[18],y60[18],y60[18],y60[18],y60[18], y60[18: 0]  }, x184); 

 Register29Bit Reg796 (clk,x184, x184_1 );

 Adder29Bit Adder102(clk,  { x184_1[28: 0] },  {y61[21],y61[21],y61[21],y61[21],y61[21],y61[21],y61[21], y61[21: 0]  }, x185); 

 Register29Bit Reg797 (clk,x185, x185_1 );

 Adder29Bit Adder103(clk,  { x185_1[28: 0] },  {y62[20],y62[20],y62[20],y62[20],y62[20],y62[20],y62[20],y62[20], y62[20: 0]  }, x186); 

 Register29Bit Reg798 (clk,x186, x186_1 );

 Adder29Bit Adder104(clk,  { x186_1[28: 0] },  {y63[21],y63[21],y63[21],y63[21],y63[21],y63[21],y63[21], y63[21: 0]  }, x187); 

 Register29Bit Reg799 (clk,x187, x187_1 );

 Adder29Bit Adder105(clk,  { x187_1[28: 0] },  {y64[20],y64[20],y64[20],y64[20],y64[20],y64[20],y64[20],y64[20], y64[20: 0]  }, x188); 

 Register29Bit Reg800 (clk,x188, x188_1 );

 Adder29Bit Adder106(clk,  { x188_1[28: 0] },  {y65[21],y65[21],y65[21],y65[21],y65[21],y65[21],y65[21], y65[21: 0]  }, x189); 

 Register29Bit Reg801 (clk,x189, x189_1 );

 Adder29Bit Adder107(clk,  { x189_1[28: 0] },  {y66[19],y66[19],y66[19],y66[19],y66[19],y66[19],y66[19],y66[19],y66[19], y66[19: 0]  }, x190); 

 Register29Bit Reg802 (clk,x190, x190_1 );

 Adder29Bit Adder108(clk,  { x190_1[28: 0] },  {y67[21],y67[21],y67[21],y67[21],y67[21],y67[21],y67[21], y67[21: 0]  }, x191); 

 Register29Bit Reg803 (clk,x191, x191_1 );

 Adder29Bit Adder109(clk,  { x191_1[28: 0] },  {y68[19],y68[19],y68[19],y68[19],y68[19],y68[19],y68[19],y68[19],y68[19], y68[19: 0]  }, x192); 

 Register29Bit Reg804 (clk,x192, x192_1 );

 Adder29Bit Adder110(clk,  { x192_1[28: 0] },  {y69[21],y69[21],y69[21],y69[21],y69[21],y69[21],y69[21], y69[21: 0]  }, x193); 

 Register29Bit Reg805 (clk,x193, x193_1 );

 Adder29Bit Adder111(clk,  { x193_1[28: 0] },  {y70[20],y70[20],y70[20],y70[20],y70[20],y70[20],y70[20],y70[20], y70[20: 0]  }, x194); 

 Register29Bit Reg806 (clk,x194, x194_1 );

 Adder29Bit Adder112(clk,  { x194_1[28: 0] },  {y71[21],y71[21],y71[21],y71[21],y71[21],y71[21],y71[21], y71[21: 0]  }, x195); 

 Register29Bit Reg807 (clk,x195, x195_1 );

 Adder29Bit Adder113(clk,  { x195_1[28: 0] },  {y72[20],y72[20],y72[20],y72[20],y72[20],y72[20],y72[20],y72[20], y72[20: 0]  }, x196); 

 Register29Bit Reg808 (clk,x196, x196_1 );

 Adder29Bit Adder114(clk,  { x196_1[28: 0] },  {y73[20],y73[20],y73[20],y73[20],y73[20],y73[20],y73[20],y73[20], y73[20: 0]  }, x197); 

 Register29Bit Reg809 (clk,x197, x197_1 );

 Adder29Bit Adder115(clk,  { x197_1[28: 0] },  {y74[21],y74[21],y74[21],y74[21],y74[21],y74[21],y74[21], y74[21: 0]  }, x198); 

 Register29Bit Reg810 (clk,x198, x198_1 );

 Adder29Bit Adder116(clk,  { x198_1[28: 0] },  {y75[21],y75[21],y75[21],y75[21],y75[21],y75[21],y75[21], y75[21: 0]  }, x199); 

 Register29Bit Reg811 (clk,x199, x199_1 );

 Adder29Bit Adder117(clk,  { x199_1[28: 0] },  {y76[20],y76[20],y76[20],y76[20],y76[20],y76[20],y76[20],y76[20], y76[20: 0]  }, x200); 

 Register29Bit Reg812 (clk,x200, x200_1 );

 Adder29Bit Adder118(clk,  { x200_1[28: 0] },  {y77[21],y77[21],y77[21],y77[21],y77[21],y77[21],y77[21], y77[21: 0]  }, x201); 

 Register29Bit Reg813 (clk,x201, x201_1 );

 Adder29Bit Adder119(clk,  { x201_1[28: 0] },  {y78[21],y78[21],y78[21],y78[21],y78[21],y78[21],y78[21], y78[21: 0]  }, x202); 

 Register29Bit Reg814 (clk,x202, x202_1 );

 Adder29Bit Adder120(clk,  { x202_1[28: 0] },  {y79[21],y79[21],y79[21],y79[21],y79[21],y79[21],y79[21], y79[21: 0]  }, x203); 

 Register29Bit Reg815 (clk,x203, x203_1 );

 Adder29Bit Adder121(clk,  { x203_1[28: 0] },  {y80[21],y80[21],y80[21],y80[21],y80[21],y80[21],y80[21], y80[21: 0]  }, x204); 

 Register29Bit Reg816 (clk,x204, x204_1 );

 Adder29Bit Adder122(clk,  { x204_1[28: 0] },  {y81[21],y81[21],y81[21],y81[21],y81[21],y81[21],y81[21], y81[21: 0]  }, x205); 

 Register29Bit Reg817 (clk,x205, x205_1 );

 Adder29Bit Adder123(clk,  { x205_1[28: 0] },  {y82[22],y82[22],y82[22],y82[22],y82[22],y82[22], y82[22: 0]  }, x206); 

 Register29Bit Reg818 (clk,x206, x206_1 );

 Adder29Bit Adder124(clk,  { x206_1[28: 0] },  {y83[21],y83[21],y83[21],y83[21],y83[21],y83[21],y83[21], y83[21: 0]  }, x207); 

 Register29Bit Reg819 (clk,x207, x207_1 );

 Adder29Bit Adder125(clk,  { x207_1[28: 0] },  {y84[22],y84[22],y84[22],y84[22],y84[22],y84[22], y84[22: 0]  }, x208); 

 Register29Bit Reg820 (clk,x208, x208_1 );

 Adder29Bit Adder126(clk,  { x208_1[28: 0] },  {y85[21],y85[21],y85[21],y85[21],y85[21],y85[21],y85[21], y85[21: 0]  }, x209); 

 Register29Bit Reg821 (clk,x209, x209_1 );

 Adder29Bit Adder127(clk,  { x209_1[28: 0] },  {y86[22],y86[22],y86[22],y86[22],y86[22],y86[22], y86[22: 0]  }, x210); 

 Register29Bit Reg822 (clk,x210, x210_1 );

 Adder29Bit Adder128(clk,  { x210_1[28: 0] },  {y87[21],y87[21],y87[21],y87[21],y87[21],y87[21],y87[21], y87[21: 0]  }, x211); 

 Register29Bit Reg823 (clk,x211, x211_1 );

 Adder29Bit Adder129(clk,  { x211_1[28: 0] },  {y88[22],y88[22],y88[22],y88[22],y88[22],y88[22], y88[22: 0]  }, x212); 

 Register29Bit Reg824 (clk,x212, x212_1 );

 Adder29Bit Adder130(clk,  { x212_1[28: 0] },  {y89[20],y89[20],y89[20],y89[20],y89[20],y89[20],y89[20],y89[20], y89[20: 0]  }, x213); 

 Register29Bit Reg825 (clk,x213, x213_1 );

 Adder29Bit Adder131(clk,  { x213_1[28: 0] },  {y90[21],y90[21],y90[21],y90[21],y90[21],y90[21],y90[21], y90[21: 0]  }, x214); 

 Register29Bit Reg826 (clk,x214, x214_1 );

 Adder29Bit Adder132(clk,  { x214_1[28: 0] },  {y91[19],y91[19],y91[19],y91[19],y91[19],y91[19],y91[19],y91[19],y91[19], y91[19: 0]  }, x215); 

 Register29Bit Reg827 (clk,x215, x215_1 );

 Adder29Bit Adder133(clk,  { x215_1[28: 0] },  {y92[22],y92[22],y92[22],y92[22],y92[22],y92[22], y92[22: 0]  }, x216); 

 Register29Bit Reg828 (clk,x216, x216_1 );

 Adder29Bit Adder134(clk,  { x216_1[28: 0] },  {y93[19],y93[19],y93[19],y93[19],y93[19],y93[19],y93[19],y93[19],y93[19], y93[19: 0]  }, x217); 

 Register29Bit Reg829 (clk,x217, x217_1 );

 Adder29Bit Adder135(clk,  { x217_1[28: 0] },  {y94[22],y94[22],y94[22],y94[22],y94[22],y94[22], y94[22: 0]  }, x218); 

 Register29Bit Reg830 (clk,x218, x218_1 );

 Adder29Bit Adder136(clk,  { x218_1[28: 0] },  {y95[20],y95[20],y95[20],y95[20],y95[20],y95[20],y95[20],y95[20], y95[20: 0]  }, x219); 

 Register29Bit Reg831 (clk,x219, x219_1 );

 Adder29Bit Adder137(clk,  { x219_1[28: 0] },  {y96[24],y96[24],y96[24],y96[24], y96[24: 0]  }, x220); 

 Register29Bit Reg832 (clk,x220, x220_1 );

 Adder29Bit Adder138(clk,  { x220_1[28: 0] },  {y97[18],y97[18],y97[18],y97[18],y97[18],y97[18],y97[18],y97[18],y97[18],y97[18], y97[18: 0]  }, x221); 

 Register29Bit Reg833 (clk,x221, x221_1 );

 Adder29Bit Adder139(clk,  { x221_1[28: 0] },  {y98[23],y98[23],y98[23],y98[23],y98[23], y98[23: 0]  }, x222); 

 Register29Bit Reg834 (clk,x222, x222_1 );

 Adder29Bit Adder140(clk,  { x222_1[28: 0] },  {y99[15],y99[15],y99[15],y99[15],y99[15],y99[15],y99[15],y99[15],y99[15],y99[15],y99[15],y99[15],y99[15], y99[15: 0]  }, x223); 

 Register29Bit Reg835 (clk,x223, x223_1 );

 Adder29Bit Adder141(clk,  { x223_1[28: 0] },  {y100[24],y100[24],y100[24],y100[24], y100[24: 0]  }, x224); 

 Register29Bit Reg836 (clk,x224, x224_1 );

 Adder29Bit Adder142(clk,  { x224_1[28: 0] },  {y101[19],y101[19],y101[19],y101[19],y101[19],y101[19],y101[19],y101[19],y101[19], y101[19: 0]  }, x225); 

 Register29Bit Reg837 (clk,x225, x225_1 );

 Adder29Bit Adder143(clk,  { x225_1[28: 0] },  {y102[22],y102[22],y102[22],y102[22],y102[22],y102[22], y102[22: 0]  }, x226); 

 Register29Bit Reg838 (clk,x226, x226_1 );

 Adder29Bit Adder144(clk,  { x226_1[28: 0] },  {y103[20],y103[20],y103[20],y103[20],y103[20],y103[20],y103[20],y103[20], y103[20: 0]  }, x227); 

 Register29Bit Reg839 (clk,x227, x227_1 );

 Adder29Bit Adder145(clk,  { x227_1[28: 0] },  {y104[22],y104[22],y104[22],y104[22],y104[22],y104[22], y104[22: 0]  }, x228); 

 Register29Bit Reg840 (clk,x228, x228_1 );

 Adder29Bit Adder146(clk,  { x228_1[28: 0] },  {y105[21],y105[21],y105[21],y105[21],y105[21],y105[21],y105[21], y105[21: 0]  }, x229); 

 Register29Bit Reg841 (clk,x229, x229_1 );

 Adder29Bit Adder147(clk,  { x229_1[28: 0] },  {y106[23],y106[23],y106[23],y106[23],y106[23], y106[23: 0]  }, x230); 

 Register29Bit Reg842 (clk,x230, x230_1 );

 Adder29Bit Adder148(clk,  { x230_1[28: 0] },  {y107[21],y107[21],y107[21],y107[21],y107[21],y107[21],y107[21], y107[21: 0]  }, x231); 

 Register29Bit Reg843 (clk,x231, x231_1 );

 Adder29Bit Adder149(clk,  { x231_1[28: 0] },  {y108[23],y108[23],y108[23],y108[23],y108[23], y108[23: 0]  }, x232); 

 Register29Bit Reg844 (clk,x232, x232_1 );

 Adder29Bit Adder150(clk,  { x232_1[28: 0] },  {y109[22],y109[22],y109[22],y109[22],y109[22],y109[22], y109[22: 0]  }, x233); 

 Register29Bit Reg845 (clk,x233, x233_1 );

 Adder29Bit Adder151(clk,  { x233_1[28: 0] },  {y110[24],y110[24],y110[24],y110[24], y110[24: 0]  }, x234); 

 Register29Bit Reg846 (clk,x234, x234_1 );

 Adder29Bit Adder152(clk,  { x234_1[28: 0] },  {y111[22],y111[22],y111[22],y111[22],y111[22],y111[22], y111[22: 0]  }, x235); 

 Register29Bit Reg847 (clk,x235, x235_1 );

 Adder29Bit Adder153(clk,  { x235_1[28: 0] },  {y112[24],y112[24],y112[24],y112[24], y112[24: 0]  }, x236); 

 Register29Bit Reg848 (clk,x236, x236_1 );

 Adder29Bit Adder154(clk,  { x236_1[28: 0] },  {y113[23],y113[23],y113[23],y113[23],y113[23], y113[23: 0]  }, x237); 

 Register29Bit Reg849 (clk,x237, x237_1 );

 Adder29Bit Adder155(clk,  { x237_1[28: 0] },  {y114[24],y114[24],y114[24],y114[24], y114[24: 0]  }, x238); 

 Register29Bit Reg850 (clk,x238, x238_1 );

 Adder29Bit Adder156(clk,  { x238_1[28: 0] },  {y115[22],y115[22],y115[22],y115[22],y115[22],y115[22], y115[22: 0]  }, x239); 

 Register29Bit Reg851 (clk,x239, x239_1 );

 Adder29Bit Adder157(clk,  { x239_1[28: 0] },  {y116[24],y116[24],y116[24],y116[24], y116[24: 0]  }, x240); 

 Register29Bit Reg852 (clk,x240, x240_1 );

 Adder29Bit Adder158(clk,  { x240_1[28: 0] },  {y117[24],y117[24],y117[24],y117[24], y117[24: 0]  }, x241); 

 Register29Bit Reg853 (clk,x241, x241_1 );

 Adder29Bit Adder159(clk,  { x241_1[28: 0] },  {y118[26],y118[26], y118[26: 0]  }, x242); 

 Register29Bit Reg854 (clk,x242, x242_1 );

 Adder29Bit Adder160(clk,  { x242_1[28: 0] },  {y119[24],y119[24],y119[24],y119[24], y119[24: 0]  }, x243); 

 Register29Bit Reg855 (clk,x243, x243_1 );

 Adder29Bit Adder161(clk,  { x243_1[28: 0] },  {y120[24],y120[24],y120[24],y120[24], y120[24: 0]  }, x244); 

 Register29Bit Reg856 (clk,x244, x244_1 );

 Adder29Bit Adder162(clk,  { x244_1[28: 0] },  {y121[25],y121[25],y121[25], y121[25: 0]  }, x245); 

 Register29Bit Reg857 (clk,x245, x245_1 );

 Adder29Bit Adder163(clk,  { x245_1[28: 0] },  {y122[26],y122[26], y122[26: 0]  }, x246); 

 Register29Bit Reg858 (clk,x246, x246_1 );

 Adder29Bit Adder164(clk,  { x246_1[28: 0] },  {y123[26],y123[26], y123[26: 0]  }, x247); 

 Register29Bit Reg859 (clk,x247, x247_1 );

 Adder29Bit Adder165(clk,  { x247_1[28: 0] },  {y124[26],y124[26], y124[26: 0]  }, x248); 

 Register29Bit Reg860 (clk,x248, x248_1 );

 Adder29Bit Adder166(clk,  { x248_1[28: 0] },  {y125[26],y125[26], y125[26: 0]  }, x249); 

 Register29Bit Reg861 (clk,x249, x249_1 );

 Adder29Bit Adder167(clk,  { x249_1[28: 0] },  {y126[26],y126[26], y126[26: 0]  }, x250); 

 Register29Bit Reg862 (clk,x250, x250_1 );

 Adder29Bit Adder168(clk,  { x250_1[28: 0] },  {y127[26],y127[26], y127[26: 0]  }, x251); 

 Register29Bit Reg863 (clk,x251, x251_1 );

 Adder29Bit Adder169(clk,  { x251_1[28: 0] },  {y128[25],y128[25],y128[25], y128[25: 0]  }, x252); 

 Register29Bit Reg864 (clk,x252, x252_1 );

 Adder29Bit Adder170(clk,  { x252_1[28: 0] },  {y129[24],y129[24],y129[24],y129[24], y129[24: 0]  }, x253); 

 Register29Bit Reg865 (clk,x253, x253_1 );

 Adder29Bit Adder171(clk,  { x253_1[28: 0] },  {y130[24],y130[24],y130[24],y130[24], y130[24: 0]  }, x254); 

 Register29Bit Reg866 (clk,x254, x254_1 );

 Adder29Bit Adder172(clk,  { x254_1[28: 0] },  {y131[26],y131[26], y131[26: 0]  }, x255); 

 Register29Bit Reg867 (clk,x255, x255_1 );

 Adder29Bit Adder173(clk,  { x255_1[28: 0] },  {y132[24],y132[24],y132[24],y132[24], y132[24: 0]  }, x256); 

 Register29Bit Reg868 (clk,x256, x256_1 );

 Adder29Bit Adder174(clk,  { x256_1[28: 0] },  {y133[24],y133[24],y133[24],y133[24], y133[24: 0]  }, x257); 

 Register29Bit Reg869 (clk,x257, x257_1 );

 Adder29Bit Adder175(clk,  { x257_1[28: 0] },  {y134[22],y134[22],y134[22],y134[22],y134[22],y134[22], y134[22: 0]  }, x258); 

 Register29Bit Reg870 (clk,x258, x258_1 );

 Adder29Bit Adder176(clk,  { x258_1[28: 0] },  {y135[24],y135[24],y135[24],y135[24], y135[24: 0]  }, x259); 

 Register29Bit Reg871 (clk,x259, x259_1 );

 Adder29Bit Adder177(clk,  { x259_1[28: 0] },  {y136[23],y136[23],y136[23],y136[23],y136[23], y136[23: 0]  }, x260); 

 Register29Bit Reg872 (clk,x260, x260_1 );

 Adder29Bit Adder178(clk,  { x260_1[28: 0] },  {y137[24],y137[24],y137[24],y137[24], y137[24: 0]  }, x261); 

 Register29Bit Reg873 (clk,x261, x261_1 );

 Adder29Bit Adder179(clk,  { x261_1[28: 0] },  {y138[22],y138[22],y138[22],y138[22],y138[22],y138[22], y138[22: 0]  }, x262); 

 Register29Bit Reg874 (clk,x262, x262_1 );

 Adder29Bit Adder180(clk,  { x262_1[28: 0] },  {y139[24],y139[24],y139[24],y139[24], y139[24: 0]  }, x263); 

 Register29Bit Reg875 (clk,x263, x263_1 );

 Adder29Bit Adder181(clk,  { x263_1[28: 0] },  {y140[22],y140[22],y140[22],y140[22],y140[22],y140[22], y140[22: 0]  }, x264); 

 Register29Bit Reg876 (clk,x264, x264_1 );

 Adder29Bit Adder182(clk,  { x264_1[28: 0] },  {y141[23],y141[23],y141[23],y141[23],y141[23], y141[23: 0]  }, x265); 

 Register29Bit Reg877 (clk,x265, x265_1 );

 Adder29Bit Adder183(clk,  { x265_1[28: 0] },  {y142[21],y142[21],y142[21],y142[21],y142[21],y142[21],y142[21], y142[21: 0]  }, x266); 

 Register29Bit Reg878 (clk,x266, x266_1 );

 Adder29Bit Adder184(clk,  { x266_1[28: 0] },  {y143[23],y143[23],y143[23],y143[23],y143[23], y143[23: 0]  }, x267); 

 Register29Bit Reg879 (clk,x267, x267_1 );

 Adder29Bit Adder185(clk,  { x267_1[28: 0] },  {y144[21],y144[21],y144[21],y144[21],y144[21],y144[21],y144[21], y144[21: 0]  }, x268); 

 Register29Bit Reg880 (clk,x268, x268_1 );

 Adder29Bit Adder186(clk,  { x268_1[28: 0] },  {y145[22],y145[22],y145[22],y145[22],y145[22],y145[22], y145[22: 0]  }, x269); 

 Register29Bit Reg881 (clk,x269, x269_1 );

 Adder29Bit Adder187(clk,  { x269_1[28: 0] },  {y146[20],y146[20],y146[20],y146[20],y146[20],y146[20],y146[20],y146[20], y146[20: 0]  }, x270); 

 Register29Bit Reg882 (clk,x270, x270_1 );

 Adder29Bit Adder188(clk,  { x270_1[28: 0] },  {y147[22],y147[22],y147[22],y147[22],y147[22],y147[22], y147[22: 0]  }, x271); 

 Register29Bit Reg883 (clk,x271, x271_1 );

 Adder29Bit Adder189(clk,  { x271_1[28: 0] },  {y148[19],y148[19],y148[19],y148[19],y148[19],y148[19],y148[19],y148[19],y148[19], y148[19: 0]  }, x272); 

 Register29Bit Reg884 (clk,x272, x272_1 );

 Adder29Bit Adder190(clk,  { x272_1[28: 0] },  {y149[24],y149[24],y149[24],y149[24], y149[24: 0]  }, x273); 

 Register29Bit Reg885 (clk,x273, x273_1 );

 Adder29Bit Adder191(clk,  { x273_1[28: 0] },  {y150[15],y150[15],y150[15],y150[15],y150[15],y150[15],y150[15],y150[15],y150[15],y150[15],y150[15],y150[15],y150[15], y150[15: 0]  }, x274); 

 Register29Bit Reg886 (clk,x274, x274_1 );

 Adder29Bit Adder192(clk,  { x274_1[28: 0] },  {y151[23],y151[23],y151[23],y151[23],y151[23], y151[23: 0]  }, x275); 

 Register29Bit Reg887 (clk,x275, x275_1 );

 Adder29Bit Adder193(clk,  { x275_1[28: 0] },  {y152[18],y152[18],y152[18],y152[18],y152[18],y152[18],y152[18],y152[18],y152[18],y152[18], y152[18: 0]  }, x276); 

 Register29Bit Reg888 (clk,x276, x276_1 );

 Adder29Bit Adder194(clk,  { x276_1[28: 0] },  {y153[24],y153[24],y153[24],y153[24], y153[24: 0]  }, x277); 

 Register29Bit Reg889 (clk,x277, x277_1 );

 Adder29Bit Adder195(clk,  { x277_1[28: 0] },  {y154[20],y154[20],y154[20],y154[20],y154[20],y154[20],y154[20],y154[20], y154[20: 0]  }, x278); 

 Register29Bit Reg890 (clk,x278, x278_1 );

 Adder29Bit Adder196(clk,  { x278_1[28: 0] },  {y155[22],y155[22],y155[22],y155[22],y155[22],y155[22], y155[22: 0]  }, x279); 

 Register29Bit Reg891 (clk,x279, x279_1 );

 Adder29Bit Adder197(clk,  { x279_1[28: 0] },  {y156[19],y156[19],y156[19],y156[19],y156[19],y156[19],y156[19],y156[19],y156[19], y156[19: 0]  }, x280); 

 Register29Bit Reg892 (clk,x280, x280_1 );

 Adder29Bit Adder198(clk,  { x280_1[28: 0] },  {y157[22],y157[22],y157[22],y157[22],y157[22],y157[22], y157[22: 0]  }, x281); 

 Register29Bit Reg893 (clk,x281, x281_1 );

 Adder29Bit Adder199(clk,  { x281_1[28: 0] },  {y158[19],y158[19],y158[19],y158[19],y158[19],y158[19],y158[19],y158[19],y158[19], y158[19: 0]  }, x282); 

 Register29Bit Reg894 (clk,x282, x282_1 );

 Adder29Bit Adder200(clk,  { x282_1[28: 0] },  {y159[21],y159[21],y159[21],y159[21],y159[21],y159[21],y159[21], y159[21: 0]  }, x283); 

 Register29Bit Reg895 (clk,x283, x283_1 );

 Adder29Bit Adder201(clk,  { x283_1[28: 0] },  {y160[20],y160[20],y160[20],y160[20],y160[20],y160[20],y160[20],y160[20], y160[20: 0]  }, x284); 

 Register29Bit Reg896 (clk,x284, x284_1 );

 Adder29Bit Adder202(clk,  { x284_1[28: 0] },  {y161[22],y161[22],y161[22],y161[22],y161[22],y161[22], y161[22: 0]  }, x285); 

 Register29Bit Reg897 (clk,x285, x285_1 );

 Adder29Bit Adder203(clk,  { x285_1[28: 0] },  {y162[21],y162[21],y162[21],y162[21],y162[21],y162[21],y162[21], y162[21: 0]  }, x286); 

 Register29Bit Reg898 (clk,x286, x286_1 );

 Adder29Bit Adder204(clk,  { x286_1[28: 0] },  {y163[22],y163[22],y163[22],y163[22],y163[22],y163[22], y163[22: 0]  }, x287); 

 Register29Bit Reg899 (clk,x287, x287_1 );

 Adder29Bit Adder205(clk,  { x287_1[28: 0] },  {y164[21],y164[21],y164[21],y164[21],y164[21],y164[21],y164[21], y164[21: 0]  }, x288); 

 Register29Bit Reg900 (clk,x288, x288_1 );

 Adder29Bit Adder206(clk,  { x288_1[28: 0] },  {y165[22],y165[22],y165[22],y165[22],y165[22],y165[22], y165[22: 0]  }, x289); 

 Register29Bit Reg901 (clk,x289, x289_1 );

 Adder29Bit Adder207(clk,  { x289_1[28: 0] },  {y166[21],y166[21],y166[21],y166[21],y166[21],y166[21],y166[21], y166[21: 0]  }, x290); 

 Register29Bit Reg902 (clk,x290, x290_1 );

 Adder29Bit Adder208(clk,  { x290_1[28: 0] },  {y167[22],y167[22],y167[22],y167[22],y167[22],y167[22], y167[22: 0]  }, x291); 

 Register29Bit Reg903 (clk,x291, x291_1 );

 Adder29Bit Adder209(clk,  { x291_1[28: 0] },  {y168[21],y168[21],y168[21],y168[21],y168[21],y168[21],y168[21], y168[21: 0]  }, x292); 

 Register29Bit Reg904 (clk,x292, x292_1 );

 Adder29Bit Adder210(clk,  { x292_1[28: 0] },  {y169[21],y169[21],y169[21],y169[21],y169[21],y169[21],y169[21], y169[21: 0]  }, x293); 

 Register29Bit Reg905 (clk,x293, x293_1 );

 Adder29Bit Adder211(clk,  { x293_1[28: 0] },  {y170[21],y170[21],y170[21],y170[21],y170[21],y170[21],y170[21], y170[21: 0]  }, x294); 

 Register29Bit Reg906 (clk,x294, x294_1 );

 Adder29Bit Adder212(clk,  { x294_1[28: 0] },  {y171[21],y171[21],y171[21],y171[21],y171[21],y171[21],y171[21], y171[21: 0]  }, x295); 

 Register29Bit Reg907 (clk,x295, x295_1 );

 Adder29Bit Adder213(clk,  { x295_1[28: 0] },  {y172[21],y172[21],y172[21],y172[21],y172[21],y172[21],y172[21], y172[21: 0]  }, x296); 

 Register29Bit Reg908 (clk,x296, x296_1 );

 Adder29Bit Adder214(clk,  { x296_1[28: 0] },  {y173[20],y173[20],y173[20],y173[20],y173[20],y173[20],y173[20],y173[20], y173[20: 0]  }, x297); 

 Register29Bit Reg909 (clk,x297, x297_1 );

 Adder29Bit Adder215(clk,  { x297_1[28: 0] },  {y174[21],y174[21],y174[21],y174[21],y174[21],y174[21],y174[21], y174[21: 0]  }, x298); 

 Register29Bit Reg910 (clk,x298, x298_1 );

 Adder29Bit Adder216(clk,  { x298_1[28: 0] },  {y175[21],y175[21],y175[21],y175[21],y175[21],y175[21],y175[21], y175[21: 0]  }, x299); 

 Register29Bit Reg911 (clk,x299, x299_1 );

 Adder29Bit Adder217(clk,  { x299_1[28: 0] },  {y176[20],y176[20],y176[20],y176[20],y176[20],y176[20],y176[20],y176[20], y176[20: 0]  }, x300); 

 Register29Bit Reg912 (clk,x300, x300_1 );

 Adder29Bit Adder218(clk,  { x300_1[28: 0] },  {y177[20],y177[20],y177[20],y177[20],y177[20],y177[20],y177[20],y177[20], y177[20: 0]  }, x301); 

 Register29Bit Reg913 (clk,x301, x301_1 );

 Adder29Bit Adder219(clk,  { x301_1[28: 0] },  {y178[21],y178[21],y178[21],y178[21],y178[21],y178[21],y178[21], y178[21: 0]  }, x302); 

 Register29Bit Reg914 (clk,x302, x302_1 );

 Adder29Bit Adder220(clk,  { x302_1[28: 0] },  {y179[20],y179[20],y179[20],y179[20],y179[20],y179[20],y179[20],y179[20], y179[20: 0]  }, x303); 

 Register29Bit Reg915 (clk,x303, x303_1 );

 Adder29Bit Adder221(clk,  { x303_1[28: 0] },  {y180[21],y180[21],y180[21],y180[21],y180[21],y180[21],y180[21], y180[21: 0]  }, x304); 

 Register29Bit Reg916 (clk,x304, x304_1 );

 Adder29Bit Adder222(clk,  { x304_1[28: 0] },  {y181[19],y181[19],y181[19],y181[19],y181[19],y181[19],y181[19],y181[19],y181[19], y181[19: 0]  }, x305); 

 Register29Bit Reg917 (clk,x305, x305_1 );

 Adder29Bit Adder223(clk,  { x305_1[28: 0] },  {y182[21],y182[21],y182[21],y182[21],y182[21],y182[21],y182[21], y182[21: 0]  }, x306); 

 Register29Bit Reg918 (clk,x306, x306_1 );

 Adder29Bit Adder224(clk,  { x306_1[28: 0] },  {y183[19],y183[19],y183[19],y183[19],y183[19],y183[19],y183[19],y183[19],y183[19], y183[19: 0]  }, x307); 

 Register29Bit Reg919 (clk,x307, x307_1 );

 Adder29Bit Adder225(clk,  { x307_1[28: 0] },  {y184[21],y184[21],y184[21],y184[21],y184[21],y184[21],y184[21], y184[21: 0]  }, x308); 

 Register29Bit Reg920 (clk,x308, x308_1 );

 Adder29Bit Adder226(clk,  { x308_1[28: 0] },  {y185[20],y185[20],y185[20],y185[20],y185[20],y185[20],y185[20],y185[20], y185[20: 0]  }, x309); 

 Register29Bit Reg921 (clk,x309, x309_1 );

 Adder29Bit Adder227(clk,  { x309_1[28: 0] },  {y186[21],y186[21],y186[21],y186[21],y186[21],y186[21],y186[21], y186[21: 0]  }, x310); 

 Register29Bit Reg922 (clk,x310, x310_1 );

 Adder29Bit Adder228(clk,  { x310_1[28: 0] },  {y187[20],y187[20],y187[20],y187[20],y187[20],y187[20],y187[20],y187[20], y187[20: 0]  }, x311); 

 Register29Bit Reg923 (clk,x311, x311_1 );

 Adder29Bit Adder229(clk,  { x311_1[28: 0] },  {y188[21],y188[21],y188[21],y188[21],y188[21],y188[21],y188[21], y188[21: 0]  }, x312); 

 Register29Bit Reg924 (clk,x312, x312_1 );

 Adder29Bit Adder230(clk,  { x312_1[28: 0] },  {y189[18],y189[18],y189[18],y189[18],y189[18],y189[18],y189[18],y189[18],y189[18],y189[18], y189[18: 0]  }, x313); 

 Register29Bit Reg925 (clk,x313, x313_1 );

 Adder29Bit Adder231(clk,  { x313_1[28: 0] },  {y190[20],y190[20],y190[20],y190[20],y190[20],y190[20],y190[20],y190[20], y190[20: 0]  }, x314); 

 Register29Bit Reg926 (clk,x314, x314_1 );

 Adder29Bit Adder232(clk,  { x314_1[28: 0] },  {y191[19],y191[19],y191[19],y191[19],y191[19],y191[19],y191[19],y191[19],y191[19], y191[19: 0]  }, x315); 

 Register29Bit Reg927 (clk,x315, x315_1 );

 Adder29Bit Adder233(clk,  { x315_1[28: 0] },  {y192[19],y192[19],y192[19],y192[19],y192[19],y192[19],y192[19],y192[19],y192[19], y192[19: 0]  }, x316); 

 Register29Bit Reg928 (clk,x316, x316_1 );

 Adder29Bit Adder234(clk,  { x316_1[28: 0] },  {y193[19],y193[19],y193[19],y193[19],y193[19],y193[19],y193[19],y193[19],y193[19], y193[19: 0]  }, x317); 

 Register29Bit Reg929 (clk,x317, x317_1 );

 Adder29Bit Adder235(clk,  { x317_1[28: 0] },  {y194[20],y194[20],y194[20],y194[20],y194[20],y194[20],y194[20],y194[20], y194[20: 0]  }, x318); 

 Register29Bit Reg930 (clk,x318, x318_1 );

 Adder29Bit Adder236(clk,  { x318_1[28: 0] },  {y195[17],y195[17],y195[17],y195[17],y195[17],y195[17],y195[17],y195[17],y195[17],y195[17],y195[17], y195[17: 0]  }, x319); 

 Register29Bit Reg931 (clk,x319, x319_1 );

 Adder29Bit Adder237(clk,  { x319_1[28: 0] },  {y196[20],y196[20],y196[20],y196[20],y196[20],y196[20],y196[20],y196[20], y196[20: 0]  }, x320); 

 Register29Bit Reg932 (clk,x320, x320_1 );

 Adder29Bit Adder238(clk,  { x320_1[28: 0] },  {y197[18],y197[18],y197[18],y197[18],y197[18],y197[18],y197[18],y197[18],y197[18],y197[18], y197[18: 0]  }, x321); 

 Register29Bit Reg933 (clk,x321, x321_1 );

 Adder29Bit Adder239(clk,  { x321_1[28: 0] },  {y198[19],y198[19],y198[19],y198[19],y198[19],y198[19],y198[19],y198[19],y198[19], y198[19: 0]  }, x322); 

 Register29Bit Reg934 (clk,x322, x322_1 );

 Adder29Bit Adder240(clk,  { x322_1[28: 0] },  {y199[16],y199[16],y199[16],y199[16],y199[16],y199[16],y199[16],y199[16],y199[16],y199[16],y199[16],y199[16], y199[16: 0]  }, x323); 

 Register29Bit Reg935 (clk,x323, x323_1 );

 Adder29Bit Adder241(clk,  { x323_1[28: 0] },  {y200[19],y200[19],y200[19],y200[19],y200[19],y200[19],y200[19],y200[19],y200[19], y200[19: 0]  }, x324); 

 Register29Bit Reg936 (clk,x324, x324_1 );

 Adder29Bit Adder242(clk,  { x324_1[28: 0] },  {y201[15],y201[15],y201[15],y201[15],y201[15],y201[15],y201[15],y201[15],y201[15],y201[15],y201[15],y201[15],y201[15], y201[15: 0]  }, x325); 

 Register29Bit Reg937 (clk,x325, x325_1 );

 Adder29Bit Adder243(clk,  { x325_1[28: 0] },  {y202[20],y202[20],y202[20],y202[20],y202[20],y202[20],y202[20],y202[20], y202[20: 0]  }, x326); 

 Register29Bit Reg938 (clk,x326, x326_1 );

 Adder29Bit Adder244(clk,  { x326_1[28: 0] },  {y203[11],y203[11],y203[11],y203[11],y203[11],y203[11],y203[11],y203[11],y203[11],y203[11],y203[11],y203[11],y203[11],y203[11],y203[11],y203[11],y203[11], y203[11: 0]  }, x327); 

 Register29Bit Reg939 (clk,x327, x327_1 );

 Adder29Bit Adder245(clk,  { x327_1[28: 0] },  {y204[20],y204[20],y204[20],y204[20],y204[20],y204[20],y204[20],y204[20], y204[20: 0]  }, x328); 

 Register29Bit Reg940 (clk,x328, x328_1 );

 Adder29Bit Adder246(clk,  { x328_1[28: 0] },  {y205[15],y205[15],y205[15],y205[15],y205[15],y205[15],y205[15],y205[15],y205[15],y205[15],y205[15],y205[15],y205[15], y205[15: 0]  }, x329); 

 Register29Bit Reg941 (clk,x329, x329_1 );

 Adder29Bit Adder247(clk,  { x329_1[28: 0] },  {y206[20],y206[20],y206[20],y206[20],y206[20],y206[20],y206[20],y206[20], y206[20: 0]  }, x330); 

 Register29Bit Reg942 (clk,x330, x330_1 );

 Adder29Bit Adder248(clk,  { x330_1[28: 0] },  {y207[15],y207[15],y207[15],y207[15],y207[15],y207[15],y207[15],y207[15],y207[15],y207[15],y207[15],y207[15],y207[15], y207[15: 0]  }, x331); 

 Register29Bit Reg943 (clk,x331, x331_1 );

 Adder29Bit Adder249(clk,  { x331_1[28: 0] },  {y208[20],y208[20],y208[20],y208[20],y208[20],y208[20],y208[20],y208[20], y208[20: 0]  }, x332); 

 Register29Bit Reg944 (clk,x332, x332_1 );

 Adder29Bit Adder250(clk,  { x332_1[28: 0] },  {y209[16],y209[16],y209[16],y209[16],y209[16],y209[16],y209[16],y209[16],y209[16],y209[16],y209[16],y209[16], y209[16: 0]  }, x333); 

 Register29Bit Reg945 (clk,x333, x333_1 );

 Adder29Bit Adder251(clk,  { x333_1[28: 0] },  {y210[19],y210[19],y210[19],y210[19],y210[19],y210[19],y210[19],y210[19],y210[19], y210[19: 0]  }, x334); 

 Register29Bit Reg946 (clk,x334, x334_1 );

 Adder29Bit Adder252(clk,  { x334_1[28: 0] },  {y211[16],y211[16],y211[16],y211[16],y211[16],y211[16],y211[16],y211[16],y211[16],y211[16],y211[16],y211[16], y211[16: 0]  }, x335); 

 Register29Bit Reg947 (clk,x335, x335_1 );

 Adder29Bit Adder253(clk,  { x335_1[28: 0] },  {y212[19],y212[19],y212[19],y212[19],y212[19],y212[19],y212[19],y212[19],y212[19], y212[19: 0]  }, x336); 

 Register29Bit Reg948 (clk,x336, x336_1 );

 Adder29Bit Adder254(clk,  { x336_1[28: 0] },  {y213[16],y213[16],y213[16],y213[16],y213[16],y213[16],y213[16],y213[16],y213[16],y213[16],y213[16],y213[16], y213[16: 0]  }, x337); 

 Register29Bit Reg949 (clk,x337, x337_1 );

 Adder29Bit Adder255(clk,  { x337_1[28: 0] },  {y214[18],y214[18],y214[18],y214[18],y214[18],y214[18],y214[18],y214[18],y214[18],y214[18], y214[18: 0]  }, x338); 

 Register29Bit Reg950 (clk,x338, x338_1 );

 Adder29Bit Adder256(clk,  { x338_1[28: 0] },  {y215[16],y215[16],y215[16],y215[16],y215[16],y215[16],y215[16],y215[16],y215[16],y215[16],y215[16],y215[16], y215[16: 0]  }, x339); 

 Register29Bit Reg951 (clk,x339, x339_1 );

 Adder29Bit Adder257(clk,  { x339_1[28: 0] },  {y216[18],y216[18],y216[18],y216[18],y216[18],y216[18],y216[18],y216[18],y216[18],y216[18], y216[18: 0]  }, x340); 

 Register29Bit Reg952 (clk,x340, x340_1 );

 Adder29Bit Adder258(clk,  { x340_1[28: 0] },  {y217[16],y217[16],y217[16],y217[16],y217[16],y217[16],y217[16],y217[16],y217[16],y217[16],y217[16],y217[16], y217[16: 0]  }, x341); 

 Register29Bit Reg953 (clk,x341, x341_1 );

 Adder29Bit Adder259(clk,  { x341_1[28: 0] },  {y218[18],y218[18],y218[18],y218[18],y218[18],y218[18],y218[18],y218[18],y218[18],y218[18], y218[18: 0]  }, x342); 

 Register29Bit Reg954 (clk,x342, x342_1 );

 Adder29Bit Adder260(clk,  { x342_1[28: 0] },  {y219[16],y219[16],y219[16],y219[16],y219[16],y219[16],y219[16],y219[16],y219[16],y219[16],y219[16],y219[16], y219[16: 0]  }, x343); 

 Register29Bit Reg955 (clk,x343, x343_1 );

 Adder29Bit Adder261(clk,  { x343_1[28: 0] },  {y220[19],y220[19],y220[19],y220[19],y220[19],y220[19],y220[19],y220[19],y220[19], y220[19: 0]  }, x344); 

 Register29Bit Reg956 (clk,x344, x344_1 );

 Adder29Bit Adder262(clk,  { x344_1[28: 0] },  {y221[17],y221[17],y221[17],y221[17],y221[17],y221[17],y221[17],y221[17],y221[17],y221[17],y221[17], y221[17: 0]  }, x345); 

 Register29Bit Reg957 (clk,x345, x345_1 );

 Adder29Bit Adder263(clk,  { x345_1[28: 0] },  {y222[19],y222[19],y222[19],y222[19],y222[19],y222[19],y222[19],y222[19],y222[19], y222[19: 0]  }, x346); 

 Register29Bit Reg958 (clk,x346, x346_1 );

 Adder29Bit Adder264(clk,  { x346_1[28: 0] },  {y223[16],y223[16],y223[16],y223[16],y223[16],y223[16],y223[16],y223[16],y223[16],y223[16],y223[16],y223[16], y223[16: 0]  }, x347); 

 Register29Bit Reg959 (clk,x347, x347_1 );

 Adder29Bit Adder265(clk,  { x347_1[28: 0] },  {y224[17],y224[17],y224[17],y224[17],y224[17],y224[17],y224[17],y224[17],y224[17],y224[17],y224[17], y224[17: 0]  }, x348); 

 Register29Bit Reg960 (clk,x348, x348_1 );

 Adder29Bit Adder266(clk,  { x348_1[28: 0] },  {y225[16],y225[16],y225[16],y225[16],y225[16],y225[16],y225[16],y225[16],y225[16],y225[16],y225[16],y225[16], y225[16: 0]  }, x349); 

 Register29Bit Reg961 (clk,x349, x349_1 );

 Adder29Bit Adder267(clk,  { x349_1[28: 0] },  {y226[17],y226[17],y226[17],y226[17],y226[17],y226[17],y226[17],y226[17],y226[17],y226[17],y226[17], y226[17: 0]  }, x350); 

 Register29Bit Reg962 (clk,x350, x350_1 );

 Adder29Bit Adder268(clk,  { x350_1[28: 0] },  {y227[16],y227[16],y227[16],y227[16],y227[16],y227[16],y227[16],y227[16],y227[16],y227[16],y227[16],y227[16], y227[16: 0]  }, x351); 

 Register29Bit Reg963 (clk,x351, x351_1 );

 Adder29Bit Adder269(clk,  { x351_1[28: 0] },  {y228[17],y228[17],y228[17],y228[17],y228[17],y228[17],y228[17],y228[17],y228[17],y228[17],y228[17], y228[17: 0]  }, x352); 

 Register29Bit Reg964 (clk,x352, x352_1 );

 Adder29Bit Adder270(clk,  { x352_1[28: 0] },  {y229[16],y229[16],y229[16],y229[16],y229[16],y229[16],y229[16],y229[16],y229[16],y229[16],y229[16],y229[16], y229[16: 0]  }, x353); 

 Register29Bit Reg965 (clk,x353, x353_1 );

 Adder29Bit Adder271(clk,  { x353_1[28: 0] },  {y230[17],y230[17],y230[17],y230[17],y230[17],y230[17],y230[17],y230[17],y230[17],y230[17],y230[17], y230[17: 0]  }, x354); 

 Register29Bit Reg966 (clk,x354, x354_1 );

 Adder29Bit Adder272(clk,  { x354_1[28: 0] },  {y231[16],y231[16],y231[16],y231[16],y231[16],y231[16],y231[16],y231[16],y231[16],y231[16],y231[16],y231[16], y231[16: 0]  }, x355); 

 Register29Bit Reg967 (clk,x355, x355_1 );

 Adder29Bit Adder273(clk,  { x355_1[28: 0] },  {y232[18],y232[18],y232[18],y232[18],y232[18],y232[18],y232[18],y232[18],y232[18],y232[18], y232[18: 0]  }, x356); 

 Register29Bit Reg968 (clk,x356, x356_1 );

 Adder29Bit Adder274(clk,  { x356_1[28: 0] },  {y233[16],y233[16],y233[16],y233[16],y233[16],y233[16],y233[16],y233[16],y233[16],y233[16],y233[16],y233[16], y233[16: 0]  }, x357); 

 Register29Bit Reg969 (clk,x357, x357_1 );

 Adder29Bit Adder275(clk,  { x357_1[28: 0] },  {y234[17],y234[17],y234[17],y234[17],y234[17],y234[17],y234[17],y234[17],y234[17],y234[17],y234[17], y234[17: 0]  }, x358); 

 Register29Bit Reg970 (clk,x358, x358_1 );

 Adder29Bit Adder276(clk,  { x358_1[28: 0] },  {y235[16],y235[16],y235[16],y235[16],y235[16],y235[16],y235[16],y235[16],y235[16],y235[16],y235[16],y235[16], y235[16: 0]  }, x359); 

 Register29Bit Reg971 (clk,x359, x359_1 );

 Adder29Bit Adder277(clk,  { x359_1[28: 0] },  {y236[16],y236[16],y236[16],y236[16],y236[16],y236[16],y236[16],y236[16],y236[16],y236[16],y236[16],y236[16], y236[16: 0]  }, x360); 

 Register29Bit Reg972 (clk,x360, x360_1 );

 Adder29Bit Adder278(clk,  { x360_1[28: 0] },  {y237[16],y237[16],y237[16],y237[16],y237[16],y237[16],y237[16],y237[16],y237[16],y237[16],y237[16],y237[16], y237[16: 0]  }, x361); 

 Register29Bit Reg973 (clk,x361, x361_1 );

 Adder29Bit Adder279(clk,  { x361_1[28: 0] },  {y238[16],y238[16],y238[16],y238[16],y238[16],y238[16],y238[16],y238[16],y238[16],y238[16],y238[16],y238[16], y238[16: 0]  }, x362); 

 Register29Bit Reg974 (clk,x362, x362_1 );

 Adder29Bit Adder280(clk,  { x362_1[28: 0] },  {y239[15],y239[15],y239[15],y239[15],y239[15],y239[15],y239[15],y239[15],y239[15],y239[15],y239[15],y239[15],y239[15], y239[15: 0]  }, x363); 

 Register29Bit Reg975 (clk,x363, x363_1 );

 Adder29Bit Adder281(clk,  { x363_1[28: 0] },  {y240[16],y240[16],y240[16],y240[16],y240[16],y240[16],y240[16],y240[16],y240[16],y240[16],y240[16],y240[16], y240[16: 0]  }, x364); 

 Register29Bit Reg976 (clk,x364, x364_1 );

 Adder29Bit Adder282(clk,  { x364_1[28: 0] },  {y241[14],y241[14],y241[14],y241[14],y241[14],y241[14],y241[14],y241[14],y241[14],y241[14],y241[14],y241[14],y241[14],y241[14], y241[14: 0]  }, x365); 

 Register29Bit Reg977 (clk,x365, x365_1 );

 Adder29Bit Adder283(clk,  { x365_1[28: 0] },  {y242[16],y242[16],y242[16],y242[16],y242[16],y242[16],y242[16],y242[16],y242[16],y242[16],y242[16],y242[16], y242[16: 0]  }, x366); 

 Register29Bit Reg978 (clk,x366, x366_1 );

 Adder29Bit Adder284(clk,  { x366_1[28: 0] },  {y243[14],y243[14],y243[14],y243[14],y243[14],y243[14],y243[14],y243[14],y243[14],y243[14],y243[14],y243[14],y243[14],y243[14], y243[14: 0]  }, x367); 

 Register29Bit Reg979 (clk,x367, x367_1 );

 Adder29Bit Adder285(clk,  { x367_1[28: 0] },  {y244[16],y244[16],y244[16],y244[16],y244[16],y244[16],y244[16],y244[16],y244[16],y244[16],y244[16],y244[16], y244[16: 0]  }, x368); 

 Register29Bit Reg980 (clk,x368, x368_1 );

 Adder29Bit Adder286(clk,  { x368_1[28: 0] },  {y245[14],y245[14],y245[14],y245[14],y245[14],y245[14],y245[14],y245[14],y245[14],y245[14],y245[14],y245[14],y245[14],y245[14], y245[14: 0]  }, x369); 

 Register29Bit Reg981 (clk,x369, x369_1 );

 Adder29Bit Adder287(clk,  { x369_1[28: 0] },  {y246[17],y246[17],y246[17],y246[17],y246[17],y246[17],y246[17],y246[17],y246[17],y246[17],y246[17], y246[17: 0]  }, x370); 

 Register29Bit Reg982 (clk,x370, x370_1 );

 Adder29Bit Adder288(clk,  { x370_1[28: 0] },  {y247[12],y247[12],y247[12],y247[12],y247[12],y247[12],y247[12],y247[12],y247[12],y247[12],y247[12],y247[12],y247[12],y247[12],y247[12],y247[12], y247[12: 0]  }, x371); 

 Register29Bit Reg983 (clk,x371, x371_1 );

 Adder29Bit Adder289(clk,  { x371_1[28: 0] },  {y248[15],y248[15],y248[15],y248[15],y248[15],y248[15],y248[15],y248[15],y248[15],y248[15],y248[15],y248[15],y248[15], y248[15: 0]  }, x372); 

 Register29Bit Reg984 (clk,x372, x372_1 );

 Adder29Bit Adder290(clk,  { x372_1[28: 0] },  {y249[14],y249[14],y249[14],y249[14],y249[14],y249[14],y249[14],y249[14],y249[14],y249[14],y249[14],y249[14],y249[14],y249[14], y249[14: 0]  }, Out_Y_wire); 

 endmodule 



module Adder17Bit (clk, In1, In2, AddOut);
 input clk;
 input [16:0] In1, In2; 

 output [17:0] AddOut;

 reg [17 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder24Bit (clk, In1, In2, AddOut);
 input clk;
 input [23:0] In1, In2; 

 output [24:0] AddOut;

 reg [24 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder22Bit (clk, In1, In2, AddOut);
 input clk;
 input [21:0] In1, In2; 

 output [22:0] AddOut;

 reg [22 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder25Bit (clk, In1, In2, AddOut);
 input clk;
 input [24:0] In1, In2; 

 output [25:0] AddOut;

 reg [25 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder19Bit (clk, In1, In2, AddOut);
 input clk;
 input [18:0] In1, In2; 

 output [19:0] AddOut;

 reg [19 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder18Bit (clk, In1, In2, AddOut);
 input clk;
 input [17:0] In1, In2; 

 output [18:0] AddOut;

 reg [18 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder20Bit (clk, In1, In2, AddOut);
 input clk;
 input [19:0] In1, In2; 

 output [20:0] AddOut;

 reg [20 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder23Bit (clk, In1, In2, AddOut);
 input clk;
 input [22:0] In1, In2; 

 output [23:0] AddOut;

 reg [23 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder21Bit (clk, In1, In2, AddOut);
 input clk;
 input [20:0] In1, In2; 

 output [21:0] AddOut;

 reg [21 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder14Bit (clk, In1, In2, AddOut);
 input clk;
 input [13:0] In1, In2; 

 output [14:0] AddOut;

 reg [14 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder15Bit (clk, In1, In2, AddOut);
 input clk;
 input [14:0] In1, In2; 

 output [15:0] AddOut;

 reg [15 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder16Bit (clk, In1, In2, AddOut);
 input clk;
 input [15:0] In1, In2; 

 output [16:0] AddOut;

 reg [16 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder26Bit (clk, In1, In2, AddOut);
 input clk;
 input [25:0] In1, In2; 

 output [26:0] AddOut;

 reg [26 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder27Bit (clk, In1, In2, AddOut);
 input clk;
 input [26:0] In1, In2; 

 output [27:0] AddOut;

 reg [27 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder28Bit (clk, In1, In2, AddOut);
 input clk;
 input [27:0] In1, In2; 

 output [28:0] AddOut;

 reg [28 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule

module Adder29Bit (clk, In1, In2, AddOut);
 input clk;
 input [28:0] In1, In2; 

 output [28:0] AddOut;

 reg [28 :0] AddOut; 

always @(posedge clk)
begin
AddOut <= (In1 + In2);
end
endmodule



module Subtractor14Bit (clk, In1, In2, SubOut);
 input clk;
 input [13:0] In1, In2;
 output [14 :0] SubOut;

 reg [14 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule

module Subtractor21Bit (clk, In1, In2, SubOut);
 input clk;
 input [20:0] In1, In2;
 output [21 :0] SubOut;

 reg [21 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule

module Subtractor19Bit (clk, In1, In2, SubOut);
 input clk;
 input [18:0] In1, In2;
 output [19 :0] SubOut;

 reg [19 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule

module Subtractor24Bit (clk, In1, In2, SubOut);
 input clk;
 input [23:0] In1, In2;
 output [24 :0] SubOut;

 reg [24 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule

module Subtractor20Bit (clk, In1, In2, SubOut);
 input clk;
 input [19:0] In1, In2;
 output [20 :0] SubOut;

 reg [20 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule

module Subtractor22Bit (clk, In1, In2, SubOut);
 input clk;
 input [21:0] In1, In2;
 output [22 :0] SubOut;

 reg [22 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule

module Subtractor16Bit (clk, In1, In2, SubOut);
 input clk;
 input [15:0] In1, In2;
 output [16 :0] SubOut;

 reg [16 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule

module Subtractor18Bit (clk, In1, In2, SubOut);
 input clk;
 input [17:0] In1, In2;
 output [18 :0] SubOut;

 reg [18 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule

module Subtractor17Bit (clk, In1, In2, SubOut);
 input clk;
 input [16:0] In1, In2;
 output [17 :0] SubOut;

 reg [17 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule

module Subtractor23Bit (clk, In1, In2, SubOut);
 input clk;
 input [22:0] In1, In2;
 output [23 :0] SubOut;

 reg [23 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule

module Subtractor15Bit (clk, In1, In2, SubOut);
 input clk;
 input [14:0] In1, In2;
 output [15 :0] SubOut;

 reg [15 :0] SubOut; 

always @(posedge clk)
begin
SubOut <= (In1 - In2);
end
endmodule



module Register25Bit (clk, In1, RegOut);
 input clk;
 input [24:0] In1;
 output [24 :0] RegOut;

 reg [24 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register23Bit (clk, In1, RegOut);
 input clk;
 input [22:0] In1;
 output [22 :0] RegOut;

 reg [22 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register26Bit (clk, In1, RegOut);
 input clk;
 input [25:0] In1;
 output [25 :0] RegOut;

 reg [25 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register27Bit (clk, In1, RegOut);
 input clk;
 input [26:0] In1;
 output [26 :0] RegOut;

 reg [26 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register18Bit (clk, In1, RegOut);
 input clk;
 input [17:0] In1;
 output [17 :0] RegOut;

 reg [17 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register21Bit (clk, In1, RegOut);
 input clk;
 input [20:0] In1;
 output [20 :0] RegOut;

 reg [20 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register19Bit (clk, In1, RegOut);
 input clk;
 input [18:0] In1;
 output [18 :0] RegOut;

 reg [18 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register22Bit (clk, In1, RegOut);
 input clk;
 input [21:0] In1;
 output [21 :0] RegOut;

 reg [21 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register20Bit (clk, In1, RegOut);
 input clk;
 input [19:0] In1;
 output [19 :0] RegOut;

 reg [19 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register17Bit (clk, In1, RegOut);
 input clk;
 input [16:0] In1;
 output [16 :0] RegOut;

 reg [16 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register24Bit (clk, In1, RegOut);
 input clk;
 input [23:0] In1;
 output [23 :0] RegOut;

 reg [23 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register15Bit (clk, In1, RegOut);
 input clk;
 input [14:0] In1;
 output [14 :0] RegOut;

 reg [14 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register16Bit (clk, In1, RegOut);
 input clk;
 input [15:0] In1;
 output [15 :0] RegOut;

 reg [15 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register12Bit (clk, In1, RegOut);
 input clk;
 input [11:0] In1;
 output [11 :0] RegOut;

 reg [11 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register13Bit (clk, In1, RegOut);
 input clk;
 input [12:0] In1;
 output [12 :0] RegOut;

 reg [12 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register28Bit (clk, In1, RegOut);
 input clk;
 input [27:0] In1;
 output [27 :0] RegOut;

 reg [27 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule

module Register29Bit (clk, In1, RegOut);
 input clk;
 input [28:0] In1;
 output [28 :0] RegOut;

 reg [28 :0] RegOut; 

always @(posedge clk)
begin
RegOut <= (In1);
end
endmodule



module Negator25Bit (clk, In1, NegOut);
 input clk;
 input [24:0] In1;
 output [24 :0] NegOut;

 reg [24 :0] NegOut; 

always @(posedge clk)
begin
NegOut <= -(In1);
end
endmodule

module Negator23Bit (clk, In1, NegOut);
 input clk;
 input [22:0] In1;
 output [22 :0] NegOut;

 reg [22 :0] NegOut; 

always @(posedge clk)
begin
NegOut <= -(In1);
end
endmodule

module Negator18Bit (clk, In1, NegOut);
 input clk;
 input [17:0] In1;
 output [17 :0] NegOut;

 reg [17 :0] NegOut; 

always @(posedge clk)
begin
NegOut <= -(In1);
end
endmodule

module Negator20Bit (clk, In1, NegOut);
 input clk;
 input [19:0] In1;
 output [19 :0] NegOut;

 reg [19 :0] NegOut; 

always @(posedge clk)
begin
NegOut <= -(In1);
end
endmodule

module Negator19Bit (clk, In1, NegOut);
 input clk;
 input [18:0] In1;
 output [18 :0] NegOut;

 reg [18 :0] NegOut; 

always @(posedge clk)
begin
NegOut <= -(In1);
end
endmodule

module Negator22Bit (clk, In1, NegOut);
 input clk;
 input [21:0] In1;
 output [21 :0] NegOut;

 reg [21 :0] NegOut; 

always @(posedge clk)
begin
NegOut <= -(In1);
end
endmodule

module Negator21Bit (clk, In1, NegOut);
 input clk;
 input [20:0] In1;
 output [20 :0] NegOut;

 reg [20 :0] NegOut; 

always @(posedge clk)
begin
NegOut <= -(In1);
end
endmodule

module Negator24Bit (clk, In1, NegOut);
 input clk;
 input [23:0] In1;
 output [23 :0] NegOut;

 reg [23 :0] NegOut; 

always @(posedge clk)
begin
NegOut <= -(In1);
end
endmodule

module Negator15Bit (clk, In1, NegOut);
 input clk;
 input [14:0] In1;
 output [14 :0] NegOut;

 reg [14 :0] NegOut; 

always @(posedge clk)
begin
NegOut <= -(In1);
end
endmodule

module Negator16Bit (clk, In1, NegOut);
 input clk;
 input [15:0] In1;
 output [15 :0] NegOut;

 reg [15 :0] NegOut; 

always @(posedge clk)
begin
NegOut <= -(In1);
end
endmodule

module Negator17Bit (clk, In1, NegOut);
 input clk;
 input [16:0] In1;
 output [16 :0] NegOut;

 reg [16 :0] NegOut; 

always @(posedge clk)
begin
NegOut <= -(In1);
end
endmodule

module Negator12Bit (clk, In1, NegOut);
 input clk;
 input [11:0] In1;
 output [11 :0] NegOut;

 reg [11 :0] NegOut; 

always @(posedge clk)
begin
NegOut <= -(In1);
end
endmodule
