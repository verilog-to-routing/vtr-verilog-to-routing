/*
 * Integer wide range test
*/

`define WIDTH 32
`define operator buf
`include "range_any_width_unary_test.v"