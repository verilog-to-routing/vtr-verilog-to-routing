module simple_op(a, out);
    input   a;
    output  out;

    buf(out, a);
endmodule