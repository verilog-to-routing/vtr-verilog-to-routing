//////////////////////////////////////////////////////////////////////////////
// Author: Karan Mathur
//////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////
// This benchmark is based on ARM FixyNN DeepFreeze. It accelerates some layers
// of MobileNet.
//////////////////////////////////////////////////////////////////////////////
module top (
    input logic clk,
    input logic rstn,
    input logic valid,
    input logic [24-1:0] input_act,
    output logic [512-1:0] output_act,
    output logic ready
);

logic valid_ff;
logic [24-1:0] input_act_ff;
always_ff @(posedge clk) begin
    if (!rstn) begin
        valid_ff       <= '0;
        input_act_ff   <= '0;
    end
    else begin
        valid_ff       <= valid;
        input_act_ff   <= input_act;
    end
end

logic conv0_buf_valid;
logic [3*72-1:0] conv0_buf_act;
buffer_main #(
    .KER_SIZE (3),
    .BITWIDTH (8),
    .NFMAPS (3),
    .STRIDE (2),
    .PAD (1),
    .NW (224),
    .AW (8)
) conv0_buf_inst (
    .clk (clk),
    .rstn (rstn),
    .valid (valid_ff),
    .D (input_act_ff),
    .Q (conv0_buf_act),
    .ready (conv0_buf_valid)
);

logic conv0_valid;
logic [64-1:0] conv0_act;
conv0 conv0_inst (
    .clk (clk),
    .rstn (rstn),
    .valid (conv0_buf_valid),
    .input_act (conv0_buf_act),
    .output_act (conv0_act),
    .ready (conv0_valid)
);

logic conv1_dw_buf_valid;
logic [8*72-1:0] conv1_dw_buf_act;
buffer_main #(
    .KER_SIZE (3),
    .BITWIDTH (8),
    .NFMAPS (8),
    .STRIDE (1),
    .PAD (1),
    .NW (112),
    .AW (7)
) conv1_dw_buf_inst (
    .clk (clk),
    .rstn (rstn),
    .valid (conv0_valid),
    .D (conv0_act),
    .Q (conv1_dw_buf_act),
    .ready (conv1_dw_buf_valid)
);

logic conv1_dw_valid;
logic [64-1:0] conv1_dw_act;
conv1_dw conv1_dw_inst (
    .clk (clk),
    .rstn (rstn),
    .valid (conv1_dw_buf_valid),
    .input_act (conv1_dw_buf_act),
    .output_act (conv1_dw_act),
    .ready (conv1_dw_valid)
);

logic conv1_pw_buf_valid;

logic  [64-1:0]conv1_pw_buf_act;
assign conv1_pw_buf_act = conv1_dw_act;
assign conv1_pw_buf_valid = conv1_dw_valid ;

logic conv1_pw_valid;
logic [64-1:0] conv1_pw_act;
conv1_pw conv1_pw_inst (
    .clk (clk),
    .rstn (rstn),
    .valid (conv1_pw_buf_valid),
    .input_act (conv1_pw_buf_act),
    .output_act (conv1_pw_act),
    .ready (conv1_pw_valid)
);

logic conv2_dw_buf_valid;
logic [8*72-1:0] conv2_dw_buf_act;
buffer_main #(
    .KER_SIZE (3),
    .BITWIDTH (8),
    .NFMAPS (8),
    .STRIDE (2),
    .PAD (1),
    .NW (112),
    .AW (7)
) conv2_dw_buf_inst (
    .clk (clk),
    .rstn (rstn),
    .valid (conv1_pw_valid),
    .D (conv1_pw_act),
    .Q (conv2_dw_buf_act),
    .ready (conv2_dw_buf_valid)
);

logic conv2_dw_valid;
logic [64-1:0] conv2_dw_act;
conv2_dw conv2_dw_inst (
    .clk (clk),
    .rstn (rstn),
    .valid (conv2_dw_buf_valid),
    .input_act (conv2_dw_buf_act),
    .output_act (conv2_dw_act),
    .ready (conv2_dw_valid)
);

logic conv2_pw_buf_valid;

logic  [64-1:0]conv2_pw_buf_act;
assign conv2_pw_buf_act = conv2_dw_act;
assign conv2_pw_buf_valid = conv2_dw_valid ;

logic conv2_pw_valid;
logic [128-1:0] conv2_pw_act;
conv2_pw conv2_pw_inst (
    .clk (clk),
    .rstn (rstn),
    .valid (conv2_pw_buf_valid),
    .input_act (conv2_pw_buf_act),
    .output_act (conv2_pw_act),
    .ready (conv2_pw_valid)
);

logic conv3_dw_buf_valid;
logic [16*72-1:0] conv3_dw_buf_act;
buffer_main #(
    .KER_SIZE (3),
    .BITWIDTH (8),
    .NFMAPS (16),
    .STRIDE (1),
    .PAD (1),
    .NW (56),
    .AW (6)
) conv3_dw_buf_inst (
    .clk (clk),
    .rstn (rstn),
    .valid (conv2_pw_valid),
    .D (conv2_pw_act),
    .Q (conv3_dw_buf_act),
    .ready (conv3_dw_buf_valid)
);

logic conv3_dw_valid;
logic [128-1:0] conv3_dw_act;
conv3_dw conv3_dw_inst (
    .clk (clk),
    .rstn (rstn),
    .valid (conv3_dw_buf_valid),
    .input_act (conv3_dw_buf_act),
    .output_act (conv3_dw_act),
    .ready (conv3_dw_valid)
);

logic conv3_pw_buf_valid;

logic  [128-1:0]conv3_pw_buf_act;
assign conv3_pw_buf_act = conv3_dw_act;
assign conv3_pw_buf_valid = conv3_dw_valid ;

logic conv3_pw_valid;
logic [128-1:0] conv3_pw_act;
conv3_pw conv3_pw_inst (
    .clk (clk),
    .rstn (rstn),
    .valid (conv3_pw_buf_valid),
    .input_act (conv3_pw_buf_act),
    .output_act (conv3_pw_act),
    .ready (conv3_pw_valid)
);

logic conv4_dw_buf_valid;
logic [16*72-1:0] conv4_dw_buf_act;
buffer_main #(
    .KER_SIZE (3),
    .BITWIDTH (8),
    .NFMAPS (16),
    .STRIDE (2),
    .PAD (1),
    .NW (56),
    .AW (6)
) conv4_dw_buf_inst (
    .clk (clk),
    .rstn (rstn),
    .valid (conv3_pw_valid),
    .D (conv3_pw_act),
    .Q (conv4_dw_buf_act),
    .ready (conv4_dw_buf_valid)
);

logic conv4_dw_valid;
logic [128-1:0] conv4_dw_act;
conv4_dw conv4_dw_inst (
    .clk (clk),
    .rstn (rstn),
    .valid (conv4_dw_buf_valid),
    .input_act (conv4_dw_buf_act),
    .output_act (conv4_dw_act),
    .ready (conv4_dw_valid)
);

logic conv4_pw_buf_valid;

logic  [128-1:0]conv4_pw_buf_act;
assign conv4_pw_buf_act = conv4_dw_act;
assign conv4_pw_buf_valid = conv4_dw_valid ;

logic conv4_pw_valid;
logic [256-1:0] conv4_pw_act;
conv4_pw conv4_pw_inst (
    .clk (clk),
    .rstn (rstn),
    .valid (conv4_pw_buf_valid),
    .input_act (conv4_pw_buf_act),
    .output_act (conv4_pw_act),
    .ready (conv4_pw_valid)
);

logic conv5_dw_buf_valid;
logic [32*72-1:0] conv5_dw_buf_act;
buffer_main #(
    .KER_SIZE (3),
    .BITWIDTH (8),
    .NFMAPS (32),
    .STRIDE (1),
    .PAD (1),
    .NW (28),
    .AW (5)
) conv5_dw_buf_inst (
    .clk (clk),
    .rstn (rstn),
    .valid (conv4_pw_valid),
    .D (conv4_pw_act),
    .Q (conv5_dw_buf_act),
    .ready (conv5_dw_buf_valid)
);

logic conv5_dw_valid;
logic [256-1:0] conv5_dw_act;
conv5_dw conv5_dw_inst (
    .clk (clk),
    .rstn (rstn),
    .valid (conv5_dw_buf_valid),
    .input_act (conv5_dw_buf_act),
    .output_act (conv5_dw_act),
    .ready (conv5_dw_valid)
);

logic conv5_pw_buf_valid;

logic  [256-1:0]conv5_pw_buf_act;
assign conv5_pw_buf_act = conv5_dw_act;
assign conv5_pw_buf_valid = conv5_dw_valid ;

logic conv5_pw_valid;
logic [256-1:0] conv5_pw_act;
conv5_pw conv5_pw_inst (
    .clk (clk),
    .rstn (rstn),
    .valid (conv5_pw_buf_valid),
    .input_act (conv5_pw_buf_act),
    .output_act (conv5_pw_act),
    .ready (conv5_pw_valid)
);

logic conv6_dw_buf_valid;
logic [32*72-1:0] conv6_dw_buf_act;
buffer_main #(
    .KER_SIZE (3),
    .BITWIDTH (8),
    .NFMAPS (32),
    .STRIDE (2),
    .PAD (1),
    .NW (28),
    .AW (5)
) conv6_dw_buf_inst (
    .clk (clk),
    .rstn (rstn),
    .valid (conv5_pw_valid),
    .D (conv5_pw_act),
    .Q (conv6_dw_buf_act),
    .ready (conv6_dw_buf_valid)
);

logic conv6_dw_valid;
logic [256-1:0] conv6_dw_act;
conv6_dw conv6_dw_inst (
    .clk (clk),
    .rstn (rstn),
    .valid (conv6_dw_buf_valid),
    .input_act (conv6_dw_buf_act),
    .output_act (conv6_dw_act),
    .ready (conv6_dw_valid)
);

logic conv6_pw_buf_valid;

logic  [256-1:0]conv6_pw_buf_act;
assign conv6_pw_buf_act = conv6_dw_act;
assign conv6_pw_buf_valid = conv6_dw_valid ;

logic conv6_pw_valid;
logic [512-1:0] conv6_pw_act;
conv6_pw conv6_pw_inst (
    .clk (clk),
    .rstn (rstn),
    .valid (conv6_pw_buf_valid),
    .input_act (conv6_pw_buf_act),
    .output_act (conv6_pw_act),
    .ready (conv6_pw_valid)
);

logic conv7_dw_buf_valid;
logic [64*72-1:0] conv7_dw_buf_act;
buffer_main #(
    .KER_SIZE (3),
    .BITWIDTH (8),
    .NFMAPS (64),
    .STRIDE (1),
    .PAD (1),
    .NW (14),
    .AW (4)
) conv7_dw_buf_inst (
    .clk (clk),
    .rstn (rstn),
    .valid (conv6_pw_valid),
    .D (conv6_pw_act),
    .Q (conv7_dw_buf_act),
    .ready (conv7_dw_buf_valid)
);

logic conv7_dw_valid;
logic [512-1:0] conv7_dw_act;
conv7_dw conv7_dw_inst (
    .clk (clk),
    .rstn (rstn),
    .valid (conv7_dw_buf_valid),
    .input_act (conv7_dw_buf_act),
    .output_act (conv7_dw_act),
    .ready (conv7_dw_valid)
);

logic conv7_pw_buf_valid;

logic  [512-1:0]conv7_pw_buf_act;
assign conv7_pw_buf_act = conv7_dw_act;
assign conv7_pw_buf_valid = conv7_dw_valid ;

logic conv7_pw_valid;
logic [512-1:0] conv7_pw_act;
conv7_pw conv7_pw_inst (
    .clk (clk),
    .rstn (rstn),
    .valid (conv7_pw_buf_valid),
    .input_act (conv7_pw_buf_act),
    .output_act (conv7_pw_act),
    .ready (conv7_pw_valid)
);

logic conv8_dw_buf_valid;
logic [64*72-1:0] conv8_dw_buf_act;
buffer_main #(
    .KER_SIZE (3),
    .BITWIDTH (8),
    .NFMAPS (64),
    .STRIDE (1),
    .PAD (1),
    .NW (14),
    .AW (4)
) conv8_dw_buf_inst (
    .clk (clk),
    .rstn (rstn),
    .valid (conv7_pw_valid),
    .D (conv7_pw_act),
    .Q (conv8_dw_buf_act),
    .ready (conv8_dw_buf_valid)
);

logic conv8_dw_valid;
logic [512-1:0] conv8_dw_act;
conv8_dw conv8_dw_inst (
    .clk (clk),
    .rstn (rstn),
    .valid (conv8_dw_buf_valid),
    .input_act (conv8_dw_buf_act),
    .output_act (conv8_dw_act),
    .ready (conv8_dw_valid)
);

logic conv8_pw_buf_valid;

logic  [512-1:0]conv8_pw_buf_act;
assign conv8_pw_buf_act = conv8_dw_act;
assign conv8_pw_buf_valid = conv8_dw_valid ;

logic conv8_pw_valid;
logic [512-1:0] conv8_pw_act;
conv8_pw conv8_pw_inst (
    .clk (clk),
    .rstn (rstn),
    .valid (conv8_pw_buf_valid),
    .input_act (conv8_pw_buf_act),
    .output_act (conv8_pw_act),
    .ready (conv8_pw_valid)
);

always_ff @(posedge clk) begin
    if (!rstn) begin
        output_act <= '0;
        ready      <= '0;
    end
    else begin
        output_act <= conv8_pw_act;
        ready      <= conv8_pw_valid;
    end
end

endmodule

module buffer_main
#(
    parameter KER_SIZE = 3,
    parameter BITWIDTH = 8,
    parameter NFMAPS   = 3,
    parameter STRIDE   = 1,
    parameter PAD      = 1,
    parameter NW       = 32,
    parameter AW       = $clog2(NW)
)
(
    input logic clk,
    input logic rstn,
    input logic valid,
    input logic [NFMAPS*BITWIDTH-1:0] D,
    //output logic [KER_SIZE*KER_SIZE*BITWIDTH-1:0] Q [NFMAPS-1:0],
    output logic [NFMAPS*KER_SIZE*KER_SIZE*BITWIDTH-1:0] Q,
    output logic ready
);

localparam DW = NFMAPS*BITWIDTH;
genvar i,j;

logic [AW-1:0] address_wire                                            ;
logic [KER_SIZE-1:0] write_en_wire                                     ;
logic [KER_SIZE-1:0] read_en_wire                                      ; 
logic [(KER_SIZE)*DW-1:0] sram_read_data_wire                          ;
logic [(KER_SIZE-1)*DW-1:0] sram_km1_read_data                         ; //kernel size - 1 read data coming from SRAM
logic [DW-1:0] incoming_px                                             ; //incoming_pixel
logic [DW-1:0] incoming_px_D1                                          ; //incoming_pixel_delayed

//logic [DW-1:0] sram_read_data_rowwise [KER_SIZE-1:0]                   ;
logic [KER_SIZE*DW-1:0] sram_read_data_rowwise;

//logic [KER_SIZE*BITWIDTH-1:0] pixel_in_fmap_wise [NFMAPS-1:0]          ;
logic [NFMAPS*KER_SIZE*BITWIDTH-1:0] pixel_in_fmap_wise;

//logic [KER_SIZE*KER_SIZE*BITWIDTH-1:0] pixel_out_fmap_wise [NFMAPS-1:0];
logic [NFMAPS*KER_SIZE*KER_SIZE*BITWIDTH-1:0] pixel_out_fmap_wise;
logic [3-1:0] col_ptr_wire                                             ;
logic [3-1:0] init_col_ptr_wire                                        ;
logic [3-1:0] col_stride_counter                                       ;
logic [3-1:0] col_stride_counter_nxt                                   ;
logic sram_is_ready,sram_is_ready_D1                                   ;
logic valid_D1                                                         ;
logic ready_wire                                                       ;
logic line_buf_is_ready                                                ;
//PAD signals
logic right_pad_valid                                                  ;
logic bottom_pad_mask                                                  ;
logic [KER_SIZE-1:0] top_pad_mask	                                     ;
logic [KER_SIZE-1:0] left_pad_mask	                                   ;
logic [KER_SIZE-1:0] right_pad_mask	                                   ;
//input flops
logic valid_reg                                                        ;
logic [NFMAPS*BITWIDTH-1:0]D_reg                                       ;
logic row_complete_wire                                                ;
 
assign valid_reg = valid;
assign D_reg = bottom_pad_mask ? D & {NFMAPS*BITWIDTH{1'b0}} : D; //mask dummy data as zeros at bottom pad
assign incoming_px = D_reg;

// delay for incoming new row
always_ff @(posedge clk) 
begin
    if (!rstn) 
        incoming_px_D1 			<= 0;
    else if(sram_is_ready) 
        incoming_px_D1 			<= incoming_px;
    else 
        incoming_px_D1 			<= 0;
end

sram_controller #(
    .KER_SIZE 		(KER_SIZE	),
    .BITWIDTH 		(BITWIDTH	),
    .STRIDE 			(STRIDE		),
    .PAD 					(PAD			),
    .NFMAPS 			(NFMAPS		),
    .INPUT_X_DIM 	(NW				),
    .AW 					(AW				)
) sram_ctrl_inst (
    .clk 			 				(clk							),
    .rstn 			 			(rstn							),
    .valid 			 			(valid_reg				),
    .addr 			 			(address_wire			),
    .write_en 				(write_en_wire		),
    .read_en 		 			(read_en_wire 		),
    .row_is_complete 	(row_complete_wire),
		.top_pad_mask	 		(top_pad_mask			),
		.bottom_pad_mask 	(bottom_pad_mask	),
    .ready 			 			(sram_is_ready		)
);

// TODO: generalize sram array module to different kernel sizes
generate
if (KER_SIZE == 3)
begin
    sram_array_k3 #(
        .KER_SIZE (KER_SIZE),
        .DW 			(DW			),
        .NW 			(NW			),
        .AW 			(AW			)
    ) sram_array_k3_inst (
        .clk 	(clk								),
        .rstn (rstn								),
        .a 		(address_wire				),
        .wen 	(write_en_wire			),
        .ren 	(read_en_wire				),
        .d 		(D_reg							),
        .q 		(sram_km1_read_data	)
    );
		assign sram_read_data_wire = {incoming_px_D1,sram_km1_read_data};
end    
else if (KER_SIZE == 2) 
begin
    sram_array_k2 #(
        .KER_SIZE (KER_SIZE),
        .DW 			(DW),
        .NW 			(NW),
        .AW 			(AW)
    ) sram_array_k2_inst (
        .clk 	(clk								),
        .rstn (rstn								),
        .a 		(address_wire				),
        .wen 	(write_en_wire			),
        .ren 	(read_en_wire				),
        .d 		(D_reg							),
        .q 		(sram_km1_read_data	)
    );
		assign sram_read_data_wire = {incoming_px_D1,sram_km1_read_data};
 end        
else if(KER_SIZE == 5)
begin
    sram_array_k5 #(
         .KER_SIZE (KER_SIZE),
         .DW 			 (DW			),
         .NW 			 (NW			),
         .AW 			 (AW			)
    ) sram_array_k5_inst (
        .clk 	(clk								),
        .rstn (rstn								),
        .a 		(address_wire				),
        .wen 	(write_en_wire			),
        .ren 	(read_en_wire				),
        .d 		(D_reg							),
        .q 		(sram_km1_read_data	)
    );
		assign sram_read_data_wire = {incoming_px_D1,sram_km1_read_data};
end        
else if(KER_SIZE == 7)
begin
    sram_array_k7 #(
         .KER_SIZE (KER_SIZE),
         .DW 			 (DW			),
         .NW 			 (NW			),
         .AW 			 (AW			)
    ) sram_array_k7_inst (
        .clk 	(clk								),
        .rstn (rstn								),
        .a 		(address_wire				),
        .wen 	(write_en_wire			),
        .ren 	(read_en_wire				),
        .d 		(D_reg							),
        .q 		(sram_km1_read_data	)
    );
		assign sram_read_data_wire = {incoming_px_D1,sram_km1_read_data};
end 
endgenerate

// delay for sram read cycle, sram data is ready after a cycle when sram is ready
always_ff @(posedge clk) begin
    if (!rstn) begin
        valid_D1 			    <= '0;
        sram_is_ready_D1 	<= '0;
    end
    else begin
        valid_D1 			    <= valid_reg;
        sram_is_ready_D1 	<= sram_is_ready;
    end
end

line_buffer_controller #(
    .KER_SIZE 		(KER_SIZE	),
    .INPUT_X_DIM 	(NW			),
    .PAD 			(PAD		)
) line_buffer_controller_inst (
    .clk 						  (clk													),
    .rstn 					  (rstn													),
    .valid 					  (valid_D1 && sram_is_ready_D1	),
    .row_complete 		(row_complete_wire						),
    .col_ptr 			    (col_ptr_wire									),
    .right_pad_valid 	(right_pad_valid							),
    .left_pad_mask 		(left_pad_mask								),
    .right_pad_mask 	(right_pad_mask								),
    .init_col_ptr 		(init_col_ptr_wire						)
);

generate
    for (i = 0; i < KER_SIZE; i++) begin: genblk_0
    always@(posedge clk) begin 
       sram_read_data_rowwise[(i+1)*DW-1:i*DW] = sram_read_data_wire [(i+1)*DW-1:(i*DW)] & {KER_SIZE*DW{!top_pad_mask[i]}};
    end   
    end

    for (j = 0; j < NFMAPS; j++) begin: genblk_1
        for (i = 0; i < KER_SIZE; i++) begin: genblk_2
        always@(posedge clk) begin 
            pixel_in_fmap_wise[(j*KER_SIZE*BITWIDTH + i*BITWIDTH)+:BITWIDTH] = sram_read_data_rowwise[(j*KER_SIZE*BITWIDTH + i*BITWIDTH)+:BITWIDTH];
        end    
        end
    end

    // TODO: generalize line buffer arrays to different kernel sizes
    for (i = 0; i < NFMAPS; i++) begin: genblk_3
        if (KER_SIZE == 3) begin
            line_buffer_array_k3 #      (
                .KER_SIZE               (KER_SIZE),
                .BITWIDTH               (BITWIDTH),
								.PAD                    (PAD),
                .AW 		                (AW)) 
								line_buffer_array_k3_inst (
                .clk                    (clk),
                .rstn                   (rstn),
                .pixel_in               (pixel_in_fmap_wise[(i+1)*KER_SIZE*BITWIDTH-1:i*KER_SIZE*BITWIDTH]),
                .col_ptr                (col_ptr_wire),
                .init_col_ptr           (init_col_ptr_wire),
								.left_pad_mask 	        (left_pad_mask),
								.right_pad_mask         (right_pad_mask),
                .pixel_out              (pixel_out_fmap_wise[(i+1)*KER_SIZE*KER_SIZE*BITWIDTH-1:i*KER_SIZE*KER_SIZE*BITWIDTH])
            );
        end
        else if (KER_SIZE == 2) begin
            line_buffer_array_k2 #      (
                .KER_SIZE               (KER_SIZE),
                .BITWIDTH               (BITWIDTH),
                .AW                     (AW)
            ) line_buffer_array_k2_inst (
                .clk                    (clk),
                .rstn                   (rstn),
                .pixel_in               (pixel_in_fmap_wise [(i+1)*KER_SIZE*BITWIDTH-1:i*KER_SIZE*BITWIDTH]),
                .col_ptr                (col_ptr_wire),
                .init_col_ptr           (init_col_ptr_wire),
                .pixel_out              (pixel_out_fmap_wise [(i+1)*KER_SIZE*KER_SIZE*BITWIDTH-1:i*KER_SIZE*KER_SIZE*BITWIDTH])
            );
        end
        else if (KER_SIZE == 5) begin
            line_buffer_array_k5 #      (
                .KER_SIZE               (KER_SIZE),
                .PAD                    (PAD),
                .BITWIDTH               (BITWIDTH),
                .AW                     (AW)
            ) line_buffer_array_k5_inst (
                .clk 			              (clk),
                .rstn 			            (rstn),
                .pixel_in 		          (pixel_in_fmap_wise [(i+1)*KER_SIZE*BITWIDTH-1:i*KER_SIZE*BITWIDTH]),
                .col_ptr 		            (col_ptr_wire),
                .init_col_ptr 	        (init_col_ptr_wire),
                .left_pad_mask 	        (left_pad_mask),
                .right_pad_mask         (right_pad_mask),
                .pixel_out 		          (pixel_out_fmap_wise [(i+1)*KER_SIZE*KER_SIZE*BITWIDTH-1:i*KER_SIZE*KER_SIZE*BITWIDTH])
            );
        end
        else if (KER_SIZE == 7) begin
            line_buffer_array_k7 #      (
                .KER_SIZE               (KER_SIZE),
                .PAD                    (PAD),
                .BITWIDTH               (BITWIDTH),
                .AW                     (AW)
            ) line_buffer_array_k7_inst (
                .clk 			              (clk),
                .rstn 			            (rstn),
                .pixel_in 		          (pixel_in_fmap_wise [(i+1)*KER_SIZE*BITWIDTH-1:i*KER_SIZE*BITWIDTH]),
                .col_ptr 		            (col_ptr_wire),
                .init_col_ptr 	        (init_col_ptr_wire),
                .left_pad_mask 	        (left_pad_mask),
                .right_pad_mask         (right_pad_mask),
                .pixel_out 		          (pixel_out_fmap_wise [(i+1)*KER_SIZE*KER_SIZE*BITWIDTH-1:i*KER_SIZE*KER_SIZE*BITWIDTH])
            );
        end
    end

    for (i = 0; i < NFMAPS; i++) begin: genblk_4
        assign Q[(i+1)*KER_SIZE*KER_SIZE*BITWIDTH-1:(i*KER_SIZE*KER_SIZE*BITWIDTH)] = pixel_out_fmap_wise[(i+1)*KER_SIZE*KER_SIZE*BITWIDTH-1:i*KER_SIZE*KER_SIZE*BITWIDTH];
    end

endgenerate

// ready_logic
always_ff @(posedge clk) begin
    if (!rstn) begin
        col_stride_counter <= '0;
    end
    else if (row_complete_wire) begin
        col_stride_counter <= '0;
    end
    else begin
        col_stride_counter <= col_stride_counter_nxt;
    end
end

// because of one cycle delay of line buffer
always_ff @(posedge clk) begin
    if (!rstn) begin
        ready_wire <= '0;
    end
    else begin
        ready_wire <= (col_stride_counter==0) && (line_buf_is_ready);
    end
end

assign line_buf_is_ready = (init_col_ptr_wire == KER_SIZE-1 && valid_D1);
assign col_stride_counter_nxt = (line_buf_is_ready) ? ((col_stride_counter<STRIDE-1'd1)?col_stride_counter+1'd1:'0 ): col_stride_counter;
assign ready = ready_wire || right_pad_valid;

endmodule


module conv0 (
    input logic clk,
    input logic rstn,
    input logic valid,
    input logic [3*72-1:0] input_act,
    output logic [64-1:0] output_act,
    output logic ready
);
logic we;
logic [8:0] zero_number; 
assign zero_number = 9'd0; 
logic [3*72-1:0] input_act_ff;
genvar i;
generate
for (i=0;i<3;i++)
    begin: genblk_5
        always_ff @(posedge clk) begin
            if (rstn == 0) begin
                input_act_ff[(i+1)*72-1:i*72] <= '0;
            end
            else begin
                input_act_ff[(i+1)*72-1:i*72] <= input_act[(i+1)*72-1:i*72];
            end
        end
    end
endgenerate
logic [71:0] input_fmap_0;
assign input_fmap_0 = input_act_ff[71:0];
logic [71:0] input_fmap_1;
assign input_fmap_1 = input_act_ff[143:72];
logic [71:0] input_fmap_2;
assign input_fmap_2 = input_act_ff[215:144];

logic [10-1:0] O0_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O0_I0_R0_C01_rom_inst (.q(O0_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O0_I0_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O0_I0_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O0_I0_R0_C01_rom_inst (.q(O0_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [10-1:0] O0_I0_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O0_I0_R0_C11_rom_inst (.q(O0_I0_R0_C1_SM1 ),.address(input_fmap_0[15:8]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R0_C1_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O0_I0_R0_C1_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O0_I0_R0_C11_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O0_I0_R0_C11_rom_inst (.q(O0_I0_R0_C1_SM1 ),.address(input_fmap_0[15:8]),.clock  (clk));
logic [10-1:0] O0_I0_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O0_I0_R0_C21_rom_inst (.q(O0_I0_R0_C2_SM1 ),.address(input_fmap_0[23:16]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R0_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O0_I0_R0_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O0_I0_R0_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O0_I0_R0_C21_rom_inst (.q(O0_I0_R0_C2_SM1 ),.address(input_fmap_0[23:16]),.clock  (clk));
logic [11-1:0] O0_I0_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O0_I0_R1_C02_rom_inst (.q(O0_I0_R1_C0_SM1 ),.address(input_fmap_0[31:24]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R1_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O0_I0_R1_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O0_I0_R1_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O0_I0_R1_C02_rom_inst (.q(O0_I0_R1_C0_SM1 ),.address(input_fmap_0[31:24]),.clock  (clk));
logic [11-1:0] O0_I0_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O0_I0_R1_C13_rom_inst (.q(O0_I0_R1_C1_SM1 ),.address(input_fmap_0[39:32]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R1_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O0_I0_R1_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O0_I0_R1_C13_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O0_I0_R1_C13_rom_inst (.q(O0_I0_R1_C1_SM1 ),.address(input_fmap_0[39:32]),.clock  (clk));
logic [11-1:0] O0_I0_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O0_I0_R1_C22_rom_inst (.q(O0_I0_R1_C2_SM1 ),.address(input_fmap_0[47:40]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R1_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O0_I0_R1_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O0_I0_R1_C22_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O0_I0_R1_C22_rom_inst (.q(O0_I0_R1_C2_SM1 ),.address(input_fmap_0[47:40]),.clock  (clk));
logic [11-1:0] O0_I0_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O0_I0_R2_C02_rom_inst (.q(O0_I0_R2_C0_SM1 ),.address(input_fmap_0[55:48]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R2_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O0_I0_R2_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O0_I0_R2_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O0_I0_R2_C02_rom_inst (.q(O0_I0_R2_C0_SM1 ),.address(input_fmap_0[55:48]),.clock  (clk));
logic [11-1:0] O0_I0_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O0_I0_R2_C12_rom_inst (.q(O0_I0_R2_C1_SM1 ),.address(input_fmap_0[63:56]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R2_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O0_I0_R2_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O0_I0_R2_C12_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O0_I0_R2_C12_rom_inst (.q(O0_I0_R2_C1_SM1 ),.address(input_fmap_0[63:56]),.clock  (clk));
logic [10-1:0] O0_I0_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O0_I0_R2_C21_rom_inst (.q(O0_I0_R2_C2_SM1 ),.address(input_fmap_0[71:64]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R2_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O0_I0_R2_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O0_I0_R2_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O0_I0_R2_C21_rom_inst (.q(O0_I0_R2_C2_SM1 ),.address(input_fmap_0[71:64]),.clock  (clk));
logic [11-1:0] O0_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O0_I1_R0_C03_rom_inst (.q(O0_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I1_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O0_I1_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O0_I1_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O0_I1_R0_C03_rom_inst (.q(O0_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [12-1:0] O0_I1_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv0_O0_I1_R0_C14_rom_inst (.q(O0_I1_R0_C1_SM1 ),.address(input_fmap_1[15:8]),.clk(clk),.d(0),.we(0));
//assign O0_I1_R0_C1_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O0_I1_R0_C1_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O0_I1_R0_C14_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv0_O0_I1_R0_C14_rom_inst (.q(O0_I1_R0_C1_SM1 ),.address(input_fmap_1[15:8]),.clock  (clk));
logic [11-1:0] O0_I1_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O0_I1_R0_C23_rom_inst (.q(O0_I1_R0_C2_SM1 ),.address(input_fmap_1[23:16]),.clk(clk),.d(0),.we(0));
//assign O0_I1_R0_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O0_I1_R0_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O0_I1_R0_C23_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O0_I1_R0_C23_rom_inst (.q(O0_I1_R0_C2_SM1 ),.address(input_fmap_1[23:16]),.clock  (clk));
logic [11-1:0] O0_I1_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O0_I1_R1_C03_rom_inst (.q(O0_I1_R1_C0_SM1 ),.address(input_fmap_1[31:24]),.clk(clk),.d(0),.we(0));
//assign O0_I1_R1_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O0_I1_R1_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O0_I1_R1_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O0_I1_R1_C03_rom_inst (.q(O0_I1_R1_C0_SM1 ),.address(input_fmap_1[31:24]),.clock  (clk));
logic [11-1:0] O0_I1_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O0_I1_R1_C13_rom_inst (.q(O0_I1_R1_C1_SM1 ),.address(input_fmap_1[39:32]),.clk(clk),.d(0),.we(0));
//assign O0_I1_R1_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O0_I1_R1_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O0_I1_R1_C13_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O0_I1_R1_C13_rom_inst (.q(O0_I1_R1_C1_SM1 ),.address(input_fmap_1[39:32]),.clock  (clk));
logic [12-1:0] O0_I1_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv0_O0_I1_R1_C24_rom_inst (.q(O0_I1_R1_C2_SM1 ),.address(input_fmap_1[47:40]),.clk(clk),.d(0),.we(0));
//assign O0_I1_R1_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O0_I1_R1_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O0_I1_R1_C24_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv0_O0_I1_R1_C24_rom_inst (.q(O0_I1_R1_C2_SM1 ),.address(input_fmap_1[47:40]),.clock  (clk));
logic [12-1:0] O0_I1_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv0_O0_I1_R2_C04_rom_inst (.q(O0_I1_R2_C0_SM1 ),.address(input_fmap_1[55:48]),.clk(clk),.d(0),.we(0));
//assign O0_I1_R2_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O0_I1_R2_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O0_I1_R2_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv0_O0_I1_R2_C04_rom_inst (.q(O0_I1_R2_C0_SM1 ),.address(input_fmap_1[55:48]),.clock  (clk));
logic [12-1:0] O0_I1_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv0_O0_I1_R2_C14_rom_inst (.q(O0_I1_R2_C1_SM1 ),.address(input_fmap_1[63:56]),.clk(clk),.d(0),.we(0));
//assign O0_I1_R2_C1_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O0_I1_R2_C1_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O0_I1_R2_C14_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv0_O0_I1_R2_C14_rom_inst (.q(O0_I1_R2_C1_SM1 ),.address(input_fmap_1[63:56]),.clock  (clk));
logic [12-1:0] O0_I1_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv0_O0_I1_R2_C25_rom_inst (.q(O0_I1_R2_C2_SM1 ),.address(input_fmap_1[71:64]),.clk(clk),.d(0),.we(0));
//assign O0_I1_R2_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O0_I1_R2_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O0_I1_R2_C25_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv0_O0_I1_R2_C25_rom_inst (.q(O0_I1_R2_C2_SM1 ),.address(input_fmap_1[71:64]),.clock  (clk));
logic [11-1:0] O0_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O0_I2_R0_C02_rom_inst (.q(O0_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I2_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O0_I2_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O0_I2_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O0_I2_R0_C02_rom_inst (.q(O0_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [11-1:0] O0_I2_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O0_I2_R0_C12_rom_inst (.q(O0_I2_R0_C1_SM1 ),.address(input_fmap_2[15:8]),.clk(clk),.d(0),.we(0));
//assign O0_I2_R0_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O0_I2_R0_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O0_I2_R0_C12_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O0_I2_R0_C12_rom_inst (.q(O0_I2_R0_C1_SM1 ),.address(input_fmap_2[15:8]),.clock  (clk));
logic [11-1:0] O0_I2_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O0_I2_R0_C22_rom_inst (.q(O0_I2_R0_C2_SM1 ),.address(input_fmap_2[23:16]),.clk(clk),.d(0),.we(0));
//assign O0_I2_R0_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O0_I2_R0_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O0_I2_R0_C22_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O0_I2_R0_C22_rom_inst (.q(O0_I2_R0_C2_SM1 ),.address(input_fmap_2[23:16]),.clock  (clk));
logic [11-1:0] O0_I2_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O0_I2_R1_C02_rom_inst (.q(O0_I2_R1_C0_SM1 ),.address(input_fmap_2[31:24]),.clk(clk),.d(0),.we(0));
//assign O0_I2_R1_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O0_I2_R1_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O0_I2_R1_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O0_I2_R1_C02_rom_inst (.q(O0_I2_R1_C0_SM1 ),.address(input_fmap_2[31:24]),.clock  (clk));
logic [11-1:0] O0_I2_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O0_I2_R1_C13_rom_inst (.q(O0_I2_R1_C1_SM1 ),.address(input_fmap_2[39:32]),.clk(clk),.d(0),.we(0));
//assign O0_I2_R1_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O0_I2_R1_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O0_I2_R1_C13_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O0_I2_R1_C13_rom_inst (.q(O0_I2_R1_C1_SM1 ),.address(input_fmap_2[39:32]),.clock  (clk));
logic [11-1:0] O0_I2_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O0_I2_R1_C22_rom_inst (.q(O0_I2_R1_C2_SM1 ),.address(input_fmap_2[47:40]),.clk(clk),.d(0),.we(0));
//assign O0_I2_R1_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O0_I2_R1_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O0_I2_R1_C22_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O0_I2_R1_C22_rom_inst (.q(O0_I2_R1_C2_SM1 ),.address(input_fmap_2[47:40]),.clock  (clk));
logic [11-1:0] O0_I2_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O0_I2_R2_C02_rom_inst (.q(O0_I2_R2_C0_SM1 ),.address(input_fmap_2[55:48]),.clk(clk),.d(0),.we(0));
//assign O0_I2_R2_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O0_I2_R2_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O0_I2_R2_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O0_I2_R2_C02_rom_inst (.q(O0_I2_R2_C0_SM1 ),.address(input_fmap_2[55:48]),.clock  (clk));
logic [11-1:0] O0_I2_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O0_I2_R2_C13_rom_inst (.q(O0_I2_R2_C1_SM1 ),.address(input_fmap_2[63:56]),.clk(clk),.d(0),.we(0));
//assign O0_I2_R2_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O0_I2_R2_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O0_I2_R2_C13_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O0_I2_R2_C13_rom_inst (.q(O0_I2_R2_C1_SM1 ),.address(input_fmap_2[63:56]),.clock  (clk));
logic [11-1:0] O0_I2_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O0_I2_R2_C22_rom_inst (.q(O0_I2_R2_C2_SM1 ),.address(input_fmap_2[71:64]),.clk(clk),.d(0),.we(0));
//assign O0_I2_R2_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O0_I2_R2_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O0_I2_R2_C22_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O0_I2_R2_C22_rom_inst (.q(O0_I2_R2_C2_SM1 ),.address(input_fmap_2[71:64]),.clock  (clk));
logic [11-1:0] O1_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O1_I0_R0_C03_rom_inst (.q(O1_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I0_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O1_I0_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O1_I0_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O1_I0_R0_C03_rom_inst (.q(O1_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [12-1:0] O1_I0_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv0_O1_I0_R0_C14_rom_inst (.q(O1_I0_R0_C1_SM1 ),.address(input_fmap_0[15:8]),.clk(clk),.d(0),.we(0));
//assign O1_I0_R0_C1_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O1_I0_R0_C1_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O1_I0_R0_C14_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv0_O1_I0_R0_C14_rom_inst (.q(O1_I0_R0_C1_SM1 ),.address(input_fmap_0[15:8]),.clock  (clk));
logic [11-1:0] O1_I0_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O1_I0_R0_C22_rom_inst (.q(O1_I0_R0_C2_SM1 ),.address(input_fmap_0[23:16]),.clk(clk),.d(0),.we(0));
//assign O1_I0_R0_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O1_I0_R0_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O1_I0_R0_C22_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O1_I0_R0_C22_rom_inst (.q(O1_I0_R0_C2_SM1 ),.address(input_fmap_0[23:16]),.clock  (clk));
logic [10-1:0] O1_I0_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O1_I0_R1_C01_rom_inst (.q(O1_I0_R1_C0_SM1 ),.address(input_fmap_0[31:24]),.clk(clk),.d(0),.we(0));
//assign O1_I0_R1_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O1_I0_R1_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O1_I0_R1_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O1_I0_R1_C01_rom_inst (.q(O1_I0_R1_C0_SM1 ),.address(input_fmap_0[31:24]),.clock  (clk));
logic [10-1:0] O1_I0_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O1_I0_R1_C11_rom_inst (.q(O1_I0_R1_C1_SM1 ),.address(input_fmap_0[39:32]),.clk(clk),.d(0),.we(0));
//assign O1_I0_R1_C1_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O1_I0_R1_C1_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O1_I0_R1_C11_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O1_I0_R1_C11_rom_inst (.q(O1_I0_R1_C1_SM1 ),.address(input_fmap_0[39:32]),.clock  (clk));
logic [10-1:0] O1_I0_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O1_I0_R1_C21_rom_inst (.q(O1_I0_R1_C2_SM1 ),.address(input_fmap_0[47:40]),.clk(clk),.d(0),.we(0));
//assign O1_I0_R1_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O1_I0_R1_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O1_I0_R1_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O1_I0_R1_C21_rom_inst (.q(O1_I0_R1_C2_SM1 ),.address(input_fmap_0[47:40]),.clock  (clk));
logic [11-1:0] O1_I0_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O1_I0_R2_C03_rom_inst (.q(O1_I0_R2_C0_SM1 ),.address(input_fmap_0[55:48]),.clk(clk),.d(0),.we(0));
//assign O1_I0_R2_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O1_I0_R2_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O1_I0_R2_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O1_I0_R2_C03_rom_inst (.q(O1_I0_R2_C0_SM1 ),.address(input_fmap_0[55:48]),.clock  (clk));
logic [12-1:0] O1_I0_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv0_O1_I0_R2_C15_rom_inst (.q(O1_I0_R2_C1_SM1 ),.address(input_fmap_0[63:56]),.clk(clk),.d(0),.we(0));
//assign O1_I0_R2_C1_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O1_I0_R2_C1_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O1_I0_R2_C15_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv0_O1_I0_R2_C15_rom_inst (.q(O1_I0_R2_C1_SM1 ),.address(input_fmap_0[63:56]),.clock  (clk));
logic [11-1:0] O1_I0_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O1_I0_R2_C22_rom_inst (.q(O1_I0_R2_C2_SM1 ),.address(input_fmap_0[71:64]),.clk(clk),.d(0),.we(0));
//assign O1_I0_R2_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O1_I0_R2_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O1_I0_R2_C22_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O1_I0_R2_C22_rom_inst (.q(O1_I0_R2_C2_SM1 ),.address(input_fmap_0[71:64]),.clock  (clk));
logic [12-1:0] O1_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv0_O1_I1_R0_C06_rom_inst (.q(O1_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O1_I1_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O1_I1_R0_C06_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv0_O1_I1_R0_C06_rom_inst (.q(O1_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [13-1:0] O1_I1_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv0_O1_I1_R0_C18_rom_inst (.q(O1_I1_R0_C1_SM1 ),.address(input_fmap_1[15:8]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R0_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O1_I1_R0_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O1_I1_R0_C18_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv0_O1_I1_R0_C18_rom_inst (.q(O1_I1_R0_C1_SM1 ),.address(input_fmap_1[15:8]),.clock  (clk));
logic [11-1:0] O1_I1_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O1_I1_R0_C23_rom_inst (.q(O1_I1_R0_C2_SM1 ),.address(input_fmap_1[23:16]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R0_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O1_I1_R0_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O1_I1_R0_C23_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O1_I1_R0_C23_rom_inst (.q(O1_I1_R0_C2_SM1 ),.address(input_fmap_1[23:16]),.clock  (clk));
logic [11-1:0] O1_I1_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O1_I1_R1_C02_rom_inst (.q(O1_I1_R1_C0_SM1 ),.address(input_fmap_1[31:24]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R1_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O1_I1_R1_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O1_I1_R1_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O1_I1_R1_C02_rom_inst (.q(O1_I1_R1_C0_SM1 ),.address(input_fmap_1[31:24]),.clock  (clk));
logic [10-1:0] O1_I1_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O1_I1_R1_C11_rom_inst (.q(O1_I1_R1_C1_SM1 ),.address(input_fmap_1[39:32]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R1_C1_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O1_I1_R1_C1_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O1_I1_R1_C11_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O1_I1_R1_C11_rom_inst (.q(O1_I1_R1_C1_SM1 ),.address(input_fmap_1[39:32]),.clock  (clk));
logic [10-1:0] O1_I1_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O1_I1_R1_C21_rom_inst (.q(O1_I1_R1_C2_SM1 ),.address(input_fmap_1[47:40]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R1_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O1_I1_R1_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O1_I1_R1_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O1_I1_R1_C21_rom_inst (.q(O1_I1_R1_C2_SM1 ),.address(input_fmap_1[47:40]),.clock  (clk));
logic [12-1:0] O1_I1_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv0_O1_I1_R2_C07_rom_inst (.q(O1_I1_R2_C0_SM1 ),.address(input_fmap_1[55:48]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R2_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O1_I1_R2_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O1_I1_R2_C07_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv0_O1_I1_R2_C07_rom_inst (.q(O1_I1_R2_C0_SM1 ),.address(input_fmap_1[55:48]),.clock  (clk));
logic [13-1:0] O1_I1_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv0_O1_I1_R2_C19_rom_inst (.q(O1_I1_R2_C1_SM1 ),.address(input_fmap_1[63:56]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R2_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O1_I1_R2_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O1_I1_R2_C19_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv0_O1_I1_R2_C19_rom_inst (.q(O1_I1_R2_C1_SM1 ),.address(input_fmap_1[63:56]),.clock  (clk));
logic [11-1:0] O1_I1_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O1_I1_R2_C23_rom_inst (.q(O1_I1_R2_C2_SM1 ),.address(input_fmap_1[71:64]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R2_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O1_I1_R2_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O1_I1_R2_C23_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O1_I1_R2_C23_rom_inst (.q(O1_I1_R2_C2_SM1 ),.address(input_fmap_1[71:64]),.clock  (clk));
logic [10-1:0] O1_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O1_I2_R0_C01_rom_inst (.q(O1_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O1_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O1_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O1_I2_R0_C01_rom_inst (.q(O1_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [10-1:0] O1_I2_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O1_I2_R0_C11_rom_inst (.q(O1_I2_R0_C1_SM1 ),.address(input_fmap_2[15:8]),.clk(clk),.d(0),.we(0));
//assign O1_I2_R0_C1_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O1_I2_R0_C1_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O1_I2_R0_C11_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O1_I2_R0_C11_rom_inst (.q(O1_I2_R0_C1_SM1 ),.address(input_fmap_2[15:8]),.clock  (clk));
logic [10-1:0] O1_I2_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O1_I2_R0_C21_rom_inst (.q(O1_I2_R0_C2_SM1 ),.address(input_fmap_2[23:16]),.clk(clk),.d(0),.we(0));
//assign O1_I2_R0_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O1_I2_R0_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O1_I2_R0_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O1_I2_R0_C21_rom_inst (.q(O1_I2_R0_C2_SM1 ),.address(input_fmap_2[23:16]),.clock  (clk));
logic [10-1:0] O1_I2_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O1_I2_R2_C01_rom_inst (.q(O1_I2_R2_C0_SM1 ),.address(input_fmap_2[55:48]),.clk(clk),.d(0),.we(0));
//assign O1_I2_R2_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O1_I2_R2_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O1_I2_R2_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O1_I2_R2_C01_rom_inst (.q(O1_I2_R2_C0_SM1 ),.address(input_fmap_2[55:48]),.clock  (clk));
logic [10-1:0] O1_I2_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O1_I2_R2_C11_rom_inst (.q(O1_I2_R2_C1_SM1 ),.address(input_fmap_2[63:56]),.clk(clk),.d(0),.we(0));
//assign O1_I2_R2_C1_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O1_I2_R2_C1_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O1_I2_R2_C11_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O1_I2_R2_C11_rom_inst (.q(O1_I2_R2_C1_SM1 ),.address(input_fmap_2[63:56]),.clock  (clk));
logic [10-1:0] O1_I2_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O1_I2_R2_C21_rom_inst (.q(O1_I2_R2_C2_SM1 ),.address(input_fmap_2[71:64]),.clk(clk),.d(0),.we(0));
//assign O1_I2_R2_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O1_I2_R2_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O1_I2_R2_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O1_I2_R2_C21_rom_inst (.q(O1_I2_R2_C2_SM1 ),.address(input_fmap_2[71:64]),.clock  (clk));
logic [10-1:0] O2_I0_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O2_I0_R1_C21_rom_inst (.q(O2_I0_R1_C2_SM1 ),.address(input_fmap_0[47:40]),.clk(clk),.d(0),.we(0));
//assign O2_I0_R1_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O2_I0_R1_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O2_I0_R1_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O2_I0_R1_C21_rom_inst (.q(O2_I0_R1_C2_SM1 ),.address(input_fmap_0[47:40]),.clock  (clk));
logic [10-1:0] O2_I0_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O2_I0_R2_C01_rom_inst (.q(O2_I0_R2_C0_SM1 ),.address(input_fmap_0[55:48]),.clk(clk),.d(0),.we(0));
//assign O2_I0_R2_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O2_I0_R2_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O2_I0_R2_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O2_I0_R2_C01_rom_inst (.q(O2_I0_R2_C0_SM1 ),.address(input_fmap_0[55:48]),.clock  (clk));
logic [10-1:0] O2_I0_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O2_I0_R2_C11_rom_inst (.q(O2_I0_R2_C1_SM1 ),.address(input_fmap_0[63:56]),.clk(clk),.d(0),.we(0));
//assign O2_I0_R2_C1_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O2_I0_R2_C1_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O2_I0_R2_C11_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O2_I0_R2_C11_rom_inst (.q(O2_I0_R2_C1_SM1 ),.address(input_fmap_0[63:56]),.clock  (clk));
logic [10-1:0] O2_I0_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O2_I0_R2_C21_rom_inst (.q(O2_I0_R2_C2_SM1 ),.address(input_fmap_0[71:64]),.clk(clk),.d(0),.we(0));
//assign O2_I0_R2_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O2_I0_R2_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O2_I0_R2_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O2_I0_R2_C21_rom_inst (.q(O2_I0_R2_C2_SM1 ),.address(input_fmap_0[71:64]),.clock  (clk));
logic [10-1:0] O2_I1_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O2_I1_R2_C21_rom_inst (.q(O2_I1_R2_C2_SM1 ),.address(input_fmap_1[71:64]),.clk(clk),.d(0),.we(0));
//assign O2_I1_R2_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O2_I1_R2_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O2_I1_R2_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O2_I1_R2_C21_rom_inst (.q(O2_I1_R2_C2_SM1 ),.address(input_fmap_1[71:64]),.clock  (clk));
logic [10-1:0] O2_I2_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O2_I2_R2_C21_rom_inst (.q(O2_I2_R2_C2_SM1 ),.address(input_fmap_2[71:64]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R2_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O2_I2_R2_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O2_I2_R2_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O2_I2_R2_C21_rom_inst (.q(O2_I2_R2_C2_SM1 ),.address(input_fmap_2[71:64]),.clock  (clk));
logic [14-1:0] O3_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv0_O3_I0_R0_C017_rom_inst (.q(O3_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I0_R0_C0_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O3_I0_R0_C0_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O3_I0_R0_C017_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv0_O3_I0_R0_C017_rom_inst (.q(O3_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [10-1:0] O3_I0_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O3_I0_R0_C11_rom_inst (.q(O3_I0_R0_C1_SM1 ),.address(input_fmap_0[15:8]),.clk(clk),.d(0),.we(0));
//assign O3_I0_R0_C1_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O3_I0_R0_C1_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O3_I0_R0_C11_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O3_I0_R0_C11_rom_inst (.q(O3_I0_R0_C1_SM1 ),.address(input_fmap_0[15:8]),.clock  (clk));
logic [14-1:0] O3_I0_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv0_O3_I0_R0_C222_rom_inst (.q(O3_I0_R0_C2_SM1 ),.address(input_fmap_0[23:16]),.clk(clk),.d(0),.we(0));
//assign O3_I0_R0_C2_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O3_I0_R0_C2_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O3_I0_R0_C222_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv0_O3_I0_R0_C222_rom_inst (.q(O3_I0_R0_C2_SM1 ),.address(input_fmap_0[23:16]),.clock  (clk));
logic [14-1:0] O3_I0_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv0_O3_I0_R1_C024_rom_inst (.q(O3_I0_R1_C0_SM1 ),.address(input_fmap_0[31:24]),.clk(clk),.d(0),.we(0));
//assign O3_I0_R1_C0_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O3_I0_R1_C0_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O3_I0_R1_C024_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv0_O3_I0_R1_C024_rom_inst (.q(O3_I0_R1_C0_SM1 ),.address(input_fmap_0[31:24]),.clock  (clk));
logic [10-1:0] O3_I0_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O3_I0_R1_C11_rom_inst (.q(O3_I0_R1_C1_SM1 ),.address(input_fmap_0[39:32]),.clk(clk),.d(0),.we(0));
//assign O3_I0_R1_C1_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O3_I0_R1_C1_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O3_I0_R1_C11_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O3_I0_R1_C11_rom_inst (.q(O3_I0_R1_C1_SM1 ),.address(input_fmap_0[39:32]),.clock  (clk));
logic [14-1:0] O3_I0_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv0_O3_I0_R1_C224_rom_inst (.q(O3_I0_R1_C2_SM1 ),.address(input_fmap_0[47:40]),.clk(clk),.d(0),.we(0));
//assign O3_I0_R1_C2_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O3_I0_R1_C2_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O3_I0_R1_C224_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv0_O3_I0_R1_C224_rom_inst (.q(O3_I0_R1_C2_SM1 ),.address(input_fmap_0[47:40]),.clock  (clk));
logic [13-1:0] O3_I0_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv0_O3_I0_R2_C010_rom_inst (.q(O3_I0_R2_C0_SM1 ),.address(input_fmap_0[55:48]),.clk(clk),.d(0),.we(0));
//assign O3_I0_R2_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O3_I0_R2_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O3_I0_R2_C010_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv0_O3_I0_R2_C010_rom_inst (.q(O3_I0_R2_C0_SM1 ),.address(input_fmap_0[55:48]),.clock  (clk));
logic [10-1:0] O3_I0_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O3_I0_R2_C11_rom_inst (.q(O3_I0_R2_C1_SM1 ),.address(input_fmap_0[63:56]),.clk(clk),.d(0),.we(0));
//assign O3_I0_R2_C1_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O3_I0_R2_C1_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O3_I0_R2_C11_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O3_I0_R2_C11_rom_inst (.q(O3_I0_R2_C1_SM1 ),.address(input_fmap_0[63:56]),.clock  (clk));
logic [13-1:0] O3_I0_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv0_O3_I0_R2_C210_rom_inst (.q(O3_I0_R2_C2_SM1 ),.address(input_fmap_0[71:64]),.clk(clk),.d(0),.we(0));
//assign O3_I0_R2_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O3_I0_R2_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O3_I0_R2_C210_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv0_O3_I0_R2_C210_rom_inst (.q(O3_I0_R2_C2_SM1 ),.address(input_fmap_0[71:64]),.clock  (clk));
logic [14-1:0] O3_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv0_O3_I1_R0_C020_rom_inst (.q(O3_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I1_R0_C0_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O3_I1_R0_C0_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O3_I1_R0_C020_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv0_O3_I1_R0_C020_rom_inst (.q(O3_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [10-1:0] O3_I1_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O3_I1_R0_C11_rom_inst (.q(O3_I1_R0_C1_SM1 ),.address(input_fmap_1[15:8]),.clk(clk),.d(0),.we(0));
//assign O3_I1_R0_C1_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O3_I1_R0_C1_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O3_I1_R0_C11_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O3_I1_R0_C11_rom_inst (.q(O3_I1_R0_C1_SM1 ),.address(input_fmap_1[15:8]),.clock  (clk));
logic [14-1:0] O3_I1_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv0_O3_I1_R0_C223_rom_inst (.q(O3_I1_R0_C2_SM1 ),.address(input_fmap_1[23:16]),.clk(clk),.d(0),.we(0));
//assign O3_I1_R0_C2_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O3_I1_R0_C2_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O3_I1_R0_C223_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv0_O3_I1_R0_C223_rom_inst (.q(O3_I1_R0_C2_SM1 ),.address(input_fmap_1[23:16]),.clock  (clk));
logic [14-1:0] O3_I1_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv0_O3_I1_R1_C030_rom_inst (.q(O3_I1_R1_C0_SM1 ),.address(input_fmap_1[31:24]),.clk(clk),.d(0),.we(0));
//assign O3_I1_R1_C0_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O3_I1_R1_C0_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O3_I1_R1_C030_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv0_O3_I1_R1_C030_rom_inst (.q(O3_I1_R1_C0_SM1 ),.address(input_fmap_1[31:24]),.clock  (clk));
logic [10-1:0] O3_I1_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O3_I1_R1_C11_rom_inst (.q(O3_I1_R1_C1_SM1 ),.address(input_fmap_1[39:32]),.clk(clk),.d(0),.we(0));
//assign O3_I1_R1_C1_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O3_I1_R1_C1_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O3_I1_R1_C11_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O3_I1_R1_C11_rom_inst (.q(O3_I1_R1_C1_SM1 ),.address(input_fmap_1[39:32]),.clock  (clk));
logic [14-1:0] O3_I1_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv0_O3_I1_R1_C226_rom_inst (.q(O3_I1_R1_C2_SM1 ),.address(input_fmap_1[47:40]),.clk(clk),.d(0),.we(0));
//assign O3_I1_R1_C2_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O3_I1_R1_C2_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O3_I1_R1_C226_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv0_O3_I1_R1_C226_rom_inst (.q(O3_I1_R1_C2_SM1 ),.address(input_fmap_1[47:40]),.clock  (clk));
logic [13-1:0] O3_I1_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv0_O3_I1_R2_C015_rom_inst (.q(O3_I1_R2_C0_SM1 ),.address(input_fmap_1[55:48]),.clk(clk),.d(0),.we(0));
//assign O3_I1_R2_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O3_I1_R2_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O3_I1_R2_C015_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv0_O3_I1_R2_C015_rom_inst (.q(O3_I1_R2_C0_SM1 ),.address(input_fmap_1[55:48]),.clock  (clk));
logic [10-1:0] O3_I1_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O3_I1_R2_C11_rom_inst (.q(O3_I1_R2_C1_SM1 ),.address(input_fmap_1[63:56]),.clk(clk),.d(0),.we(0));
//assign O3_I1_R2_C1_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O3_I1_R2_C1_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O3_I1_R2_C11_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O3_I1_R2_C11_rom_inst (.q(O3_I1_R2_C1_SM1 ),.address(input_fmap_1[63:56]),.clock  (clk));
logic [13-1:0] O3_I1_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv0_O3_I1_R2_C212_rom_inst (.q(O3_I1_R2_C2_SM1 ),.address(input_fmap_1[71:64]),.clk(clk),.d(0),.we(0));
//assign O3_I1_R2_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O3_I1_R2_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O3_I1_R2_C212_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv0_O3_I1_R2_C212_rom_inst (.q(O3_I1_R2_C2_SM1 ),.address(input_fmap_1[71:64]),.clock  (clk));
logic [13-1:0] O3_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv0_O3_I2_R0_C011_rom_inst (.q(O3_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I2_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O3_I2_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O3_I2_R0_C011_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv0_O3_I2_R0_C011_rom_inst (.q(O3_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [13-1:0] O3_I2_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv0_O3_I2_R0_C213_rom_inst (.q(O3_I2_R0_C2_SM1 ),.address(input_fmap_2[23:16]),.clk(clk),.d(0),.we(0));
//assign O3_I2_R0_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O3_I2_R0_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O3_I2_R0_C213_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv0_O3_I2_R0_C213_rom_inst (.q(O3_I2_R0_C2_SM1 ),.address(input_fmap_2[23:16]),.clock  (clk));
logic [13-1:0] O3_I2_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv0_O3_I2_R1_C015_rom_inst (.q(O3_I2_R1_C0_SM1 ),.address(input_fmap_2[31:24]),.clk(clk),.d(0),.we(0));
//assign O3_I2_R1_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O3_I2_R1_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O3_I2_R1_C015_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv0_O3_I2_R1_C015_rom_inst (.q(O3_I2_R1_C0_SM1 ),.address(input_fmap_2[31:24]),.clock  (clk));
logic [13-1:0] O3_I2_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv0_O3_I2_R1_C212_rom_inst (.q(O3_I2_R1_C2_SM1 ),.address(input_fmap_2[47:40]),.clk(clk),.d(0),.we(0));
//assign O3_I2_R1_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O3_I2_R1_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O3_I2_R1_C212_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv0_O3_I2_R1_C212_rom_inst (.q(O3_I2_R1_C2_SM1 ),.address(input_fmap_2[47:40]),.clock  (clk));
logic [12-1:0] O3_I2_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv0_O3_I2_R2_C04_rom_inst (.q(O3_I2_R2_C0_SM1 ),.address(input_fmap_2[55:48]),.clk(clk),.d(0),.we(0));
//assign O3_I2_R2_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O3_I2_R2_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O3_I2_R2_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv0_O3_I2_R2_C04_rom_inst (.q(O3_I2_R2_C0_SM1 ),.address(input_fmap_2[55:48]),.clock  (clk));
logic [11-1:0] O3_I2_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O3_I2_R2_C13_rom_inst (.q(O3_I2_R2_C1_SM1 ),.address(input_fmap_2[63:56]),.clk(clk),.d(0),.we(0));
//assign O3_I2_R2_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O3_I2_R2_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O3_I2_R2_C13_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O3_I2_R2_C13_rom_inst (.q(O3_I2_R2_C1_SM1 ),.address(input_fmap_2[63:56]),.clock  (clk));
logic [12-1:0] O3_I2_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv0_O3_I2_R2_C25_rom_inst (.q(O3_I2_R2_C2_SM1 ),.address(input_fmap_2[71:64]),.clk(clk),.d(0),.we(0));
//assign O3_I2_R2_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O3_I2_R2_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O3_I2_R2_C25_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv0_O3_I2_R2_C25_rom_inst (.q(O3_I2_R2_C2_SM1 ),.address(input_fmap_2[71:64]),.clock  (clk));
logic [10-1:0] O4_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O4_I0_R0_C01_rom_inst (.q(O4_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I0_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I0_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O4_I0_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O4_I0_R0_C01_rom_inst (.q(O4_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [10-1:0] O4_I0_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O4_I0_R0_C11_rom_inst (.q(O4_I0_R0_C1_SM1 ),.address(input_fmap_0[15:8]),.clk(clk),.d(0),.we(0));
//assign O4_I0_R0_C1_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I0_R0_C1_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O4_I0_R0_C11_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O4_I0_R0_C11_rom_inst (.q(O4_I0_R0_C1_SM1 ),.address(input_fmap_0[15:8]),.clock  (clk));
logic [11-1:0] O4_I0_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O4_I0_R0_C22_rom_inst (.q(O4_I0_R0_C2_SM1 ),.address(input_fmap_0[23:16]),.clk(clk),.d(0),.we(0));
//assign O4_I0_R0_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O4_I0_R0_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O4_I0_R0_C22_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O4_I0_R0_C22_rom_inst (.q(O4_I0_R0_C2_SM1 ),.address(input_fmap_0[23:16]),.clock  (clk));
logic [10-1:0] O4_I0_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O4_I0_R1_C01_rom_inst (.q(O4_I0_R1_C0_SM1 ),.address(input_fmap_0[31:24]),.clk(clk),.d(0),.we(0));
//assign O4_I0_R1_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I0_R1_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O4_I0_R1_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O4_I0_R1_C01_rom_inst (.q(O4_I0_R1_C0_SM1 ),.address(input_fmap_0[31:24]),.clock  (clk));
logic [11-1:0] O4_I0_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O4_I0_R1_C12_rom_inst (.q(O4_I0_R1_C1_SM1 ),.address(input_fmap_0[39:32]),.clk(clk),.d(0),.we(0));
//assign O4_I0_R1_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O4_I0_R1_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O4_I0_R1_C12_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O4_I0_R1_C12_rom_inst (.q(O4_I0_R1_C1_SM1 ),.address(input_fmap_0[39:32]),.clock  (clk));
logic [11-1:0] O4_I0_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O4_I0_R1_C23_rom_inst (.q(O4_I0_R1_C2_SM1 ),.address(input_fmap_0[47:40]),.clk(clk),.d(0),.we(0));
//assign O4_I0_R1_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O4_I0_R1_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O4_I0_R1_C23_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O4_I0_R1_C23_rom_inst (.q(O4_I0_R1_C2_SM1 ),.address(input_fmap_0[47:40]),.clock  (clk));
logic [10-1:0] O4_I0_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O4_I0_R2_C01_rom_inst (.q(O4_I0_R2_C0_SM1 ),.address(input_fmap_0[55:48]),.clk(clk),.d(0),.we(0));
//assign O4_I0_R2_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I0_R2_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O4_I0_R2_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O4_I0_R2_C01_rom_inst (.q(O4_I0_R2_C0_SM1 ),.address(input_fmap_0[55:48]),.clock  (clk));
logic [10-1:0] O4_I0_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O4_I0_R2_C11_rom_inst (.q(O4_I0_R2_C1_SM1 ),.address(input_fmap_0[63:56]),.clk(clk),.d(0),.we(0));
//assign O4_I0_R2_C1_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I0_R2_C1_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O4_I0_R2_C11_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O4_I0_R2_C11_rom_inst (.q(O4_I0_R2_C1_SM1 ),.address(input_fmap_0[63:56]),.clock  (clk));
logic [10-1:0] O4_I0_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O4_I0_R2_C21_rom_inst (.q(O4_I0_R2_C2_SM1 ),.address(input_fmap_0[71:64]),.clk(clk),.d(0),.we(0));
//assign O4_I0_R2_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I0_R2_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O4_I0_R2_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O4_I0_R2_C21_rom_inst (.q(O4_I0_R2_C2_SM1 ),.address(input_fmap_0[71:64]),.clock  (clk));
logic [11-1:0] O4_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O4_I1_R0_C02_rom_inst (.q(O4_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I1_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O4_I1_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O4_I1_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O4_I1_R0_C02_rom_inst (.q(O4_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [11-1:0] O4_I1_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O4_I1_R0_C22_rom_inst (.q(O4_I1_R0_C2_SM1 ),.address(input_fmap_1[23:16]),.clk(clk),.d(0),.we(0));
//assign O4_I1_R0_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O4_I1_R0_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O4_I1_R0_C22_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O4_I1_R0_C22_rom_inst (.q(O4_I1_R0_C2_SM1 ),.address(input_fmap_1[23:16]),.clock  (clk));
logic [11-1:0] O4_I1_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O4_I1_R1_C02_rom_inst (.q(O4_I1_R1_C0_SM1 ),.address(input_fmap_1[31:24]),.clk(clk),.d(0),.we(0));
//assign O4_I1_R1_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O4_I1_R1_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O4_I1_R1_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O4_I1_R1_C02_rom_inst (.q(O4_I1_R1_C0_SM1 ),.address(input_fmap_1[31:24]),.clock  (clk));
logic [11-1:0] O4_I1_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O4_I1_R1_C12_rom_inst (.q(O4_I1_R1_C1_SM1 ),.address(input_fmap_1[39:32]),.clk(clk),.d(0),.we(0));
//assign O4_I1_R1_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O4_I1_R1_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O4_I1_R1_C12_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O4_I1_R1_C12_rom_inst (.q(O4_I1_R1_C1_SM1 ),.address(input_fmap_1[39:32]),.clock  (clk));
logic [11-1:0] O4_I1_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O4_I1_R1_C23_rom_inst (.q(O4_I1_R1_C2_SM1 ),.address(input_fmap_1[47:40]),.clk(clk),.d(0),.we(0));
//assign O4_I1_R1_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O4_I1_R1_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O4_I1_R1_C23_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O4_I1_R1_C23_rom_inst (.q(O4_I1_R1_C2_SM1 ),.address(input_fmap_1[47:40]),.clock  (clk));
logic [10-1:0] O4_I1_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O4_I1_R2_C11_rom_inst (.q(O4_I1_R2_C1_SM1 ),.address(input_fmap_1[63:56]),.clk(clk),.d(0),.we(0));
//assign O4_I1_R2_C1_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I1_R2_C1_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O4_I1_R2_C11_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O4_I1_R2_C11_rom_inst (.q(O4_I1_R2_C1_SM1 ),.address(input_fmap_1[63:56]),.clock  (clk));
logic [10-1:0] O4_I1_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O4_I1_R2_C21_rom_inst (.q(O4_I1_R2_C2_SM1 ),.address(input_fmap_1[71:64]),.clk(clk),.d(0),.we(0));
//assign O4_I1_R2_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I1_R2_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O4_I1_R2_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O4_I1_R2_C21_rom_inst (.q(O4_I1_R2_C2_SM1 ),.address(input_fmap_1[71:64]),.clock  (clk));
logic [11-1:0] O4_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O4_I2_R0_C02_rom_inst (.q(O4_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I2_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O4_I2_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O4_I2_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O4_I2_R0_C02_rom_inst (.q(O4_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [10-1:0] O4_I2_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O4_I2_R0_C11_rom_inst (.q(O4_I2_R0_C1_SM1 ),.address(input_fmap_2[15:8]),.clk(clk),.d(0),.we(0));
//assign O4_I2_R0_C1_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I2_R0_C1_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O4_I2_R0_C11_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O4_I2_R0_C11_rom_inst (.q(O4_I2_R0_C1_SM1 ),.address(input_fmap_2[15:8]),.clock  (clk));
logic [11-1:0] O4_I2_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O4_I2_R1_C12_rom_inst (.q(O4_I2_R1_C1_SM1 ),.address(input_fmap_2[39:32]),.clk(clk),.d(0),.we(0));
//assign O4_I2_R1_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O4_I2_R1_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O4_I2_R1_C12_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O4_I2_R1_C12_rom_inst (.q(O4_I2_R1_C1_SM1 ),.address(input_fmap_2[39:32]),.clock  (clk));
logic [10-1:0] O4_I2_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O4_I2_R1_C21_rom_inst (.q(O4_I2_R1_C2_SM1 ),.address(input_fmap_2[47:40]),.clk(clk),.d(0),.we(0));
//assign O4_I2_R1_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I2_R1_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O4_I2_R1_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O4_I2_R1_C21_rom_inst (.q(O4_I2_R1_C2_SM1 ),.address(input_fmap_2[47:40]),.clock  (clk));
logic [10-1:0] O4_I2_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O4_I2_R2_C01_rom_inst (.q(O4_I2_R2_C0_SM1 ),.address(input_fmap_2[55:48]),.clk(clk),.d(0),.we(0));
//assign O4_I2_R2_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I2_R2_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O4_I2_R2_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O4_I2_R2_C01_rom_inst (.q(O4_I2_R2_C0_SM1 ),.address(input_fmap_2[55:48]),.clock  (clk));
logic [10-1:0] O4_I2_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O4_I2_R2_C11_rom_inst (.q(O4_I2_R2_C1_SM1 ),.address(input_fmap_2[63:56]),.clk(clk),.d(0),.we(0));
//assign O4_I2_R2_C1_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I2_R2_C1_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O4_I2_R2_C11_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O4_I2_R2_C11_rom_inst (.q(O4_I2_R2_C1_SM1 ),.address(input_fmap_2[63:56]),.clock  (clk));
logic [10-1:0] O4_I2_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O4_I2_R2_C21_rom_inst (.q(O4_I2_R2_C2_SM1 ),.address(input_fmap_2[71:64]),.clk(clk),.d(0),.we(0));
//assign O4_I2_R2_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I2_R2_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O4_I2_R2_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O4_I2_R2_C21_rom_inst (.q(O4_I2_R2_C2_SM1 ),.address(input_fmap_2[71:64]),.clock  (clk));
logic [10-1:0] O5_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O5_I0_R0_C01_rom_inst (.q(O5_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I0_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I0_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O5_I0_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O5_I0_R0_C01_rom_inst (.q(O5_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [10-1:0] O5_I0_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O5_I0_R0_C21_rom_inst (.q(O5_I0_R0_C2_SM1 ),.address(input_fmap_0[23:16]),.clk(clk),.d(0),.we(0));
//assign O5_I0_R0_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I0_R0_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O5_I0_R0_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O5_I0_R0_C21_rom_inst (.q(O5_I0_R0_C2_SM1 ),.address(input_fmap_0[23:16]),.clock  (clk));
logic [10-1:0] O5_I0_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O5_I0_R1_C01_rom_inst (.q(O5_I0_R1_C0_SM1 ),.address(input_fmap_0[31:24]),.clk(clk),.d(0),.we(0));
//assign O5_I0_R1_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I0_R1_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O5_I0_R1_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O5_I0_R1_C01_rom_inst (.q(O5_I0_R1_C0_SM1 ),.address(input_fmap_0[31:24]),.clock  (clk));
logic [11-1:0] O5_I0_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O5_I0_R1_C12_rom_inst (.q(O5_I0_R1_C1_SM1 ),.address(input_fmap_0[39:32]),.clk(clk),.d(0),.we(0));
//assign O5_I0_R1_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O5_I0_R1_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O5_I0_R1_C12_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O5_I0_R1_C12_rom_inst (.q(O5_I0_R1_C1_SM1 ),.address(input_fmap_0[39:32]),.clock  (clk));
logic [10-1:0] O5_I0_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O5_I0_R1_C21_rom_inst (.q(O5_I0_R1_C2_SM1 ),.address(input_fmap_0[47:40]),.clk(clk),.d(0),.we(0));
//assign O5_I0_R1_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I0_R1_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O5_I0_R1_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O5_I0_R1_C21_rom_inst (.q(O5_I0_R1_C2_SM1 ),.address(input_fmap_0[47:40]),.clock  (clk));
logic [10-1:0] O5_I0_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O5_I0_R2_C01_rom_inst (.q(O5_I0_R2_C0_SM1 ),.address(input_fmap_0[55:48]),.clk(clk),.d(0),.we(0));
//assign O5_I0_R2_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I0_R2_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O5_I0_R2_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O5_I0_R2_C01_rom_inst (.q(O5_I0_R2_C0_SM1 ),.address(input_fmap_0[55:48]),.clock  (clk));
logic [11-1:0] O5_I0_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O5_I0_R2_C12_rom_inst (.q(O5_I0_R2_C1_SM1 ),.address(input_fmap_0[63:56]),.clk(clk),.d(0),.we(0));
//assign O5_I0_R2_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O5_I0_R2_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O5_I0_R2_C12_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O5_I0_R2_C12_rom_inst (.q(O5_I0_R2_C1_SM1 ),.address(input_fmap_0[63:56]),.clock  (clk));
logic [10-1:0] O5_I0_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O5_I0_R2_C21_rom_inst (.q(O5_I0_R2_C2_SM1 ),.address(input_fmap_0[71:64]),.clk(clk),.d(0),.we(0));
//assign O5_I0_R2_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I0_R2_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O5_I0_R2_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O5_I0_R2_C21_rom_inst (.q(O5_I0_R2_C2_SM1 ),.address(input_fmap_0[71:64]),.clock  (clk));
logic [10-1:0] O5_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O5_I1_R0_C01_rom_inst (.q(O5_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I1_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I1_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O5_I1_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O5_I1_R0_C01_rom_inst (.q(O5_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [10-1:0] O5_I1_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O5_I1_R0_C11_rom_inst (.q(O5_I1_R0_C1_SM1 ),.address(input_fmap_1[15:8]),.clk(clk),.d(0),.we(0));
//assign O5_I1_R0_C1_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I1_R0_C1_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O5_I1_R0_C11_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O5_I1_R0_C11_rom_inst (.q(O5_I1_R0_C1_SM1 ),.address(input_fmap_1[15:8]),.clock  (clk));
logic [10-1:0] O5_I1_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O5_I1_R0_C21_rom_inst (.q(O5_I1_R0_C2_SM1 ),.address(input_fmap_1[23:16]),.clk(clk),.d(0),.we(0));
//assign O5_I1_R0_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I1_R0_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O5_I1_R0_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O5_I1_R0_C21_rom_inst (.q(O5_I1_R0_C2_SM1 ),.address(input_fmap_1[23:16]),.clock  (clk));
logic [10-1:0] O5_I1_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O5_I1_R1_C01_rom_inst (.q(O5_I1_R1_C0_SM1 ),.address(input_fmap_1[31:24]),.clk(clk),.d(0),.we(0));
//assign O5_I1_R1_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I1_R1_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O5_I1_R1_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O5_I1_R1_C01_rom_inst (.q(O5_I1_R1_C0_SM1 ),.address(input_fmap_1[31:24]),.clock  (clk));
logic [11-1:0] O5_I1_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O5_I1_R1_C12_rom_inst (.q(O5_I1_R1_C1_SM1 ),.address(input_fmap_1[39:32]),.clk(clk),.d(0),.we(0));
//assign O5_I1_R1_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O5_I1_R1_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O5_I1_R1_C12_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O5_I1_R1_C12_rom_inst (.q(O5_I1_R1_C1_SM1 ),.address(input_fmap_1[39:32]),.clock  (clk));
logic [11-1:0] O5_I1_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O5_I1_R1_C23_rom_inst (.q(O5_I1_R1_C2_SM1 ),.address(input_fmap_1[47:40]),.clk(clk),.d(0),.we(0));
//assign O5_I1_R1_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O5_I1_R1_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O5_I1_R1_C23_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O5_I1_R1_C23_rom_inst (.q(O5_I1_R1_C2_SM1 ),.address(input_fmap_1[47:40]),.clock  (clk));
logic [10-1:0] O5_I1_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O5_I1_R2_C01_rom_inst (.q(O5_I1_R2_C0_SM1 ),.address(input_fmap_1[55:48]),.clk(clk),.d(0),.we(0));
//assign O5_I1_R2_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I1_R2_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O5_I1_R2_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O5_I1_R2_C01_rom_inst (.q(O5_I1_R2_C0_SM1 ),.address(input_fmap_1[55:48]),.clock  (clk));
logic [11-1:0] O5_I1_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O5_I1_R2_C12_rom_inst (.q(O5_I1_R2_C1_SM1 ),.address(input_fmap_1[63:56]),.clk(clk),.d(0),.we(0));
//assign O5_I1_R2_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O5_I1_R2_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O5_I1_R2_C12_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O5_I1_R2_C12_rom_inst (.q(O5_I1_R2_C1_SM1 ),.address(input_fmap_1[63:56]),.clock  (clk));
logic [11-1:0] O5_I1_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O5_I1_R2_C22_rom_inst (.q(O5_I1_R2_C2_SM1 ),.address(input_fmap_1[71:64]),.clk(clk),.d(0),.we(0));
//assign O5_I1_R2_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O5_I1_R2_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O5_I1_R2_C22_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O5_I1_R2_C22_rom_inst (.q(O5_I1_R2_C2_SM1 ),.address(input_fmap_1[71:64]),.clock  (clk));
logic [10-1:0] O5_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O5_I2_R0_C01_rom_inst (.q(O5_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O5_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O5_I2_R0_C01_rom_inst (.q(O5_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [10-1:0] O5_I2_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O5_I2_R1_C01_rom_inst (.q(O5_I2_R1_C0_SM1 ),.address(input_fmap_2[31:24]),.clk(clk),.d(0),.we(0));
//assign O5_I2_R1_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I2_R1_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O5_I2_R1_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O5_I2_R1_C01_rom_inst (.q(O5_I2_R1_C0_SM1 ),.address(input_fmap_2[31:24]),.clock  (clk));
logic [10-1:0] O5_I2_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O5_I2_R1_C11_rom_inst (.q(O5_I2_R1_C1_SM1 ),.address(input_fmap_2[39:32]),.clk(clk),.d(0),.we(0));
//assign O5_I2_R1_C1_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I2_R1_C1_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O5_I2_R1_C11_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O5_I2_R1_C11_rom_inst (.q(O5_I2_R1_C1_SM1 ),.address(input_fmap_2[39:32]),.clock  (clk));
logic [10-1:0] O5_I2_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O5_I2_R1_C21_rom_inst (.q(O5_I2_R1_C2_SM1 ),.address(input_fmap_2[47:40]),.clk(clk),.d(0),.we(0));
//assign O5_I2_R1_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I2_R1_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O5_I2_R1_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O5_I2_R1_C21_rom_inst (.q(O5_I2_R1_C2_SM1 ),.address(input_fmap_2[47:40]),.clock  (clk));
logic [10-1:0] O5_I2_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O5_I2_R2_C11_rom_inst (.q(O5_I2_R2_C1_SM1 ),.address(input_fmap_2[63:56]),.clk(clk),.d(0),.we(0));
//assign O5_I2_R2_C1_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I2_R2_C1_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O5_I2_R2_C11_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O5_I2_R2_C11_rom_inst (.q(O5_I2_R2_C1_SM1 ),.address(input_fmap_2[63:56]),.clock  (clk));
logic [10-1:0] O6_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O6_I0_R0_C01_rom_inst (.q(O6_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I0_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O6_I0_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O6_I0_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O6_I0_R0_C01_rom_inst (.q(O6_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [11-1:0] O6_I0_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O6_I0_R0_C12_rom_inst (.q(O6_I0_R0_C1_SM1 ),.address(input_fmap_0[15:8]),.clk(clk),.d(0),.we(0));
//assign O6_I0_R0_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O6_I0_R0_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O6_I0_R0_C12_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O6_I0_R0_C12_rom_inst (.q(O6_I0_R0_C1_SM1 ),.address(input_fmap_0[15:8]),.clock  (clk));
logic [10-1:0] O6_I0_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O6_I0_R0_C21_rom_inst (.q(O6_I0_R0_C2_SM1 ),.address(input_fmap_0[23:16]),.clk(clk),.d(0),.we(0));
//assign O6_I0_R0_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O6_I0_R0_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O6_I0_R0_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O6_I0_R0_C21_rom_inst (.q(O6_I0_R0_C2_SM1 ),.address(input_fmap_0[23:16]),.clock  (clk));
logic [11-1:0] O6_I0_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O6_I0_R1_C02_rom_inst (.q(O6_I0_R1_C0_SM1 ),.address(input_fmap_0[31:24]),.clk(clk),.d(0),.we(0));
//assign O6_I0_R1_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O6_I0_R1_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O6_I0_R1_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O6_I0_R1_C02_rom_inst (.q(O6_I0_R1_C0_SM1 ),.address(input_fmap_0[31:24]),.clock  (clk));
logic [11-1:0] O6_I0_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O6_I0_R1_C12_rom_inst (.q(O6_I0_R1_C1_SM1 ),.address(input_fmap_0[39:32]),.clk(clk),.d(0),.we(0));
//assign O6_I0_R1_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O6_I0_R1_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O6_I0_R1_C12_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O6_I0_R1_C12_rom_inst (.q(O6_I0_R1_C1_SM1 ),.address(input_fmap_0[39:32]),.clock  (clk));
logic [10-1:0] O6_I0_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O6_I0_R1_C21_rom_inst (.q(O6_I0_R1_C2_SM1 ),.address(input_fmap_0[47:40]),.clk(clk),.d(0),.we(0));
//assign O6_I0_R1_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O6_I0_R1_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O6_I0_R1_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O6_I0_R1_C21_rom_inst (.q(O6_I0_R1_C2_SM1 ),.address(input_fmap_0[47:40]),.clock  (clk));
logic [11-1:0] O6_I0_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O6_I0_R2_C02_rom_inst (.q(O6_I0_R2_C0_SM1 ),.address(input_fmap_0[55:48]),.clk(clk),.d(0),.we(0));
//assign O6_I0_R2_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O6_I0_R2_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O6_I0_R2_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O6_I0_R2_C02_rom_inst (.q(O6_I0_R2_C0_SM1 ),.address(input_fmap_0[55:48]),.clock  (clk));
logic [11-1:0] O6_I0_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O6_I0_R2_C12_rom_inst (.q(O6_I0_R2_C1_SM1 ),.address(input_fmap_0[63:56]),.clk(clk),.d(0),.we(0));
//assign O6_I0_R2_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O6_I0_R2_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O6_I0_R2_C12_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O6_I0_R2_C12_rom_inst (.q(O6_I0_R2_C1_SM1 ),.address(input_fmap_0[63:56]),.clock  (clk));
logic [10-1:0] O6_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O6_I1_R0_C01_rom_inst (.q(O6_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I1_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O6_I1_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O6_I1_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O6_I1_R0_C01_rom_inst (.q(O6_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [10-1:0] O6_I1_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O6_I1_R0_C21_rom_inst (.q(O6_I1_R0_C2_SM1 ),.address(input_fmap_1[23:16]),.clk(clk),.d(0),.we(0));
//assign O6_I1_R0_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O6_I1_R0_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O6_I1_R0_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O6_I1_R0_C21_rom_inst (.q(O6_I1_R0_C2_SM1 ),.address(input_fmap_1[23:16]),.clock  (clk));
logic [10-1:0] O6_I1_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O6_I1_R1_C01_rom_inst (.q(O6_I1_R1_C0_SM1 ),.address(input_fmap_1[31:24]),.clk(clk),.d(0),.we(0));
//assign O6_I1_R1_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O6_I1_R1_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O6_I1_R1_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O6_I1_R1_C01_rom_inst (.q(O6_I1_R1_C0_SM1 ),.address(input_fmap_1[31:24]),.clock  (clk));
logic [10-1:0] O6_I1_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O6_I1_R1_C11_rom_inst (.q(O6_I1_R1_C1_SM1 ),.address(input_fmap_1[39:32]),.clk(clk),.d(0),.we(0));
//assign O6_I1_R1_C1_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O6_I1_R1_C1_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O6_I1_R1_C11_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O6_I1_R1_C11_rom_inst (.q(O6_I1_R1_C1_SM1 ),.address(input_fmap_1[39:32]),.clock  (clk));
logic [10-1:0] O6_I1_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O6_I1_R1_C21_rom_inst (.q(O6_I1_R1_C2_SM1 ),.address(input_fmap_1[47:40]),.clk(clk),.d(0),.we(0));
//assign O6_I1_R1_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O6_I1_R1_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O6_I1_R1_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O6_I1_R1_C21_rom_inst (.q(O6_I1_R1_C2_SM1 ),.address(input_fmap_1[47:40]),.clock  (clk));
logic [10-1:0] O6_I1_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O6_I1_R2_C01_rom_inst (.q(O6_I1_R2_C0_SM1 ),.address(input_fmap_1[55:48]),.clk(clk),.d(0),.we(0));
//assign O6_I1_R2_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O6_I1_R2_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O6_I1_R2_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O6_I1_R2_C01_rom_inst (.q(O6_I1_R2_C0_SM1 ),.address(input_fmap_1[55:48]),.clock  (clk));
logic [11-1:0] O6_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O6_I2_R0_C02_rom_inst (.q(O6_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I2_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O6_I2_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O6_I2_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O6_I2_R0_C02_rom_inst (.q(O6_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [11-1:0] O6_I2_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O6_I2_R0_C12_rom_inst (.q(O6_I2_R0_C1_SM1 ),.address(input_fmap_2[15:8]),.clk(clk),.d(0),.we(0));
//assign O6_I2_R0_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O6_I2_R0_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O6_I2_R0_C12_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O6_I2_R0_C12_rom_inst (.q(O6_I2_R0_C1_SM1 ),.address(input_fmap_2[15:8]),.clock  (clk));
logic [10-1:0] O6_I2_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O6_I2_R0_C21_rom_inst (.q(O6_I2_R0_C2_SM1 ),.address(input_fmap_2[23:16]),.clk(clk),.d(0),.we(0));
//assign O6_I2_R0_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O6_I2_R0_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O6_I2_R0_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O6_I2_R0_C21_rom_inst (.q(O6_I2_R0_C2_SM1 ),.address(input_fmap_2[23:16]),.clock  (clk));
logic [11-1:0] O6_I2_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O6_I2_R1_C03_rom_inst (.q(O6_I2_R1_C0_SM1 ),.address(input_fmap_2[31:24]),.clk(clk),.d(0),.we(0));
//assign O6_I2_R1_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O6_I2_R1_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O6_I2_R1_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O6_I2_R1_C03_rom_inst (.q(O6_I2_R1_C0_SM1 ),.address(input_fmap_2[31:24]),.clock  (clk));
logic [11-1:0] O6_I2_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O6_I2_R1_C12_rom_inst (.q(O6_I2_R1_C1_SM1 ),.address(input_fmap_2[39:32]),.clk(clk),.d(0),.we(0));
//assign O6_I2_R1_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O6_I2_R1_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O6_I2_R1_C12_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O6_I2_R1_C12_rom_inst (.q(O6_I2_R1_C1_SM1 ),.address(input_fmap_2[39:32]),.clock  (clk));
logic [10-1:0] O6_I2_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O6_I2_R1_C21_rom_inst (.q(O6_I2_R1_C2_SM1 ),.address(input_fmap_2[47:40]),.clk(clk),.d(0),.we(0));
//assign O6_I2_R1_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O6_I2_R1_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O6_I2_R1_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O6_I2_R1_C21_rom_inst (.q(O6_I2_R1_C2_SM1 ),.address(input_fmap_2[47:40]),.clock  (clk));
logic [11-1:0] O6_I2_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O6_I2_R2_C03_rom_inst (.q(O6_I2_R2_C0_SM1 ),.address(input_fmap_2[55:48]),.clk(clk),.d(0),.we(0));
//assign O6_I2_R2_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O6_I2_R2_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O6_I2_R2_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O6_I2_R2_C03_rom_inst (.q(O6_I2_R2_C0_SM1 ),.address(input_fmap_2[55:48]),.clock  (clk));
logic [11-1:0] O6_I2_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O6_I2_R2_C12_rom_inst (.q(O6_I2_R2_C1_SM1 ),.address(input_fmap_2[63:56]),.clk(clk),.d(0),.we(0));
//assign O6_I2_R2_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O6_I2_R2_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O6_I2_R2_C12_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O6_I2_R2_C12_rom_inst (.q(O6_I2_R2_C1_SM1 ),.address(input_fmap_2[63:56]),.clock  (clk));
logic [10-1:0] O6_I2_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O6_I2_R2_C21_rom_inst (.q(O6_I2_R2_C2_SM1 ),.address(input_fmap_2[71:64]),.clk(clk),.d(0),.we(0));
//assign O6_I2_R2_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O6_I2_R2_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O6_I2_R2_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O6_I2_R2_C21_rom_inst (.q(O6_I2_R2_C2_SM1 ),.address(input_fmap_2[71:64]),.clock  (clk));
logic [10-1:0] O7_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O7_I0_R0_C01_rom_inst (.q(O7_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I0_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O7_I0_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O7_I0_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O7_I0_R0_C01_rom_inst (.q(O7_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [10-1:0] O7_I0_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O7_I0_R0_C11_rom_inst (.q(O7_I0_R0_C1_SM1 ),.address(input_fmap_0[15:8]),.clk(clk),.d(0),.we(0));
//assign O7_I0_R0_C1_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O7_I0_R0_C1_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O7_I0_R0_C11_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O7_I0_R0_C11_rom_inst (.q(O7_I0_R0_C1_SM1 ),.address(input_fmap_0[15:8]),.clock  (clk));
logic [11-1:0] O7_I0_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O7_I0_R0_C22_rom_inst (.q(O7_I0_R0_C2_SM1 ),.address(input_fmap_0[23:16]),.clk(clk),.d(0),.we(0));
//assign O7_I0_R0_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O7_I0_R0_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O7_I0_R0_C22_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O7_I0_R0_C22_rom_inst (.q(O7_I0_R0_C2_SM1 ),.address(input_fmap_0[23:16]),.clock  (clk));
logic [11-1:0] O7_I0_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O7_I0_R1_C02_rom_inst (.q(O7_I0_R1_C0_SM1 ),.address(input_fmap_0[31:24]),.clk(clk),.d(0),.we(0));
//assign O7_I0_R1_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O7_I0_R1_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O7_I0_R1_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O7_I0_R1_C02_rom_inst (.q(O7_I0_R1_C0_SM1 ),.address(input_fmap_0[31:24]),.clock  (clk));
logic [11-1:0] O7_I0_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O7_I0_R1_C12_rom_inst (.q(O7_I0_R1_C1_SM1 ),.address(input_fmap_0[39:32]),.clk(clk),.d(0),.we(0));
//assign O7_I0_R1_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O7_I0_R1_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O7_I0_R1_C12_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O7_I0_R1_C12_rom_inst (.q(O7_I0_R1_C1_SM1 ),.address(input_fmap_0[39:32]),.clock  (clk));
logic [11-1:0] O7_I0_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O7_I0_R1_C22_rom_inst (.q(O7_I0_R1_C2_SM1 ),.address(input_fmap_0[47:40]),.clk(clk),.d(0),.we(0));
//assign O7_I0_R1_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O7_I0_R1_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O7_I0_R1_C22_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O7_I0_R1_C22_rom_inst (.q(O7_I0_R1_C2_SM1 ),.address(input_fmap_0[47:40]),.clock  (clk));
logic [11-1:0] O7_I0_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O7_I0_R2_C02_rom_inst (.q(O7_I0_R2_C0_SM1 ),.address(input_fmap_0[55:48]),.clk(clk),.d(0),.we(0));
//assign O7_I0_R2_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O7_I0_R2_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O7_I0_R2_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O7_I0_R2_C02_rom_inst (.q(O7_I0_R2_C0_SM1 ),.address(input_fmap_0[55:48]),.clock  (clk));
logic [11-1:0] O7_I0_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O7_I0_R2_C12_rom_inst (.q(O7_I0_R2_C1_SM1 ),.address(input_fmap_0[63:56]),.clk(clk),.d(0),.we(0));
//assign O7_I0_R2_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O7_I0_R2_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O7_I0_R2_C12_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O7_I0_R2_C12_rom_inst (.q(O7_I0_R2_C1_SM1 ),.address(input_fmap_0[63:56]),.clock  (clk));
logic [11-1:0] O7_I0_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O7_I0_R2_C22_rom_inst (.q(O7_I0_R2_C2_SM1 ),.address(input_fmap_0[71:64]),.clk(clk),.d(0),.we(0));
//assign O7_I0_R2_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O7_I0_R2_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O7_I0_R2_C22_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O7_I0_R2_C22_rom_inst (.q(O7_I0_R2_C2_SM1 ),.address(input_fmap_0[71:64]),.clock  (clk));
logic [11-1:0] O7_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O7_I1_R0_C02_rom_inst (.q(O7_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I1_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O7_I1_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O7_I1_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O7_I1_R0_C02_rom_inst (.q(O7_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [11-1:0] O7_I1_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O7_I1_R0_C12_rom_inst (.q(O7_I1_R0_C1_SM1 ),.address(input_fmap_1[15:8]),.clk(clk),.d(0),.we(0));
//assign O7_I1_R0_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O7_I1_R0_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O7_I1_R0_C12_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O7_I1_R0_C12_rom_inst (.q(O7_I1_R0_C1_SM1 ),.address(input_fmap_1[15:8]),.clock  (clk));
logic [11-1:0] O7_I1_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O7_I1_R0_C22_rom_inst (.q(O7_I1_R0_C2_SM1 ),.address(input_fmap_1[23:16]),.clk(clk),.d(0),.we(0));
//assign O7_I1_R0_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O7_I1_R0_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O7_I1_R0_C22_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O7_I1_R0_C22_rom_inst (.q(O7_I1_R0_C2_SM1 ),.address(input_fmap_1[23:16]),.clock  (clk));
logic [10-1:0] O7_I1_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O7_I1_R1_C01_rom_inst (.q(O7_I1_R1_C0_SM1 ),.address(input_fmap_1[31:24]),.clk(clk),.d(0),.we(0));
//assign O7_I1_R1_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O7_I1_R1_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O7_I1_R1_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O7_I1_R1_C01_rom_inst (.q(O7_I1_R1_C0_SM1 ),.address(input_fmap_1[31:24]),.clock  (clk));
logic [11-1:0] O7_I1_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O7_I1_R1_C12_rom_inst (.q(O7_I1_R1_C1_SM1 ),.address(input_fmap_1[39:32]),.clk(clk),.d(0),.we(0));
//assign O7_I1_R1_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O7_I1_R1_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O7_I1_R1_C12_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O7_I1_R1_C12_rom_inst (.q(O7_I1_R1_C1_SM1 ),.address(input_fmap_1[39:32]),.clock  (clk));
logic [11-1:0] O7_I1_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O7_I1_R1_C22_rom_inst (.q(O7_I1_R1_C2_SM1 ),.address(input_fmap_1[47:40]),.clk(clk),.d(0),.we(0));
//assign O7_I1_R1_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O7_I1_R1_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O7_I1_R1_C22_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O7_I1_R1_C22_rom_inst (.q(O7_I1_R1_C2_SM1 ),.address(input_fmap_1[47:40]),.clock  (clk));
logic [11-1:0] O7_I1_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O7_I1_R2_C02_rom_inst (.q(O7_I1_R2_C0_SM1 ),.address(input_fmap_1[55:48]),.clk(clk),.d(0),.we(0));
//assign O7_I1_R2_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O7_I1_R2_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O7_I1_R2_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O7_I1_R2_C02_rom_inst (.q(O7_I1_R2_C0_SM1 ),.address(input_fmap_1[55:48]),.clock  (clk));
logic [11-1:0] O7_I1_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O7_I1_R2_C12_rom_inst (.q(O7_I1_R2_C1_SM1 ),.address(input_fmap_1[63:56]),.clk(clk),.d(0),.we(0));
//assign O7_I1_R2_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O7_I1_R2_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O7_I1_R2_C12_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O7_I1_R2_C12_rom_inst (.q(O7_I1_R2_C1_SM1 ),.address(input_fmap_1[63:56]),.clock  (clk));
logic [11-1:0] O7_I1_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv0_O7_I1_R2_C22_rom_inst (.q(O7_I1_R2_C2_SM1 ),.address(input_fmap_1[71:64]),.clk(clk),.d(0),.we(0));
//assign O7_I1_R2_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O7_I1_R2_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O7_I1_R2_C22_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv0_O7_I1_R2_C22_rom_inst (.q(O7_I1_R2_C2_SM1 ),.address(input_fmap_1[71:64]),.clock  (clk));
logic [10-1:0] O7_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv0_O7_I2_R0_C01_rom_inst (.q(O7_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O7_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv0_O7_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv0_O7_I2_R0_C01_rom_inst (.q(O7_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic signed [31:0] conv_mac_0;
logic signed [31:0] O0_N0_S0;		always @(posedge clk) O0_N0_S0 <=     O0_I0_R0_C0_SM1   +  O0_I0_R0_C1_SM1  ;
 logic signed [31:0] O0_N2_S0;		always @(posedge clk) O0_N2_S0 <=     O0_I0_R0_C2_SM1   +  O0_I0_R1_C0_SM1  ;
 logic signed [31:0] O0_N4_S0;		always @(posedge clk) O0_N4_S0 <=     O0_I0_R1_C1_SM1   +  O0_I0_R1_C2_SM1  ;
 logic signed [31:0] O0_N6_S0;		always @(posedge clk) O0_N6_S0 <=     O0_I0_R2_C0_SM1   +  O0_I0_R2_C1_SM1  ;
 logic signed [31:0] O0_N8_S0;		always @(posedge clk) O0_N8_S0 <=     O0_I0_R2_C2_SM1   +  O0_I1_R0_C0_SM1  ;
 logic signed [31:0] O0_N10_S0;		always @(posedge clk) O0_N10_S0 <=     O0_I1_R0_C1_SM1   +  O0_I1_R0_C2_SM1  ;
 logic signed [31:0] O0_N12_S0;		always @(posedge clk) O0_N12_S0 <=     O0_I1_R1_C0_SM1   +  O0_I1_R1_C1_SM1  ;
 logic signed [31:0] O0_N14_S0;		always @(posedge clk) O0_N14_S0 <=     O0_I1_R1_C2_SM1   +  O0_I1_R2_C0_SM1  ;
 logic signed [31:0] O0_N16_S0;		always @(posedge clk) O0_N16_S0 <=     O0_I1_R2_C1_SM1   +  O0_I1_R2_C2_SM1  ;
 logic signed [31:0] O0_N18_S0;		always @(posedge clk) O0_N18_S0 <=     O0_I2_R0_C0_SM1   +  O0_I2_R0_C1_SM1  ;
 logic signed [31:0] O0_N20_S0;		always @(posedge clk) O0_N20_S0 <=     O0_I2_R0_C2_SM1   +  O0_I2_R1_C0_SM1  ;
 logic signed [31:0] O0_N22_S0;		always @(posedge clk) O0_N22_S0 <=     O0_I2_R1_C1_SM1   +  O0_I2_R1_C2_SM1  ;
 logic signed [31:0] O0_N24_S0;		always @(posedge clk) O0_N24_S0 <=     O0_I2_R2_C0_SM1   +  O0_I2_R2_C1_SM1  ;
 logic signed [31:0] O0_N26_S0;		always @(posedge clk) O0_N26_S0 <=     O0_I2_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O0_N0_S1;		always @(posedge clk) O0_N0_S1 <=     O0_N0_S0  +  O0_N2_S0 ;
 logic signed [31:0] O0_N2_S1;		always @(posedge clk) O0_N2_S1 <=     O0_N4_S0  +  O0_N6_S0 ;
 logic signed [31:0] O0_N4_S1;		always @(posedge clk) O0_N4_S1 <=     O0_N8_S0  +  O0_N10_S0 ;
 logic signed [31:0] O0_N6_S1;		always @(posedge clk) O0_N6_S1 <=     O0_N12_S0  +  O0_N14_S0 ;
 logic signed [31:0] O0_N8_S1;		always @(posedge clk) O0_N8_S1 <=     O0_N16_S0  +  O0_N18_S0 ;
 logic signed [31:0] O0_N10_S1;		always @(posedge clk) O0_N10_S1 <=     O0_N20_S0  +  O0_N22_S0 ;
 logic signed [31:0] O0_N12_S1;		always @(posedge clk) O0_N12_S1 <=     O0_N24_S0  +  O0_N26_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O0_N0_S2;		always @(posedge clk) O0_N0_S2 <=     O0_N0_S1  +  O0_N2_S1 ;
 logic signed [31:0] O0_N2_S2;		always @(posedge clk) O0_N2_S2 <=     O0_N4_S1  +  O0_N6_S1 ;
 logic signed [31:0] O0_N4_S2;		always @(posedge clk) O0_N4_S2 <=     O0_N8_S1  +  O0_N10_S1 ;
 logic signed [31:0] O0_N6_S2;		always @(posedge clk) O0_N6_S2 <=     O0_N12_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O0_N0_S3;		always @(posedge clk) O0_N0_S3 <=     O0_N0_S2  +  O0_N2_S2 ;
 logic signed [31:0] O0_N2_S3;		always @(posedge clk) O0_N2_S3 <=     O0_N4_S2  +  O0_N6_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O0_N0_S4;		always @(posedge clk) O0_N0_S4 <=     O0_N0_S3  +  O0_N2_S3 ;
 assign conv_mac_0 = O0_N0_S4;

logic signed [31:0] conv_mac_1;
logic signed [31:0] O1_N0_S0;		always @(posedge clk) O1_N0_S0 <=     O1_I0_R0_C0_SM1   +  O1_I0_R0_C1_SM1  ;
 logic signed [31:0] O1_N2_S0;		always @(posedge clk) O1_N2_S0 <=     O1_I0_R0_C2_SM1   +  O1_I0_R1_C0_SM1  ;
 logic signed [31:0] O1_N4_S0;		always @(posedge clk) O1_N4_S0 <=     O1_I0_R1_C1_SM1   +  O1_I0_R1_C2_SM1  ;
 logic signed [31:0] O1_N6_S0;		always @(posedge clk) O1_N6_S0 <=     O1_I0_R2_C0_SM1   +  O1_I0_R2_C1_SM1  ;
 logic signed [31:0] O1_N8_S0;		always @(posedge clk) O1_N8_S0 <=     O1_I0_R2_C2_SM1   +  O1_I1_R0_C0_SM1  ;
 logic signed [31:0] O1_N10_S0;		always @(posedge clk) O1_N10_S0 <=     O1_I1_R0_C1_SM1   +  O1_I1_R0_C2_SM1  ;
 logic signed [31:0] O1_N12_S0;		always @(posedge clk) O1_N12_S0 <=     O1_I1_R1_C0_SM1   +  O1_I1_R1_C1_SM1  ;
 logic signed [31:0] O1_N14_S0;		always @(posedge clk) O1_N14_S0 <=     O1_I1_R1_C2_SM1   +  O1_I1_R2_C0_SM1  ;
 logic signed [31:0] O1_N16_S0;		always @(posedge clk) O1_N16_S0 <=     O1_I1_R2_C1_SM1   +  O1_I1_R2_C2_SM1  ;
 logic signed [31:0] O1_N18_S0;		always @(posedge clk) O1_N18_S0 <=     O1_I2_R0_C0_SM1   +  O1_I2_R0_C1_SM1  ;
 logic signed [31:0] O1_N20_S0;		always @(posedge clk) O1_N20_S0 <=     O1_I2_R0_C2_SM1   +  O1_I2_R2_C0_SM1  ;
 logic signed [31:0] O1_N22_S0;		always @(posedge clk) O1_N22_S0 <=     O1_I2_R2_C1_SM1   +  O1_I2_R2_C2_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O1_N0_S1;		always @(posedge clk) O1_N0_S1 <=     O1_N0_S0  +  O1_N2_S0 ;
 logic signed [31:0] O1_N2_S1;		always @(posedge clk) O1_N2_S1 <=     O1_N4_S0  +  O1_N6_S0 ;
 logic signed [31:0] O1_N4_S1;		always @(posedge clk) O1_N4_S1 <=     O1_N8_S0  +  O1_N10_S0 ;
 logic signed [31:0] O1_N6_S1;		always @(posedge clk) O1_N6_S1 <=     O1_N12_S0  +  O1_N14_S0 ;
 logic signed [31:0] O1_N8_S1;		always @(posedge clk) O1_N8_S1 <=     O1_N16_S0  +  O1_N18_S0 ;
 logic signed [31:0] O1_N10_S1;		always @(posedge clk) O1_N10_S1 <=     O1_N20_S0  +  O1_N22_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O1_N0_S2;		always @(posedge clk) O1_N0_S2 <=     O1_N0_S1  +  O1_N2_S1 ;
 logic signed [31:0] O1_N2_S2;		always @(posedge clk) O1_N2_S2 <=     O1_N4_S1  +  O1_N6_S1 ;
 logic signed [31:0] O1_N4_S2;		always @(posedge clk) O1_N4_S2 <=     O1_N8_S1  +  O1_N10_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O1_N0_S3;		always @(posedge clk) O1_N0_S3 <=     O1_N0_S2  +  O1_N2_S2 ;
 logic signed [31:0] O1_N2_S3;		always @(posedge clk) O1_N2_S3 <=     O1_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O1_N0_S4;		always @(posedge clk) O1_N0_S4 <=     O1_N0_S3  +  O1_N2_S3 ;
 assign conv_mac_1 = O1_N0_S4;

logic signed [31:0] conv_mac_2;
logic signed [31:0] O2_N0_S0;		always @(posedge clk) O2_N0_S0 <=     O2_I0_R1_C2_SM1   +  O2_I0_R2_C0_SM1  ;
 logic signed [31:0] O2_N2_S0;		always @(posedge clk) O2_N2_S0 <=     O2_I0_R2_C1_SM1   +  O2_I0_R2_C2_SM1  ;
 logic signed [31:0] O2_N4_S0;		always @(posedge clk) O2_N4_S0 <=     O2_I1_R2_C2_SM1   +  O2_I2_R2_C2_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O2_N0_S1;		always @(posedge clk) O2_N0_S1 <=     O2_N0_S0  +  O2_N2_S0 ;
 logic signed [31:0] O2_N2_S1;		always @(posedge clk) O2_N2_S1 <=     O2_N4_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O2_N0_S2;		always @(posedge clk) O2_N0_S2 <=     O2_N0_S1  +  O2_N2_S1 ;
 assign conv_mac_2 = O2_N0_S2;

logic signed [31:0] conv_mac_3;
logic signed [31:0] O3_N0_S0;		always @(posedge clk) O3_N0_S0 <=     O3_I0_R0_C0_SM1   +  O3_I0_R0_C1_SM1  ;
 logic signed [31:0] O3_N2_S0;		always @(posedge clk) O3_N2_S0 <=     O3_I0_R0_C2_SM1   +  O3_I0_R1_C0_SM1  ;
 logic signed [31:0] O3_N4_S0;		always @(posedge clk) O3_N4_S0 <=     O3_I0_R1_C1_SM1   +  O3_I0_R1_C2_SM1  ;
 logic signed [31:0] O3_N6_S0;		always @(posedge clk) O3_N6_S0 <=     O3_I0_R2_C0_SM1   +  O3_I0_R2_C1_SM1  ;
 logic signed [31:0] O3_N8_S0;		always @(posedge clk) O3_N8_S0 <=     O3_I0_R2_C2_SM1   +  O3_I1_R0_C0_SM1  ;
 logic signed [31:0] O3_N10_S0;		always @(posedge clk) O3_N10_S0 <=     O3_I1_R0_C1_SM1   +  O3_I1_R0_C2_SM1  ;
 logic signed [31:0] O3_N12_S0;		always @(posedge clk) O3_N12_S0 <=     O3_I1_R1_C0_SM1   +  O3_I1_R1_C1_SM1  ;
 logic signed [31:0] O3_N14_S0;		always @(posedge clk) O3_N14_S0 <=     O3_I1_R1_C2_SM1   +  O3_I1_R2_C0_SM1  ;
 logic signed [31:0] O3_N16_S0;		always @(posedge clk) O3_N16_S0 <=     O3_I1_R2_C1_SM1   +  O3_I1_R2_C2_SM1  ;
 logic signed [31:0] O3_N18_S0;		always @(posedge clk) O3_N18_S0 <=     O3_I2_R0_C0_SM1   +  O3_I2_R0_C2_SM1  ;
 logic signed [31:0] O3_N20_S0;		always @(posedge clk) O3_N20_S0 <=     O3_I2_R1_C0_SM1   +  O3_I2_R1_C2_SM1  ;
 logic signed [31:0] O3_N22_S0;		always @(posedge clk) O3_N22_S0 <=     O3_I2_R2_C0_SM1   +  O3_I2_R2_C1_SM1  ;
 logic signed [31:0] O3_N24_S0;		always @(posedge clk) O3_N24_S0 <=     O3_I2_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O3_N0_S1;		always @(posedge clk) O3_N0_S1 <=     O3_N0_S0  +  O3_N2_S0 ;
 logic signed [31:0] O3_N2_S1;		always @(posedge clk) O3_N2_S1 <=     O3_N4_S0  +  O3_N6_S0 ;
 logic signed [31:0] O3_N4_S1;		always @(posedge clk) O3_N4_S1 <=     O3_N8_S0  +  O3_N10_S0 ;
 logic signed [31:0] O3_N6_S1;		always @(posedge clk) O3_N6_S1 <=     O3_N12_S0  +  O3_N14_S0 ;
 logic signed [31:0] O3_N8_S1;		always @(posedge clk) O3_N8_S1 <=     O3_N16_S0  +  O3_N18_S0 ;
 logic signed [31:0] O3_N10_S1;		always @(posedge clk) O3_N10_S1 <=     O3_N20_S0  +  O3_N22_S0 ;
 logic signed [31:0] O3_N12_S1;		always @(posedge clk) O3_N12_S1 <=     O3_N24_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O3_N0_S2;		always @(posedge clk) O3_N0_S2 <=     O3_N0_S1  +  O3_N2_S1 ;
 logic signed [31:0] O3_N2_S2;		always @(posedge clk) O3_N2_S2 <=     O3_N4_S1  +  O3_N6_S1 ;
 logic signed [31:0] O3_N4_S2;		always @(posedge clk) O3_N4_S2 <=     O3_N8_S1  +  O3_N10_S1 ;
 logic signed [31:0] O3_N6_S2;		always @(posedge clk) O3_N6_S2 <=     O3_N12_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O3_N0_S3;		always @(posedge clk) O3_N0_S3 <=     O3_N0_S2  +  O3_N2_S2 ;
 logic signed [31:0] O3_N2_S3;		always @(posedge clk) O3_N2_S3 <=     O3_N4_S2  +  O3_N6_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O3_N0_S4;		always @(posedge clk) O3_N0_S4 <=     O3_N0_S3  +  O3_N2_S3 ;
 assign conv_mac_3 = O3_N0_S4;

logic signed [31:0] conv_mac_4;
logic signed [31:0] O4_N0_S0;		always @(posedge clk) O4_N0_S0 <=     O4_I0_R0_C0_SM1   +  O4_I0_R0_C1_SM1  ;
 logic signed [31:0] O4_N2_S0;		always @(posedge clk) O4_N2_S0 <=     O4_I0_R0_C2_SM1   +  O4_I0_R1_C0_SM1  ;
 logic signed [31:0] O4_N4_S0;		always @(posedge clk) O4_N4_S0 <=     O4_I0_R1_C1_SM1   +  O4_I0_R1_C2_SM1  ;
 logic signed [31:0] O4_N6_S0;		always @(posedge clk) O4_N6_S0 <=     O4_I0_R2_C0_SM1   +  O4_I0_R2_C1_SM1  ;
 logic signed [31:0] O4_N8_S0;		always @(posedge clk) O4_N8_S0 <=     O4_I0_R2_C2_SM1   +  O4_I1_R0_C0_SM1  ;
 logic signed [31:0] O4_N10_S0;		always @(posedge clk) O4_N10_S0 <=     O4_I1_R0_C2_SM1   +  O4_I1_R1_C0_SM1  ;
 logic signed [31:0] O4_N12_S0;		always @(posedge clk) O4_N12_S0 <=     O4_I1_R1_C1_SM1   +  O4_I1_R1_C2_SM1  ;
 logic signed [31:0] O4_N14_S0;		always @(posedge clk) O4_N14_S0 <=     O4_I1_R2_C1_SM1   +  O4_I1_R2_C2_SM1  ;
 logic signed [31:0] O4_N16_S0;		always @(posedge clk) O4_N16_S0 <=     O4_I2_R0_C0_SM1   +  O4_I2_R0_C1_SM1  ;
 logic signed [31:0] O4_N18_S0;		always @(posedge clk) O4_N18_S0 <=     O4_I2_R1_C1_SM1   +  O4_I2_R1_C2_SM1  ;
 logic signed [31:0] O4_N20_S0;		always @(posedge clk) O4_N20_S0 <=     O4_I2_R2_C0_SM1   +  O4_I2_R2_C1_SM1  ;
 logic signed [31:0] O4_N22_S0;		always @(posedge clk) O4_N22_S0 <=     O4_I2_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O4_N0_S1;		always @(posedge clk) O4_N0_S1 <=     O4_N0_S0  +  O4_N2_S0 ;
 logic signed [31:0] O4_N2_S1;		always @(posedge clk) O4_N2_S1 <=     O4_N4_S0  +  O4_N6_S0 ;
 logic signed [31:0] O4_N4_S1;		always @(posedge clk) O4_N4_S1 <=     O4_N8_S0  +  O4_N10_S0 ;
 logic signed [31:0] O4_N6_S1;		always @(posedge clk) O4_N6_S1 <=     O4_N12_S0  +  O4_N14_S0 ;
 logic signed [31:0] O4_N8_S1;		always @(posedge clk) O4_N8_S1 <=     O4_N16_S0  +  O4_N18_S0 ;
 logic signed [31:0] O4_N10_S1;		always @(posedge clk) O4_N10_S1 <=     O4_N20_S0  +  O4_N22_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O4_N0_S2;		always @(posedge clk) O4_N0_S2 <=     O4_N0_S1  +  O4_N2_S1 ;
 logic signed [31:0] O4_N2_S2;		always @(posedge clk) O4_N2_S2 <=     O4_N4_S1  +  O4_N6_S1 ;
 logic signed [31:0] O4_N4_S2;		always @(posedge clk) O4_N4_S2 <=     O4_N8_S1  +  O4_N10_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O4_N0_S3;		always @(posedge clk) O4_N0_S3 <=     O4_N0_S2  +  O4_N2_S2 ;
 logic signed [31:0] O4_N2_S3;		always @(posedge clk) O4_N2_S3 <=     O4_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O4_N0_S4;		always @(posedge clk) O4_N0_S4 <=     O4_N0_S3  +  O4_N2_S3 ;
 assign conv_mac_4 = O4_N0_S4;

logic signed [31:0] conv_mac_5;
logic signed [31:0] O5_N0_S0;		always @(posedge clk) O5_N0_S0 <=     O5_I0_R0_C0_SM1   +  O5_I0_R0_C2_SM1  ;
 logic signed [31:0] O5_N2_S0;		always @(posedge clk) O5_N2_S0 <=     O5_I0_R1_C0_SM1   +  O5_I0_R1_C1_SM1  ;
 logic signed [31:0] O5_N4_S0;		always @(posedge clk) O5_N4_S0 <=     O5_I0_R1_C2_SM1   +  O5_I0_R2_C0_SM1  ;
 logic signed [31:0] O5_N6_S0;		always @(posedge clk) O5_N6_S0 <=     O5_I0_R2_C1_SM1   +  O5_I0_R2_C2_SM1  ;
 logic signed [31:0] O5_N8_S0;		always @(posedge clk) O5_N8_S0 <=     O5_I1_R0_C0_SM1   +  O5_I1_R0_C1_SM1  ;
 logic signed [31:0] O5_N10_S0;		always @(posedge clk) O5_N10_S0 <=     O5_I1_R0_C2_SM1   +  O5_I1_R1_C0_SM1  ;
 logic signed [31:0] O5_N12_S0;		always @(posedge clk) O5_N12_S0 <=     O5_I1_R1_C1_SM1   +  O5_I1_R1_C2_SM1  ;
 logic signed [31:0] O5_N14_S0;		always @(posedge clk) O5_N14_S0 <=     O5_I1_R2_C0_SM1   +  O5_I1_R2_C1_SM1  ;
 logic signed [31:0] O5_N16_S0;		always @(posedge clk) O5_N16_S0 <=     O5_I1_R2_C2_SM1   +  O5_I2_R0_C0_SM1  ;
 logic signed [31:0] O5_N18_S0;		always @(posedge clk) O5_N18_S0 <=     O5_I2_R1_C0_SM1   +  O5_I2_R1_C1_SM1  ;
 logic signed [31:0] O5_N20_S0;		always @(posedge clk) O5_N20_S0 <=     O5_I2_R1_C2_SM1   +  O5_I2_R2_C1_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O5_N0_S1;		always @(posedge clk) O5_N0_S1 <=     O5_N0_S0  +  O5_N2_S0 ;
 logic signed [31:0] O5_N2_S1;		always @(posedge clk) O5_N2_S1 <=     O5_N4_S0  +  O5_N6_S0 ;
 logic signed [31:0] O5_N4_S1;		always @(posedge clk) O5_N4_S1 <=     O5_N8_S0  +  O5_N10_S0 ;
 logic signed [31:0] O5_N6_S1;		always @(posedge clk) O5_N6_S1 <=     O5_N12_S0  +  O5_N14_S0 ;
 logic signed [31:0] O5_N8_S1;		always @(posedge clk) O5_N8_S1 <=     O5_N16_S0  +  O5_N18_S0 ;
 logic signed [31:0] O5_N10_S1;		always @(posedge clk) O5_N10_S1 <=     O5_N20_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O5_N0_S2;		always @(posedge clk) O5_N0_S2 <=     O5_N0_S1  +  O5_N2_S1 ;
 logic signed [31:0] O5_N2_S2;		always @(posedge clk) O5_N2_S2 <=     O5_N4_S1  +  O5_N6_S1 ;
 logic signed [31:0] O5_N4_S2;		always @(posedge clk) O5_N4_S2 <=     O5_N8_S1  +  O5_N10_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O5_N0_S3;		always @(posedge clk) O5_N0_S3 <=     O5_N0_S2  +  O5_N2_S2 ;
 logic signed [31:0] O5_N2_S3;		always @(posedge clk) O5_N2_S3 <=     O5_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O5_N0_S4;		always @(posedge clk) O5_N0_S4 <=     O5_N0_S3  +  O5_N2_S3 ;
 assign conv_mac_5 = O5_N0_S4;

logic signed [31:0] conv_mac_6;
logic signed [31:0] O6_N0_S0;		always @(posedge clk) O6_N0_S0 <=     O6_I0_R0_C0_SM1   +  O6_I0_R0_C1_SM1  ;
 logic signed [31:0] O6_N2_S0;		always @(posedge clk) O6_N2_S0 <=     O6_I0_R0_C2_SM1   +  O6_I0_R1_C0_SM1  ;
 logic signed [31:0] O6_N4_S0;		always @(posedge clk) O6_N4_S0 <=     O6_I0_R1_C1_SM1   +  O6_I0_R1_C2_SM1  ;
 logic signed [31:0] O6_N6_S0;		always @(posedge clk) O6_N6_S0 <=     O6_I0_R2_C0_SM1   +  O6_I0_R2_C1_SM1  ;
 logic signed [31:0] O6_N8_S0;		always @(posedge clk) O6_N8_S0 <=     O6_I1_R0_C0_SM1   +  O6_I1_R0_C2_SM1  ;
 logic signed [31:0] O6_N10_S0;		always @(posedge clk) O6_N10_S0 <=     O6_I1_R1_C0_SM1   +  O6_I1_R1_C1_SM1  ;
 logic signed [31:0] O6_N12_S0;		always @(posedge clk) O6_N12_S0 <=     O6_I1_R1_C2_SM1   +  O6_I1_R2_C0_SM1  ;
 logic signed [31:0] O6_N14_S0;		always @(posedge clk) O6_N14_S0 <=     O6_I2_R0_C0_SM1   +  O6_I2_R0_C1_SM1  ;
 logic signed [31:0] O6_N16_S0;		always @(posedge clk) O6_N16_S0 <=     O6_I2_R0_C2_SM1   +  O6_I2_R1_C0_SM1  ;
 logic signed [31:0] O6_N18_S0;		always @(posedge clk) O6_N18_S0 <=     O6_I2_R1_C1_SM1   +  O6_I2_R1_C2_SM1  ;
 logic signed [31:0] O6_N20_S0;		always @(posedge clk) O6_N20_S0 <=     O6_I2_R2_C0_SM1   +  O6_I2_R2_C1_SM1  ;
 logic signed [31:0] O6_N22_S0;		always @(posedge clk) O6_N22_S0 <=     O6_I2_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O6_N0_S1;		always @(posedge clk) O6_N0_S1 <=     O6_N0_S0  +  O6_N2_S0 ;
 logic signed [31:0] O6_N2_S1;		always @(posedge clk) O6_N2_S1 <=     O6_N4_S0  +  O6_N6_S0 ;
 logic signed [31:0] O6_N4_S1;		always @(posedge clk) O6_N4_S1 <=     O6_N8_S0  +  O6_N10_S0 ;
 logic signed [31:0] O6_N6_S1;		always @(posedge clk) O6_N6_S1 <=     O6_N12_S0  +  O6_N14_S0 ;
 logic signed [31:0] O6_N8_S1;		always @(posedge clk) O6_N8_S1 <=     O6_N16_S0  +  O6_N18_S0 ;
 logic signed [31:0] O6_N10_S1;		always @(posedge clk) O6_N10_S1 <=     O6_N20_S0  +  O6_N22_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O6_N0_S2;		always @(posedge clk) O6_N0_S2 <=     O6_N0_S1  +  O6_N2_S1 ;
 logic signed [31:0] O6_N2_S2;		always @(posedge clk) O6_N2_S2 <=     O6_N4_S1  +  O6_N6_S1 ;
 logic signed [31:0] O6_N4_S2;		always @(posedge clk) O6_N4_S2 <=     O6_N8_S1  +  O6_N10_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O6_N0_S3;		always @(posedge clk) O6_N0_S3 <=     O6_N0_S2  +  O6_N2_S2 ;
 logic signed [31:0] O6_N2_S3;		always @(posedge clk) O6_N2_S3 <=     O6_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O6_N0_S4;		always @(posedge clk) O6_N0_S4 <=     O6_N0_S3  +  O6_N2_S3 ;
 assign conv_mac_6 = O6_N0_S4;

logic signed [31:0] conv_mac_7;
logic signed [31:0] O7_N0_S0;		always @(posedge clk) O7_N0_S0 <=     O7_I0_R0_C0_SM1   +  O7_I0_R0_C1_SM1  ;
 logic signed [31:0] O7_N2_S0;		always @(posedge clk) O7_N2_S0 <=     O7_I0_R0_C2_SM1   +  O7_I0_R1_C0_SM1  ;
 logic signed [31:0] O7_N4_S0;		always @(posedge clk) O7_N4_S0 <=     O7_I0_R1_C1_SM1   +  O7_I0_R1_C2_SM1  ;
 logic signed [31:0] O7_N6_S0;		always @(posedge clk) O7_N6_S0 <=     O7_I0_R2_C0_SM1   +  O7_I0_R2_C1_SM1  ;
 logic signed [31:0] O7_N8_S0;		always @(posedge clk) O7_N8_S0 <=     O7_I0_R2_C2_SM1   +  O7_I1_R0_C0_SM1  ;
 logic signed [31:0] O7_N10_S0;		always @(posedge clk) O7_N10_S0 <=     O7_I1_R0_C1_SM1   +  O7_I1_R0_C2_SM1  ;
 logic signed [31:0] O7_N12_S0;		always @(posedge clk) O7_N12_S0 <=     O7_I1_R1_C0_SM1   +  O7_I1_R1_C1_SM1  ;
 logic signed [31:0] O7_N14_S0;		always @(posedge clk) O7_N14_S0 <=     O7_I1_R1_C2_SM1   +  O7_I1_R2_C0_SM1  ;
 logic signed [31:0] O7_N16_S0;		always @(posedge clk) O7_N16_S0 <=     O7_I1_R2_C1_SM1   +  O7_I1_R2_C2_SM1  ;
 logic signed [31:0] O7_N18_S0;		always @(posedge clk) O7_N18_S0 <=     O7_I2_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O7_N0_S1;		always @(posedge clk) O7_N0_S1 <=     O7_N0_S0  +  O7_N2_S0 ;
 logic signed [31:0] O7_N2_S1;		always @(posedge clk) O7_N2_S1 <=     O7_N4_S0  +  O7_N6_S0 ;
 logic signed [31:0] O7_N4_S1;		always @(posedge clk) O7_N4_S1 <=     O7_N8_S0  +  O7_N10_S0 ;
 logic signed [31:0] O7_N6_S1;		always @(posedge clk) O7_N6_S1 <=     O7_N12_S0  +  O7_N14_S0 ;
 logic signed [31:0] O7_N8_S1;		always @(posedge clk) O7_N8_S1 <=     O7_N16_S0  +  O7_N18_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O7_N0_S2;		always @(posedge clk) O7_N0_S2 <=     O7_N0_S1  +  O7_N2_S1 ;
 logic signed [31:0] O7_N2_S2;		always @(posedge clk) O7_N2_S2 <=     O7_N4_S1  +  O7_N6_S1 ;
 logic signed [31:0] O7_N4_S2;		always @(posedge clk) O7_N4_S2 <=     O7_N8_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O7_N0_S3;		always @(posedge clk) O7_N0_S3 <=     O7_N0_S2  +  O7_N2_S2 ;
 logic signed [31:0] O7_N2_S3;		always @(posedge clk) O7_N2_S3 <=     O7_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O7_N0_S4;		always @(posedge clk) O7_N0_S4 <=     O7_N0_S3  +  O7_N2_S3 ;
 assign conv_mac_7 = O7_N0_S4;

logic valid_D1;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D1<= 0 ;
	else valid_D1<=valid;
end
logic valid_D2;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D2<= 0 ;
	else valid_D2<=valid_D1;
end
logic valid_D3;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D3<= 0 ;
	else valid_D3<=valid_D2;
end
logic valid_D4;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D4<= 0 ;
	else valid_D4<=valid_D3;
end
logic valid_D5;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D5<= 0 ;
	else valid_D5<=valid_D4;
end
logic valid_D6;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D6<= 0 ;
	else valid_D6<=valid_D5;
end
always_ff @(posedge clk) begin
	if (rstn == 0) ready <= 0 ;
	else ready <=valid_D6;
end
logic [31:0] bias_add_0;
assign bias_add_0 = conv_mac_0 + 7'd35;
logic [31:0] bias_add_1;
assign bias_add_1 = conv_mac_1 + 6'd30;
logic [31:0] bias_add_2;
assign bias_add_2 = conv_mac_2 + 6'd17;
logic [31:0] bias_add_3;
assign bias_add_3 = conv_mac_3 + 6'd17;
logic [31:0] bias_add_4;
assign bias_add_4 = conv_mac_4 - 5'd13;
logic [31:0] bias_add_5;
assign bias_add_5 = conv_mac_5 + 6'd31;
logic [31:0] bias_add_6;
assign bias_add_6 = conv_mac_6 + 5'd14;
logic [31:0] bias_add_7;
assign bias_add_7 = conv_mac_7 + 7'd32;

logic [7:0] relu_0;
assign relu_0[7:0] = (bias_add_0[31]==0) ? ((bias_add_0<3'd6) ? {{bias_add_0[31],bias_add_0[10:4]}} :'d6) : '0;
logic [7:0] relu_1;
assign relu_1[7:0] = (bias_add_1[31]==0) ? ((bias_add_1<3'd6) ? {{bias_add_1[31],bias_add_1[10:4]}} :'d6) : '0;
logic [7:0] relu_2;
assign relu_2[7:0] = (bias_add_2[31]==0) ? ((bias_add_2<3'd6) ? {{bias_add_2[31],bias_add_2[10:4]}} :'d6) : '0;
logic [7:0] relu_3;
assign relu_3[7:0] = (bias_add_3[31]==0) ? ((bias_add_3<3'd6) ? {{bias_add_3[31],bias_add_3[10:4]}} :'d6) : '0;
logic [7:0] relu_4;
assign relu_4[7:0] = (bias_add_4[31]==0) ? ((bias_add_4<3'd6) ? {{bias_add_4[31],bias_add_4[10:4]}} :'d6) : '0;
logic [7:0] relu_5;
assign relu_5[7:0] = (bias_add_5[31]==0) ? ((bias_add_5<3'd6) ? {{bias_add_5[31],bias_add_5[10:4]}} :'d6) : '0;
logic [7:0] relu_6;
assign relu_6[7:0] = (bias_add_6[31]==0) ? ((bias_add_6<3'd6) ? {{bias_add_6[31],bias_add_6[10:4]}} :'d6) : '0;
logic [7:0] relu_7;
assign relu_7[7:0] = (bias_add_7[31]==0) ? ((bias_add_7<3'd6) ? {{bias_add_7[31],bias_add_7[10:4]}} :'d6) : '0;

assign output_act = {
	relu_7,
	relu_6,
	relu_5,
	relu_4,
	relu_3,
	relu_2,
	relu_1,
	relu_0
};

endmodule
module conv1_dw (
    input logic clk,
    input logic rstn,
    input logic valid,
    input logic [8*72-1:0] input_act,
    output logic [64-1:0] output_act,
    output logic ready
);
logic we;
logic [8:0] zero_number; 
assign zero_number = 9'd0; 
logic [8*72-1:0] input_act_ff;
genvar i;
generate
for (i=0;i<8;i++)
    begin: genblk_6
        always_ff @(posedge clk) begin
            if (rstn == 0) begin
                input_act_ff[(i+1)*72-1:i*72] <= '0;
            end
            else begin
                input_act_ff[(i+1)*72-1:i*72] <= input_act[(i+1)*72-1:i*72];
            end
        end
    end
endgenerate
logic [71:0] input_fmap_0;
assign input_fmap_0 = input_act_ff[71:0];
logic [71:0] input_fmap_1;
assign input_fmap_1 = input_act_ff[143:72];
logic [71:0] input_fmap_2;
assign input_fmap_2 = input_act_ff[215:144];
logic [71:0] input_fmap_3;
assign input_fmap_3 = input_act_ff[287:216];
logic [71:0] input_fmap_4;
assign input_fmap_4 = input_act_ff[359:288];
logic [71:0] input_fmap_5;
assign input_fmap_5 = input_act_ff[431:360];
logic [71:0] input_fmap_6;
assign input_fmap_6 = input_act_ff[503:432];
logic [71:0] input_fmap_7;
assign input_fmap_7 = input_act_ff[575:504];

logic [14-1:0] O0_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv1_dw_O0_I0_R0_C019_rom_inst (.q(O0_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R0_C0_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O0_I0_R0_C0_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O0_I0_R0_C019_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv1_dw_O0_I0_R0_C019_rom_inst (.q(O0_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [15-1:0] O0_I0_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(15),.INIT_FILE("deepfreeze_rom/deepfreeze_8_15.txt"))
    conv1_dw_O0_I0_R0_C151_rom_inst (.q(O0_I0_R0_C1_SM1 ),.address(input_fmap_0[15:8]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R0_C1_SM1  = 15'h1234;
//always@(posedge clk) begin 
//O0_I0_R0_C1_SM1  <= 15'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O0_I0_R0_C151_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(15))
//    conv1_dw_O0_I0_R0_C151_rom_inst (.q(O0_I0_R0_C1_SM1 ),.address(input_fmap_0[15:8]),.clock  (clk));
logic [14-1:0] O0_I0_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv1_dw_O0_I0_R0_C219_rom_inst (.q(O0_I0_R0_C2_SM1 ),.address(input_fmap_0[23:16]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R0_C2_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O0_I0_R0_C2_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O0_I0_R0_C219_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv1_dw_O0_I0_R0_C219_rom_inst (.q(O0_I0_R0_C2_SM1 ),.address(input_fmap_0[23:16]),.clock  (clk));
logic [13-1:0] O0_I0_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv1_dw_O0_I0_R1_C010_rom_inst (.q(O0_I0_R1_C0_SM1 ),.address(input_fmap_0[31:24]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R1_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O0_I0_R1_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O0_I0_R1_C010_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv1_dw_O0_I0_R1_C010_rom_inst (.q(O0_I0_R1_C0_SM1 ),.address(input_fmap_0[31:24]),.clock  (clk));
logic [12-1:0] O0_I0_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv1_dw_O0_I0_R1_C15_rom_inst (.q(O0_I0_R1_C1_SM1 ),.address(input_fmap_0[39:32]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R1_C1_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O0_I0_R1_C1_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O0_I0_R1_C15_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv1_dw_O0_I0_R1_C15_rom_inst (.q(O0_I0_R1_C1_SM1 ),.address(input_fmap_0[39:32]),.clock  (clk));
logic [13-1:0] O0_I0_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv1_dw_O0_I0_R1_C28_rom_inst (.q(O0_I0_R1_C2_SM1 ),.address(input_fmap_0[47:40]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R1_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O0_I0_R1_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O0_I0_R1_C28_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv1_dw_O0_I0_R1_C28_rom_inst (.q(O0_I0_R1_C2_SM1 ),.address(input_fmap_0[47:40]),.clock  (clk));
logic [14-1:0] O0_I0_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv1_dw_O0_I0_R2_C019_rom_inst (.q(O0_I0_R2_C0_SM1 ),.address(input_fmap_0[55:48]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R2_C0_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O0_I0_R2_C0_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O0_I0_R2_C019_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv1_dw_O0_I0_R2_C019_rom_inst (.q(O0_I0_R2_C0_SM1 ),.address(input_fmap_0[55:48]),.clock  (clk));
logic [14-1:0] O0_I0_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv1_dw_O0_I0_R2_C123_rom_inst (.q(O0_I0_R2_C1_SM1 ),.address(input_fmap_0[63:56]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R2_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O0_I0_R2_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O0_I0_R2_C123_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv1_dw_O0_I0_R2_C123_rom_inst (.q(O0_I0_R2_C1_SM1 ),.address(input_fmap_0[63:56]),.clock  (clk));
logic [14-1:0] O0_I0_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv1_dw_O0_I0_R2_C219_rom_inst (.q(O0_I0_R2_C2_SM1 ),.address(input_fmap_0[71:64]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R2_C2_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O0_I0_R2_C2_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O0_I0_R2_C219_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv1_dw_O0_I0_R2_C219_rom_inst (.q(O0_I0_R2_C2_SM1 ),.address(input_fmap_0[71:64]),.clock  (clk));
logic [13-1:0] O1_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv1_dw_O1_I1_R0_C013_rom_inst (.q(O1_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O1_I1_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O1_I1_R0_C013_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv1_dw_O1_I1_R0_C013_rom_inst (.q(O1_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [16-1:0] O1_I1_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(16),.INIT_FILE("deepfreeze_rom/deepfreeze_8_16.txt"))
    conv1_dw_O1_I1_R0_C169_rom_inst (.q(O1_I1_R0_C1_SM1 ),.address(input_fmap_1[15:8]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R0_C1_SM1  = 16'h1234;
//always@(posedge clk) begin 
//O1_I1_R0_C1_SM1  <= 16'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O1_I1_R0_C169_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(16))
//    conv1_dw_O1_I1_R0_C169_rom_inst (.q(O1_I1_R0_C1_SM1 ),.address(input_fmap_1[15:8]),.clock  (clk));
logic [13-1:0] O1_I1_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv1_dw_O1_I1_R1_C08_rom_inst (.q(O1_I1_R1_C0_SM1 ),.address(input_fmap_1[31:24]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R1_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O1_I1_R1_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O1_I1_R1_C08_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv1_dw_O1_I1_R1_C08_rom_inst (.q(O1_I1_R1_C0_SM1 ),.address(input_fmap_1[31:24]),.clock  (clk));
logic [16-1:0] O1_I1_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(16),.INIT_FILE("deepfreeze_rom/deepfreeze_8_16.txt"))
    conv1_dw_O1_I1_R1_C174_rom_inst (.q(O1_I1_R1_C1_SM1 ),.address(input_fmap_1[39:32]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R1_C1_SM1  = 16'h1234;
//always@(posedge clk) begin 
//O1_I1_R1_C1_SM1  <= 16'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O1_I1_R1_C174_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(16))
//    conv1_dw_O1_I1_R1_C174_rom_inst (.q(O1_I1_R1_C1_SM1 ),.address(input_fmap_1[39:32]),.clock  (clk));
logic [12-1:0] O1_I1_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv1_dw_O1_I1_R1_C24_rom_inst (.q(O1_I1_R1_C2_SM1 ),.address(input_fmap_1[47:40]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R1_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O1_I1_R1_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O1_I1_R1_C24_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv1_dw_O1_I1_R1_C24_rom_inst (.q(O1_I1_R1_C2_SM1 ),.address(input_fmap_1[47:40]),.clock  (clk));
logic [12-1:0] O1_I1_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv1_dw_O1_I1_R2_C06_rom_inst (.q(O1_I1_R2_C0_SM1 ),.address(input_fmap_1[55:48]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R2_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O1_I1_R2_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O1_I1_R2_C06_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv1_dw_O1_I1_R2_C06_rom_inst (.q(O1_I1_R2_C0_SM1 ),.address(input_fmap_1[55:48]),.clock  (clk));
logic [12-1:0] O1_I1_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv1_dw_O1_I1_R2_C17_rom_inst (.q(O1_I1_R2_C1_SM1 ),.address(input_fmap_1[63:56]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R2_C1_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O1_I1_R2_C1_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O1_I1_R2_C17_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv1_dw_O1_I1_R2_C17_rom_inst (.q(O1_I1_R2_C1_SM1 ),.address(input_fmap_1[63:56]),.clock  (clk));
logic [12-1:0] O1_I1_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv1_dw_O1_I1_R2_C25_rom_inst (.q(O1_I1_R2_C2_SM1 ),.address(input_fmap_1[71:64]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R2_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O1_I1_R2_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O1_I1_R2_C25_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv1_dw_O1_I1_R2_C25_rom_inst (.q(O1_I1_R2_C2_SM1 ),.address(input_fmap_1[71:64]),.clock  (clk));
logic [12-1:0] O2_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv1_dw_O2_I2_R0_C05_rom_inst (.q(O2_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O2_I2_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O2_I2_R0_C05_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv1_dw_O2_I2_R0_C05_rom_inst (.q(O2_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [13-1:0] O2_I2_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv1_dw_O2_I2_R0_C19_rom_inst (.q(O2_I2_R0_C1_SM1 ),.address(input_fmap_2[15:8]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R0_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O2_I2_R0_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O2_I2_R0_C19_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv1_dw_O2_I2_R0_C19_rom_inst (.q(O2_I2_R0_C1_SM1 ),.address(input_fmap_2[15:8]),.clock  (clk));
logic [13-1:0] O2_I2_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv1_dw_O2_I2_R0_C28_rom_inst (.q(O2_I2_R0_C2_SM1 ),.address(input_fmap_2[23:16]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R0_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O2_I2_R0_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O2_I2_R0_C28_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv1_dw_O2_I2_R0_C28_rom_inst (.q(O2_I2_R0_C2_SM1 ),.address(input_fmap_2[23:16]),.clock  (clk));
logic [11-1:0] O2_I2_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv1_dw_O2_I2_R1_C03_rom_inst (.q(O2_I2_R1_C0_SM1 ),.address(input_fmap_2[31:24]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R1_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O2_I2_R1_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O2_I2_R1_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv1_dw_O2_I2_R1_C03_rom_inst (.q(O2_I2_R1_C0_SM1 ),.address(input_fmap_2[31:24]),.clock  (clk));
logic [11-1:0] O2_I2_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv1_dw_O2_I2_R1_C12_rom_inst (.q(O2_I2_R1_C1_SM1 ),.address(input_fmap_2[39:32]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R1_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O2_I2_R1_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O2_I2_R1_C12_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv1_dw_O2_I2_R1_C12_rom_inst (.q(O2_I2_R1_C1_SM1 ),.address(input_fmap_2[39:32]),.clock  (clk));
logic [12-1:0] O2_I2_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv1_dw_O2_I2_R1_C27_rom_inst (.q(O2_I2_R1_C2_SM1 ),.address(input_fmap_2[47:40]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R1_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O2_I2_R1_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O2_I2_R1_C27_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv1_dw_O2_I2_R1_C27_rom_inst (.q(O2_I2_R1_C2_SM1 ),.address(input_fmap_2[47:40]),.clock  (clk));
logic [14-1:0] O2_I2_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv1_dw_O2_I2_R2_C017_rom_inst (.q(O2_I2_R2_C0_SM1 ),.address(input_fmap_2[55:48]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R2_C0_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O2_I2_R2_C0_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O2_I2_R2_C017_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv1_dw_O2_I2_R2_C017_rom_inst (.q(O2_I2_R2_C0_SM1 ),.address(input_fmap_2[55:48]),.clock  (clk));
logic [13-1:0] O2_I2_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv1_dw_O2_I2_R2_C114_rom_inst (.q(O2_I2_R2_C1_SM1 ),.address(input_fmap_2[63:56]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R2_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O2_I2_R2_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O2_I2_R2_C114_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv1_dw_O2_I2_R2_C114_rom_inst (.q(O2_I2_R2_C1_SM1 ),.address(input_fmap_2[63:56]),.clock  (clk));
logic [11-1:0] O2_I2_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv1_dw_O2_I2_R2_C23_rom_inst (.q(O2_I2_R2_C2_SM1 ),.address(input_fmap_2[71:64]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R2_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O2_I2_R2_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O2_I2_R2_C23_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv1_dw_O2_I2_R2_C23_rom_inst (.q(O2_I2_R2_C2_SM1 ),.address(input_fmap_2[71:64]),.clock  (clk));
logic [14-1:0] O3_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv1_dw_O3_I3_R0_C031_rom_inst (.q(O3_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R0_C0_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O3_I3_R0_C0_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O3_I3_R0_C031_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv1_dw_O3_I3_R0_C031_rom_inst (.q(O3_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [11-1:0] O3_I3_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv1_dw_O3_I3_R0_C13_rom_inst (.q(O3_I3_R0_C1_SM1 ),.address(input_fmap_3[15:8]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R0_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O3_I3_R0_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O3_I3_R0_C13_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv1_dw_O3_I3_R0_C13_rom_inst (.q(O3_I3_R0_C1_SM1 ),.address(input_fmap_3[15:8]),.clock  (clk));
logic [15-1:0] O3_I3_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(15),.INIT_FILE("deepfreeze_rom/deepfreeze_8_15.txt"))
    conv1_dw_O3_I3_R0_C235_rom_inst (.q(O3_I3_R0_C2_SM1 ),.address(input_fmap_3[23:16]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R0_C2_SM1  = 15'h1234;
//always@(posedge clk) begin 
//O3_I3_R0_C2_SM1  <= 15'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O3_I3_R0_C235_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(15))
//    conv1_dw_O3_I3_R0_C235_rom_inst (.q(O3_I3_R0_C2_SM1 ),.address(input_fmap_3[23:16]),.clock  (clk));
logic [14-1:0] O3_I3_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv1_dw_O3_I3_R1_C016_rom_inst (.q(O3_I3_R1_C0_SM1 ),.address(input_fmap_3[31:24]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R1_C0_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O3_I3_R1_C0_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O3_I3_R1_C016_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv1_dw_O3_I3_R1_C016_rom_inst (.q(O3_I3_R1_C0_SM1 ),.address(input_fmap_3[31:24]),.clock  (clk));
logic [12-1:0] O3_I3_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv1_dw_O3_I3_R1_C16_rom_inst (.q(O3_I3_R1_C1_SM1 ),.address(input_fmap_3[39:32]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R1_C1_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O3_I3_R1_C1_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O3_I3_R1_C16_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv1_dw_O3_I3_R1_C16_rom_inst (.q(O3_I3_R1_C1_SM1 ),.address(input_fmap_3[39:32]),.clock  (clk));
logic [14-1:0] O3_I3_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv1_dw_O3_I3_R1_C231_rom_inst (.q(O3_I3_R1_C2_SM1 ),.address(input_fmap_3[47:40]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R1_C2_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O3_I3_R1_C2_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O3_I3_R1_C231_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv1_dw_O3_I3_R1_C231_rom_inst (.q(O3_I3_R1_C2_SM1 ),.address(input_fmap_3[47:40]),.clock  (clk));
logic [12-1:0] O3_I3_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv1_dw_O3_I3_R2_C04_rom_inst (.q(O3_I3_R2_C0_SM1 ),.address(input_fmap_3[55:48]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R2_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O3_I3_R2_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O3_I3_R2_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv1_dw_O3_I3_R2_C04_rom_inst (.q(O3_I3_R2_C0_SM1 ),.address(input_fmap_3[55:48]),.clock  (clk));
logic [13-1:0] O3_I3_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv1_dw_O3_I3_R2_C18_rom_inst (.q(O3_I3_R2_C1_SM1 ),.address(input_fmap_3[63:56]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R2_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O3_I3_R2_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O3_I3_R2_C18_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv1_dw_O3_I3_R2_C18_rom_inst (.q(O3_I3_R2_C1_SM1 ),.address(input_fmap_3[63:56]),.clock  (clk));
logic [13-1:0] O3_I3_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv1_dw_O3_I3_R2_C211_rom_inst (.q(O3_I3_R2_C2_SM1 ),.address(input_fmap_3[71:64]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R2_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O3_I3_R2_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O3_I3_R2_C211_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv1_dw_O3_I3_R2_C211_rom_inst (.q(O3_I3_R2_C2_SM1 ),.address(input_fmap_3[71:64]),.clock  (clk));
logic [11-1:0] O4_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv1_dw_O4_I4_R0_C02_rom_inst (.q(O4_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O4_I4_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O4_I4_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv1_dw_O4_I4_R0_C02_rom_inst (.q(O4_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [10-1:0] O4_I4_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv1_dw_O4_I4_R0_C11_rom_inst (.q(O4_I4_R0_C1_SM1 ),.address(input_fmap_4[15:8]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R0_C1_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I4_R0_C1_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O4_I4_R0_C11_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv1_dw_O4_I4_R0_C11_rom_inst (.q(O4_I4_R0_C1_SM1 ),.address(input_fmap_4[15:8]),.clock  (clk));
logic [14-1:0] O4_I4_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv1_dw_O4_I4_R0_C219_rom_inst (.q(O4_I4_R0_C2_SM1 ),.address(input_fmap_4[23:16]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R0_C2_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O4_I4_R0_C2_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O4_I4_R0_C219_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv1_dw_O4_I4_R0_C219_rom_inst (.q(O4_I4_R0_C2_SM1 ),.address(input_fmap_4[23:16]),.clock  (clk));
logic [13-1:0] O4_I4_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv1_dw_O4_I4_R1_C08_rom_inst (.q(O4_I4_R1_C0_SM1 ),.address(input_fmap_4[31:24]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R1_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O4_I4_R1_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O4_I4_R1_C08_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv1_dw_O4_I4_R1_C08_rom_inst (.q(O4_I4_R1_C0_SM1 ),.address(input_fmap_4[31:24]),.clock  (clk));
logic [13-1:0] O4_I4_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv1_dw_O4_I4_R1_C18_rom_inst (.q(O4_I4_R1_C1_SM1 ),.address(input_fmap_4[39:32]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R1_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O4_I4_R1_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O4_I4_R1_C18_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv1_dw_O4_I4_R1_C18_rom_inst (.q(O4_I4_R1_C1_SM1 ),.address(input_fmap_4[39:32]),.clock  (clk));
logic [12-1:0] O4_I4_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv1_dw_O4_I4_R1_C27_rom_inst (.q(O4_I4_R1_C2_SM1 ),.address(input_fmap_4[47:40]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R1_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O4_I4_R1_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O4_I4_R1_C27_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv1_dw_O4_I4_R1_C27_rom_inst (.q(O4_I4_R1_C2_SM1 ),.address(input_fmap_4[47:40]),.clock  (clk));
logic [12-1:0] O4_I4_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv1_dw_O4_I4_R2_C06_rom_inst (.q(O4_I4_R2_C0_SM1 ),.address(input_fmap_4[55:48]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R2_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O4_I4_R2_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O4_I4_R2_C06_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv1_dw_O4_I4_R2_C06_rom_inst (.q(O4_I4_R2_C0_SM1 ),.address(input_fmap_4[55:48]),.clock  (clk));
logic [12-1:0] O4_I4_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv1_dw_O4_I4_R2_C14_rom_inst (.q(O4_I4_R2_C1_SM1 ),.address(input_fmap_4[63:56]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R2_C1_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O4_I4_R2_C1_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O4_I4_R2_C14_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv1_dw_O4_I4_R2_C14_rom_inst (.q(O4_I4_R2_C1_SM1 ),.address(input_fmap_4[63:56]),.clock  (clk));
logic [12-1:0] O4_I4_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv1_dw_O4_I4_R2_C25_rom_inst (.q(O4_I4_R2_C2_SM1 ),.address(input_fmap_4[71:64]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R2_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O4_I4_R2_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O4_I4_R2_C25_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv1_dw_O4_I4_R2_C25_rom_inst (.q(O4_I4_R2_C2_SM1 ),.address(input_fmap_4[71:64]),.clock  (clk));
logic [12-1:0] O5_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv1_dw_O5_I5_R0_C04_rom_inst (.q(O5_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O5_I5_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O5_I5_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv1_dw_O5_I5_R0_C04_rom_inst (.q(O5_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [16-1:0] O5_I5_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(16),.INIT_FILE("deepfreeze_rom/deepfreeze_8_16.txt"))
    conv1_dw_O5_I5_R0_C166_rom_inst (.q(O5_I5_R0_C1_SM1 ),.address(input_fmap_5[15:8]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R0_C1_SM1  = 16'h1234;
//always@(posedge clk) begin 
//O5_I5_R0_C1_SM1  <= 16'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O5_I5_R0_C166_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(16))
//    conv1_dw_O5_I5_R0_C166_rom_inst (.q(O5_I5_R0_C1_SM1 ),.address(input_fmap_5[15:8]),.clock  (clk));
logic [15-1:0] O5_I5_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(15),.INIT_FILE("deepfreeze_rom/deepfreeze_8_15.txt"))
    conv1_dw_O5_I5_R0_C237_rom_inst (.q(O5_I5_R0_C2_SM1 ),.address(input_fmap_5[23:16]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R0_C2_SM1  = 15'h1234;
//always@(posedge clk) begin 
//O5_I5_R0_C2_SM1  <= 15'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O5_I5_R0_C237_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(15))
//    conv1_dw_O5_I5_R0_C237_rom_inst (.q(O5_I5_R0_C2_SM1 ),.address(input_fmap_5[23:16]),.clock  (clk));
logic [13-1:0] O5_I5_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv1_dw_O5_I5_R1_C09_rom_inst (.q(O5_I5_R1_C0_SM1 ),.address(input_fmap_5[31:24]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R1_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O5_I5_R1_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O5_I5_R1_C09_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv1_dw_O5_I5_R1_C09_rom_inst (.q(O5_I5_R1_C0_SM1 ),.address(input_fmap_5[31:24]),.clock  (clk));
logic [15-1:0] O5_I5_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(15),.INIT_FILE("deepfreeze_rom/deepfreeze_8_15.txt"))
    conv1_dw_O5_I5_R1_C145_rom_inst (.q(O5_I5_R1_C1_SM1 ),.address(input_fmap_5[39:32]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R1_C1_SM1  = 15'h1234;
//always@(posedge clk) begin 
//O5_I5_R1_C1_SM1  <= 15'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O5_I5_R1_C145_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(15))
//    conv1_dw_O5_I5_R1_C145_rom_inst (.q(O5_I5_R1_C1_SM1 ),.address(input_fmap_5[39:32]),.clock  (clk));
logic [12-1:0] O5_I5_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv1_dw_O5_I5_R1_C25_rom_inst (.q(O5_I5_R1_C2_SM1 ),.address(input_fmap_5[47:40]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R1_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O5_I5_R1_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O5_I5_R1_C25_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv1_dw_O5_I5_R1_C25_rom_inst (.q(O5_I5_R1_C2_SM1 ),.address(input_fmap_5[47:40]),.clock  (clk));
logic [14-1:0] O5_I5_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv1_dw_O5_I5_R2_C020_rom_inst (.q(O5_I5_R2_C0_SM1 ),.address(input_fmap_5[55:48]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R2_C0_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O5_I5_R2_C0_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O5_I5_R2_C020_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv1_dw_O5_I5_R2_C020_rom_inst (.q(O5_I5_R2_C0_SM1 ),.address(input_fmap_5[55:48]),.clock  (clk));
logic [15-1:0] O5_I5_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(15),.INIT_FILE("deepfreeze_rom/deepfreeze_8_15.txt"))
    conv1_dw_O5_I5_R2_C136_rom_inst (.q(O5_I5_R2_C1_SM1 ),.address(input_fmap_5[63:56]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R2_C1_SM1  = 15'h1234;
//always@(posedge clk) begin 
//O5_I5_R2_C1_SM1  <= 15'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O5_I5_R2_C136_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(15))
//    conv1_dw_O5_I5_R2_C136_rom_inst (.q(O5_I5_R2_C1_SM1 ),.address(input_fmap_5[63:56]),.clock  (clk));
logic [12-1:0] O5_I5_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv1_dw_O5_I5_R2_C25_rom_inst (.q(O5_I5_R2_C2_SM1 ),.address(input_fmap_5[71:64]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R2_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O5_I5_R2_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O5_I5_R2_C25_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv1_dw_O5_I5_R2_C25_rom_inst (.q(O5_I5_R2_C2_SM1 ),.address(input_fmap_5[71:64]),.clock  (clk));
logic [15-1:0] O6_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(15),.INIT_FILE("deepfreeze_rom/deepfreeze_8_15.txt"))
    conv1_dw_O6_I6_R0_C035_rom_inst (.q(O6_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R0_C0_SM1  = 15'h1234;
//always@(posedge clk) begin 
//O6_I6_R0_C0_SM1  <= 15'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O6_I6_R0_C035_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(15))
//    conv1_dw_O6_I6_R0_C035_rom_inst (.q(O6_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [14-1:0] O6_I6_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv1_dw_O6_I6_R0_C131_rom_inst (.q(O6_I6_R0_C1_SM1 ),.address(input_fmap_6[15:8]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R0_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O6_I6_R0_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O6_I6_R0_C131_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv1_dw_O6_I6_R0_C131_rom_inst (.q(O6_I6_R0_C1_SM1 ),.address(input_fmap_6[15:8]),.clock  (clk));
logic [15-1:0] O6_I6_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(15),.INIT_FILE("deepfreeze_rom/deepfreeze_8_15.txt"))
    conv1_dw_O6_I6_R0_C250_rom_inst (.q(O6_I6_R0_C2_SM1 ),.address(input_fmap_6[23:16]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R0_C2_SM1  = 15'h1234;
//always@(posedge clk) begin 
//O6_I6_R0_C2_SM1  <= 15'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O6_I6_R0_C250_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(15))
//    conv1_dw_O6_I6_R0_C250_rom_inst (.q(O6_I6_R0_C2_SM1 ),.address(input_fmap_6[23:16]),.clock  (clk));
logic [10-1:0] O6_I6_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv1_dw_O6_I6_R1_C01_rom_inst (.q(O6_I6_R1_C0_SM1 ),.address(input_fmap_6[31:24]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R1_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O6_I6_R1_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O6_I6_R1_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv1_dw_O6_I6_R1_C01_rom_inst (.q(O6_I6_R1_C0_SM1 ),.address(input_fmap_6[31:24]),.clock  (clk));
logic [14-1:0] O6_I6_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv1_dw_O6_I6_R1_C127_rom_inst (.q(O6_I6_R1_C1_SM1 ),.address(input_fmap_6[39:32]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R1_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O6_I6_R1_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O6_I6_R1_C127_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv1_dw_O6_I6_R1_C127_rom_inst (.q(O6_I6_R1_C1_SM1 ),.address(input_fmap_6[39:32]),.clock  (clk));
logic [13-1:0] O6_I6_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv1_dw_O6_I6_R1_C213_rom_inst (.q(O6_I6_R1_C2_SM1 ),.address(input_fmap_6[47:40]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R1_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O6_I6_R1_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O6_I6_R1_C213_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv1_dw_O6_I6_R1_C213_rom_inst (.q(O6_I6_R1_C2_SM1 ),.address(input_fmap_6[47:40]),.clock  (clk));
logic [11-1:0] O6_I6_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv1_dw_O6_I6_R2_C02_rom_inst (.q(O6_I6_R2_C0_SM1 ),.address(input_fmap_6[55:48]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R2_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O6_I6_R2_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O6_I6_R2_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv1_dw_O6_I6_R2_C02_rom_inst (.q(O6_I6_R2_C0_SM1 ),.address(input_fmap_6[55:48]),.clock  (clk));
logic [14-1:0] O6_I6_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv1_dw_O6_I6_R2_C129_rom_inst (.q(O6_I6_R2_C1_SM1 ),.address(input_fmap_6[63:56]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R2_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O6_I6_R2_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O6_I6_R2_C129_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv1_dw_O6_I6_R2_C129_rom_inst (.q(O6_I6_R2_C1_SM1 ),.address(input_fmap_6[63:56]),.clock  (clk));
logic [15-1:0] O6_I6_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(15),.INIT_FILE("deepfreeze_rom/deepfreeze_8_15.txt"))
    conv1_dw_O6_I6_R2_C243_rom_inst (.q(O6_I6_R2_C2_SM1 ),.address(input_fmap_6[71:64]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R2_C2_SM1  = 15'h1234;
//always@(posedge clk) begin 
//O6_I6_R2_C2_SM1  <= 15'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O6_I6_R2_C243_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(15))
//    conv1_dw_O6_I6_R2_C243_rom_inst (.q(O6_I6_R2_C2_SM1 ),.address(input_fmap_6[71:64]),.clock  (clk));
logic [12-1:0] O7_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv1_dw_O7_I7_R0_C06_rom_inst (.q(O7_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O7_I7_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O7_I7_R0_C06_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv1_dw_O7_I7_R0_C06_rom_inst (.q(O7_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [14-1:0] O7_I7_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv1_dw_O7_I7_R0_C131_rom_inst (.q(O7_I7_R0_C1_SM1 ),.address(input_fmap_7[15:8]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R0_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O7_I7_R0_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O7_I7_R0_C131_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv1_dw_O7_I7_R0_C131_rom_inst (.q(O7_I7_R0_C1_SM1 ),.address(input_fmap_7[15:8]),.clock  (clk));
logic [14-1:0] O7_I7_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv1_dw_O7_I7_R0_C230_rom_inst (.q(O7_I7_R0_C2_SM1 ),.address(input_fmap_7[23:16]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R0_C2_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O7_I7_R0_C2_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O7_I7_R0_C230_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv1_dw_O7_I7_R0_C230_rom_inst (.q(O7_I7_R0_C2_SM1 ),.address(input_fmap_7[23:16]),.clock  (clk));
logic [12-1:0] O7_I7_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv1_dw_O7_I7_R1_C06_rom_inst (.q(O7_I7_R1_C0_SM1 ),.address(input_fmap_7[31:24]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R1_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O7_I7_R1_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O7_I7_R1_C06_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv1_dw_O7_I7_R1_C06_rom_inst (.q(O7_I7_R1_C0_SM1 ),.address(input_fmap_7[31:24]),.clock  (clk));
logic [13-1:0] O7_I7_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv1_dw_O7_I7_R1_C113_rom_inst (.q(O7_I7_R1_C1_SM1 ),.address(input_fmap_7[39:32]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R1_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O7_I7_R1_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O7_I7_R1_C113_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv1_dw_O7_I7_R1_C113_rom_inst (.q(O7_I7_R1_C1_SM1 ),.address(input_fmap_7[39:32]),.clock  (clk));
logic [13-1:0] O7_I7_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv1_dw_O7_I7_R1_C212_rom_inst (.q(O7_I7_R1_C2_SM1 ),.address(input_fmap_7[47:40]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R1_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O7_I7_R1_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O7_I7_R1_C212_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv1_dw_O7_I7_R1_C212_rom_inst (.q(O7_I7_R1_C2_SM1 ),.address(input_fmap_7[47:40]),.clock  (clk));
logic [12-1:0] O7_I7_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv1_dw_O7_I7_R2_C04_rom_inst (.q(O7_I7_R2_C0_SM1 ),.address(input_fmap_7[55:48]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R2_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O7_I7_R2_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O7_I7_R2_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv1_dw_O7_I7_R2_C04_rom_inst (.q(O7_I7_R2_C0_SM1 ),.address(input_fmap_7[55:48]),.clock  (clk));
logic [15-1:0] O7_I7_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(15),.INIT_FILE("deepfreeze_rom/deepfreeze_8_15.txt"))
    conv1_dw_O7_I7_R2_C134_rom_inst (.q(O7_I7_R2_C1_SM1 ),.address(input_fmap_7[63:56]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R2_C1_SM1  = 15'h1234;
//always@(posedge clk) begin 
//O7_I7_R2_C1_SM1  <= 15'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O7_I7_R2_C134_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(15))
//    conv1_dw_O7_I7_R2_C134_rom_inst (.q(O7_I7_R2_C1_SM1 ),.address(input_fmap_7[63:56]),.clock  (clk));
logic [14-1:0] O7_I7_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv1_dw_O7_I7_R2_C224_rom_inst (.q(O7_I7_R2_C2_SM1 ),.address(input_fmap_7[71:64]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R2_C2_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O7_I7_R2_C2_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_dw_O7_I7_R2_C224_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv1_dw_O7_I7_R2_C224_rom_inst (.q(O7_I7_R2_C2_SM1 ),.address(input_fmap_7[71:64]),.clock  (clk));
logic signed [31:0] conv_mac_0;
logic signed [31:0] O0_N0_S0;		always @(posedge clk) O0_N0_S0 <=     O0_I0_R0_C0_SM1   +  O0_I0_R0_C1_SM1  ;
 logic signed [31:0] O0_N2_S0;		always @(posedge clk) O0_N2_S0 <=     O0_I0_R0_C2_SM1   +  O0_I0_R1_C0_SM1  ;
 logic signed [31:0] O0_N4_S0;		always @(posedge clk) O0_N4_S0 <=     O0_I0_R1_C1_SM1   +  O0_I0_R1_C2_SM1  ;
 logic signed [31:0] O0_N6_S0;		always @(posedge clk) O0_N6_S0 <=     O0_I0_R2_C0_SM1   +  O0_I0_R2_C1_SM1  ;
 logic signed [31:0] O0_N8_S0;		always @(posedge clk) O0_N8_S0 <=     O0_I0_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O0_N0_S1;		always @(posedge clk) O0_N0_S1 <=     O0_N0_S0  +  O0_N2_S0 ;
 logic signed [31:0] O0_N2_S1;		always @(posedge clk) O0_N2_S1 <=     O0_N4_S0  +  O0_N6_S0 ;
 logic signed [31:0] O0_N4_S1;		always @(posedge clk) O0_N4_S1 <=     O0_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O0_N0_S2;		always @(posedge clk) O0_N0_S2 <=     O0_N0_S1  +  O0_N2_S1 ;
 logic signed [31:0] O0_N2_S2;		always @(posedge clk) O0_N2_S2 <=     O0_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O0_N0_S3;		always @(posedge clk) O0_N0_S3 <=     O0_N0_S2  +  O0_N2_S2 ;
 assign conv_mac_0 = O0_N0_S3;

logic signed [31:0] conv_mac_1;
logic signed [31:0] O1_N0_S0;		always @(posedge clk) O1_N0_S0 <=     O1_I1_R0_C0_SM1   +  O1_I1_R0_C1_SM1  ;
 logic signed [31:0] O1_N2_S0;		always @(posedge clk) O1_N2_S0 <=     O1_I1_R1_C0_SM1   +  O1_I1_R1_C1_SM1  ;
 logic signed [31:0] O1_N4_S0;		always @(posedge clk) O1_N4_S0 <=     O1_I1_R1_C2_SM1   +  O1_I1_R2_C0_SM1  ;
 logic signed [31:0] O1_N6_S0;		always @(posedge clk) O1_N6_S0 <=     O1_I1_R2_C1_SM1   +  O1_I1_R2_C2_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O1_N0_S1;		always @(posedge clk) O1_N0_S1 <=     O1_N0_S0  +  O1_N2_S0 ;
 logic signed [31:0] O1_N2_S1;		always @(posedge clk) O1_N2_S1 <=     O1_N4_S0  +  O1_N6_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O1_N0_S2;		always @(posedge clk) O1_N0_S2 <=     O1_N0_S1  +  O1_N2_S1 ;
 assign conv_mac_1 = O1_N0_S2;

logic signed [31:0] conv_mac_2;
logic signed [31:0] O2_N0_S0;		always @(posedge clk) O2_N0_S0 <=     O2_I2_R0_C0_SM1   +  O2_I2_R0_C1_SM1  ;
 logic signed [31:0] O2_N2_S0;		always @(posedge clk) O2_N2_S0 <=     O2_I2_R0_C2_SM1   +  O2_I2_R1_C0_SM1  ;
 logic signed [31:0] O2_N4_S0;		always @(posedge clk) O2_N4_S0 <=     O2_I2_R1_C1_SM1   +  O2_I2_R1_C2_SM1  ;
 logic signed [31:0] O2_N6_S0;		always @(posedge clk) O2_N6_S0 <=     O2_I2_R2_C0_SM1   +  O2_I2_R2_C1_SM1  ;
 logic signed [31:0] O2_N8_S0;		always @(posedge clk) O2_N8_S0 <=     O2_I2_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O2_N0_S1;		always @(posedge clk) O2_N0_S1 <=     O2_N0_S0  +  O2_N2_S0 ;
 logic signed [31:0] O2_N2_S1;		always @(posedge clk) O2_N2_S1 <=     O2_N4_S0  +  O2_N6_S0 ;
 logic signed [31:0] O2_N4_S1;		always @(posedge clk) O2_N4_S1 <=     O2_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O2_N0_S2;		always @(posedge clk) O2_N0_S2 <=     O2_N0_S1  +  O2_N2_S1 ;
 logic signed [31:0] O2_N2_S2;		always @(posedge clk) O2_N2_S2 <=     O2_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O2_N0_S3;		always @(posedge clk) O2_N0_S3 <=     O2_N0_S2  +  O2_N2_S2 ;
 assign conv_mac_2 = O2_N0_S3;

logic signed [31:0] conv_mac_3;
logic signed [31:0] O3_N0_S0;		always @(posedge clk) O3_N0_S0 <=     O3_I3_R0_C0_SM1   +  O3_I3_R0_C1_SM1  ;
 logic signed [31:0] O3_N2_S0;		always @(posedge clk) O3_N2_S0 <=     O3_I3_R0_C2_SM1   +  O3_I3_R1_C0_SM1  ;
 logic signed [31:0] O3_N4_S0;		always @(posedge clk) O3_N4_S0 <=     O3_I3_R1_C1_SM1   +  O3_I3_R1_C2_SM1  ;
 logic signed [31:0] O3_N6_S0;		always @(posedge clk) O3_N6_S0 <=     O3_I3_R2_C0_SM1   +  O3_I3_R2_C1_SM1  ;
 logic signed [31:0] O3_N8_S0;		always @(posedge clk) O3_N8_S0 <=     O3_I3_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O3_N0_S1;		always @(posedge clk) O3_N0_S1 <=     O3_N0_S0  +  O3_N2_S0 ;
 logic signed [31:0] O3_N2_S1;		always @(posedge clk) O3_N2_S1 <=     O3_N4_S0  +  O3_N6_S0 ;
 logic signed [31:0] O3_N4_S1;		always @(posedge clk) O3_N4_S1 <=     O3_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O3_N0_S2;		always @(posedge clk) O3_N0_S2 <=     O3_N0_S1  +  O3_N2_S1 ;
 logic signed [31:0] O3_N2_S2;		always @(posedge clk) O3_N2_S2 <=     O3_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O3_N0_S3;		always @(posedge clk) O3_N0_S3 <=     O3_N0_S2  +  O3_N2_S2 ;
 assign conv_mac_3 = O3_N0_S3;

logic signed [31:0] conv_mac_4;
logic signed [31:0] O4_N0_S0;		always @(posedge clk) O4_N0_S0 <=     O4_I4_R0_C0_SM1   +  O4_I4_R0_C1_SM1  ;
 logic signed [31:0] O4_N2_S0;		always @(posedge clk) O4_N2_S0 <=     O4_I4_R0_C2_SM1   +  O4_I4_R1_C0_SM1  ;
 logic signed [31:0] O4_N4_S0;		always @(posedge clk) O4_N4_S0 <=     O4_I4_R1_C1_SM1   +  O4_I4_R1_C2_SM1  ;
 logic signed [31:0] O4_N6_S0;		always @(posedge clk) O4_N6_S0 <=     O4_I4_R2_C0_SM1   +  O4_I4_R2_C1_SM1  ;
 logic signed [31:0] O4_N8_S0;		always @(posedge clk) O4_N8_S0 <=     O4_I4_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O4_N0_S1;		always @(posedge clk) O4_N0_S1 <=     O4_N0_S0  +  O4_N2_S0 ;
 logic signed [31:0] O4_N2_S1;		always @(posedge clk) O4_N2_S1 <=     O4_N4_S0  +  O4_N6_S0 ;
 logic signed [31:0] O4_N4_S1;		always @(posedge clk) O4_N4_S1 <=     O4_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O4_N0_S2;		always @(posedge clk) O4_N0_S2 <=     O4_N0_S1  +  O4_N2_S1 ;
 logic signed [31:0] O4_N2_S2;		always @(posedge clk) O4_N2_S2 <=     O4_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O4_N0_S3;		always @(posedge clk) O4_N0_S3 <=     O4_N0_S2  +  O4_N2_S2 ;
 assign conv_mac_4 = O4_N0_S3;

logic signed [31:0] conv_mac_5;
logic signed [31:0] O5_N0_S0;		always @(posedge clk) O5_N0_S0 <=     O5_I5_R0_C0_SM1   +  O5_I5_R0_C1_SM1  ;
 logic signed [31:0] O5_N2_S0;		always @(posedge clk) O5_N2_S0 <=     O5_I5_R0_C2_SM1   +  O5_I5_R1_C0_SM1  ;
 logic signed [31:0] O5_N4_S0;		always @(posedge clk) O5_N4_S0 <=     O5_I5_R1_C1_SM1   +  O5_I5_R1_C2_SM1  ;
 logic signed [31:0] O5_N6_S0;		always @(posedge clk) O5_N6_S0 <=     O5_I5_R2_C0_SM1   +  O5_I5_R2_C1_SM1  ;
 logic signed [31:0] O5_N8_S0;		always @(posedge clk) O5_N8_S0 <=     O5_I5_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O5_N0_S1;		always @(posedge clk) O5_N0_S1 <=     O5_N0_S0  +  O5_N2_S0 ;
 logic signed [31:0] O5_N2_S1;		always @(posedge clk) O5_N2_S1 <=     O5_N4_S0  +  O5_N6_S0 ;
 logic signed [31:0] O5_N4_S1;		always @(posedge clk) O5_N4_S1 <=     O5_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O5_N0_S2;		always @(posedge clk) O5_N0_S2 <=     O5_N0_S1  +  O5_N2_S1 ;
 logic signed [31:0] O5_N2_S2;		always @(posedge clk) O5_N2_S2 <=     O5_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O5_N0_S3;		always @(posedge clk) O5_N0_S3 <=     O5_N0_S2  +  O5_N2_S2 ;
 assign conv_mac_5 = O5_N0_S3;

logic signed [31:0] conv_mac_6;
logic signed [31:0] O6_N0_S0;		always @(posedge clk) O6_N0_S0 <=     O6_I6_R0_C0_SM1   +  O6_I6_R0_C1_SM1  ;
 logic signed [31:0] O6_N2_S0;		always @(posedge clk) O6_N2_S0 <=     O6_I6_R0_C2_SM1   +  O6_I6_R1_C0_SM1  ;
 logic signed [31:0] O6_N4_S0;		always @(posedge clk) O6_N4_S0 <=     O6_I6_R1_C1_SM1   +  O6_I6_R1_C2_SM1  ;
 logic signed [31:0] O6_N6_S0;		always @(posedge clk) O6_N6_S0 <=     O6_I6_R2_C0_SM1   +  O6_I6_R2_C1_SM1  ;
 logic signed [31:0] O6_N8_S0;		always @(posedge clk) O6_N8_S0 <=     O6_I6_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O6_N0_S1;		always @(posedge clk) O6_N0_S1 <=     O6_N0_S0  +  O6_N2_S0 ;
 logic signed [31:0] O6_N2_S1;		always @(posedge clk) O6_N2_S1 <=     O6_N4_S0  +  O6_N6_S0 ;
 logic signed [31:0] O6_N4_S1;		always @(posedge clk) O6_N4_S1 <=     O6_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O6_N0_S2;		always @(posedge clk) O6_N0_S2 <=     O6_N0_S1  +  O6_N2_S1 ;
 logic signed [31:0] O6_N2_S2;		always @(posedge clk) O6_N2_S2 <=     O6_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O6_N0_S3;		always @(posedge clk) O6_N0_S3 <=     O6_N0_S2  +  O6_N2_S2 ;
 assign conv_mac_6 = O6_N0_S3;

logic signed [31:0] conv_mac_7;
logic signed [31:0] O7_N0_S0;		always @(posedge clk) O7_N0_S0 <=     O7_I7_R0_C0_SM1   +  O7_I7_R0_C1_SM1  ;
 logic signed [31:0] O7_N2_S0;		always @(posedge clk) O7_N2_S0 <=     O7_I7_R0_C2_SM1   +  O7_I7_R1_C0_SM1  ;
 logic signed [31:0] O7_N4_S0;		always @(posedge clk) O7_N4_S0 <=     O7_I7_R1_C1_SM1   +  O7_I7_R1_C2_SM1  ;
 logic signed [31:0] O7_N6_S0;		always @(posedge clk) O7_N6_S0 <=     O7_I7_R2_C0_SM1   +  O7_I7_R2_C1_SM1  ;
 logic signed [31:0] O7_N8_S0;		always @(posedge clk) O7_N8_S0 <=     O7_I7_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O7_N0_S1;		always @(posedge clk) O7_N0_S1 <=     O7_N0_S0  +  O7_N2_S0 ;
 logic signed [31:0] O7_N2_S1;		always @(posedge clk) O7_N2_S1 <=     O7_N4_S0  +  O7_N6_S0 ;
 logic signed [31:0] O7_N4_S1;		always @(posedge clk) O7_N4_S1 <=     O7_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O7_N0_S2;		always @(posedge clk) O7_N0_S2 <=     O7_N0_S1  +  O7_N2_S1 ;
 logic signed [31:0] O7_N2_S2;		always @(posedge clk) O7_N2_S2 <=     O7_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O7_N0_S3;		always @(posedge clk) O7_N0_S3 <=     O7_N0_S2  +  O7_N2_S2 ;
 assign conv_mac_7 = O7_N0_S3;

logic valid_D1;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D1<= 0 ;
	else valid_D1<=valid;
end
logic valid_D2;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D2<= 0 ;
	else valid_D2<=valid_D1;
end
logic valid_D3;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D3<= 0 ;
	else valid_D3<=valid_D2;
end
logic valid_D4;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D4<= 0 ;
	else valid_D4<=valid_D3;
end
logic valid_D5;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D5<= 0 ;
	else valid_D5<=valid_D4;
end
always_ff @(posedge clk) begin
	if (rstn == 0) ready <= 0 ;
	else ready <=valid_D5;
end
logic [31:0] bias_add_0;
assign bias_add_0 = conv_mac_0 + 7'd41;
logic [31:0] bias_add_1;
assign bias_add_1 = conv_mac_1 + 6'd19;
logic [31:0] bias_add_2;
assign bias_add_2 = conv_mac_2 - 4'd7;
logic [31:0] bias_add_3;
assign bias_add_3 = conv_mac_3 + 7'd46;
logic [31:0] bias_add_4;
assign bias_add_4 = conv_mac_4 - 6'd22;
logic [31:0] bias_add_5;
assign bias_add_5 = conv_mac_5 + 6'd27;
logic [31:0] bias_add_6;
assign bias_add_6 = conv_mac_6 + 5'd14;
logic [31:0] bias_add_7;
assign bias_add_7 = conv_mac_7 + 7'd34;

logic [7:0] relu_0;
assign relu_0[7:0] = (bias_add_0[31]==0) ? ((bias_add_0<3'd6) ? {{bias_add_0[31],bias_add_0[10:4]}} :'d6) : '0;
logic [7:0] relu_1;
assign relu_1[7:0] = (bias_add_1[31]==0) ? ((bias_add_1<3'd6) ? {{bias_add_1[31],bias_add_1[10:4]}} :'d6) : '0;
logic [7:0] relu_2;
assign relu_2[7:0] = (bias_add_2[31]==0) ? ((bias_add_2<3'd6) ? {{bias_add_2[31],bias_add_2[10:4]}} :'d6) : '0;
logic [7:0] relu_3;
assign relu_3[7:0] = (bias_add_3[31]==0) ? ((bias_add_3<3'd6) ? {{bias_add_3[31],bias_add_3[10:4]}} :'d6) : '0;
logic [7:0] relu_4;
assign relu_4[7:0] = (bias_add_4[31]==0) ? ((bias_add_4<3'd6) ? {{bias_add_4[31],bias_add_4[10:4]}} :'d6) : '0;
logic [7:0] relu_5;
assign relu_5[7:0] = (bias_add_5[31]==0) ? ((bias_add_5<3'd6) ? {{bias_add_5[31],bias_add_5[10:4]}} :'d6) : '0;
logic [7:0] relu_6;
assign relu_6[7:0] = (bias_add_6[31]==0) ? ((bias_add_6<3'd6) ? {{bias_add_6[31],bias_add_6[10:4]}} :'d6) : '0;
logic [7:0] relu_7;
assign relu_7[7:0] = (bias_add_7[31]==0) ? ((bias_add_7<3'd6) ? {{bias_add_7[31],bias_add_7[10:4]}} :'d6) : '0;

assign output_act = {
	relu_7,
	relu_6,
	relu_5,
	relu_4,
	relu_3,
	relu_2,
	relu_1,
	relu_0
};

endmodule
module conv2_dw (
    input logic clk,
    input logic rstn,
    input logic valid,
    input logic [8*72-1:0] input_act,
    output logic [64-1:0] output_act,
    output logic ready
);
logic we;
logic [8:0] zero_number; 
assign zero_number = 9'd0; 
logic [8*72-1:0] input_act_ff;
genvar i;
generate
for (i=0;i<8;i++)
    begin: genblk_7
        always_ff @(posedge clk) begin
            if (rstn == 0) begin
                input_act_ff[(i+1)*72-1:i*72] <= '0;
            end
            else begin
                input_act_ff[(i+1)*72-1:i*72] <= input_act[(i+1)*72-1:i*72];
            end
        end
    end
endgenerate
logic [71:0] input_fmap_0;
assign input_fmap_0 = input_act_ff[71:0];
logic [71:0] input_fmap_1;
assign input_fmap_1 = input_act_ff[143:72];
logic [71:0] input_fmap_2;
assign input_fmap_2 = input_act_ff[215:144];
logic [71:0] input_fmap_3;
assign input_fmap_3 = input_act_ff[287:216];
logic [71:0] input_fmap_4;
assign input_fmap_4 = input_act_ff[359:288];
logic [71:0] input_fmap_5;
assign input_fmap_5 = input_act_ff[431:360];
logic [71:0] input_fmap_6;
assign input_fmap_6 = input_act_ff[503:432];
logic [71:0] input_fmap_7;
assign input_fmap_7 = input_act_ff[575:504];

logic [13-1:0] O0_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_dw_O0_I0_R0_C09_rom_inst (.q(O0_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O0_I0_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O0_I0_R0_C09_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_dw_O0_I0_R0_C09_rom_inst (.q(O0_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [11-1:0] O0_I0_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_dw_O0_I0_R0_C13_rom_inst (.q(O0_I0_R0_C1_SM1 ),.address(input_fmap_0[15:8]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R0_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O0_I0_R0_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O0_I0_R0_C13_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_dw_O0_I0_R0_C13_rom_inst (.q(O0_I0_R0_C1_SM1 ),.address(input_fmap_0[15:8]),.clock  (clk));
logic [10-1:0] O0_I0_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv2_dw_O0_I0_R0_C21_rom_inst (.q(O0_I0_R0_C2_SM1 ),.address(input_fmap_0[23:16]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R0_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O0_I0_R0_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O0_I0_R0_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv2_dw_O0_I0_R0_C21_rom_inst (.q(O0_I0_R0_C2_SM1 ),.address(input_fmap_0[23:16]),.clock  (clk));
logic [12-1:0] O0_I0_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv2_dw_O0_I0_R1_C06_rom_inst (.q(O0_I0_R1_C0_SM1 ),.address(input_fmap_0[31:24]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R1_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O0_I0_R1_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O0_I0_R1_C06_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv2_dw_O0_I0_R1_C06_rom_inst (.q(O0_I0_R1_C0_SM1 ),.address(input_fmap_0[31:24]),.clock  (clk));
logic [14-1:0] O0_I0_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv2_dw_O0_I0_R1_C120_rom_inst (.q(O0_I0_R1_C1_SM1 ),.address(input_fmap_0[39:32]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R1_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O0_I0_R1_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O0_I0_R1_C120_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv2_dw_O0_I0_R1_C120_rom_inst (.q(O0_I0_R1_C1_SM1 ),.address(input_fmap_0[39:32]),.clock  (clk));
logic [13-1:0] O0_I0_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_dw_O0_I0_R1_C28_rom_inst (.q(O0_I0_R1_C2_SM1 ),.address(input_fmap_0[47:40]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R1_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O0_I0_R1_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O0_I0_R1_C28_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_dw_O0_I0_R1_C28_rom_inst (.q(O0_I0_R1_C2_SM1 ),.address(input_fmap_0[47:40]),.clock  (clk));
logic [13-1:0] O0_I0_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_dw_O0_I0_R2_C011_rom_inst (.q(O0_I0_R2_C0_SM1 ),.address(input_fmap_0[55:48]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R2_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O0_I0_R2_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O0_I0_R2_C011_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_dw_O0_I0_R2_C011_rom_inst (.q(O0_I0_R2_C0_SM1 ),.address(input_fmap_0[55:48]),.clock  (clk));
logic [14-1:0] O0_I0_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv2_dw_O0_I0_R2_C128_rom_inst (.q(O0_I0_R2_C1_SM1 ),.address(input_fmap_0[63:56]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R2_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O0_I0_R2_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O0_I0_R2_C128_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv2_dw_O0_I0_R2_C128_rom_inst (.q(O0_I0_R2_C1_SM1 ),.address(input_fmap_0[63:56]),.clock  (clk));
logic [12-1:0] O0_I0_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv2_dw_O0_I0_R2_C26_rom_inst (.q(O0_I0_R2_C2_SM1 ),.address(input_fmap_0[71:64]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R2_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O0_I0_R2_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O0_I0_R2_C26_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv2_dw_O0_I0_R2_C26_rom_inst (.q(O0_I0_R2_C2_SM1 ),.address(input_fmap_0[71:64]),.clock  (clk));
logic [14-1:0] O1_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv2_dw_O1_I1_R0_C016_rom_inst (.q(O1_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R0_C0_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O1_I1_R0_C0_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O1_I1_R0_C016_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv2_dw_O1_I1_R0_C016_rom_inst (.q(O1_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [14-1:0] O1_I1_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv2_dw_O1_I1_R0_C127_rom_inst (.q(O1_I1_R0_C1_SM1 ),.address(input_fmap_1[15:8]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R0_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O1_I1_R0_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O1_I1_R0_C127_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv2_dw_O1_I1_R0_C127_rom_inst (.q(O1_I1_R0_C1_SM1 ),.address(input_fmap_1[15:8]),.clock  (clk));
logic [13-1:0] O1_I1_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_dw_O1_I1_R0_C28_rom_inst (.q(O1_I1_R0_C2_SM1 ),.address(input_fmap_1[23:16]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R0_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O1_I1_R0_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O1_I1_R0_C28_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_dw_O1_I1_R0_C28_rom_inst (.q(O1_I1_R0_C2_SM1 ),.address(input_fmap_1[23:16]),.clock  (clk));
logic [14-1:0] O1_I1_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv2_dw_O1_I1_R1_C024_rom_inst (.q(O1_I1_R1_C0_SM1 ),.address(input_fmap_1[31:24]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R1_C0_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O1_I1_R1_C0_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O1_I1_R1_C024_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv2_dw_O1_I1_R1_C024_rom_inst (.q(O1_I1_R1_C0_SM1 ),.address(input_fmap_1[31:24]),.clock  (clk));
logic [15-1:0] O1_I1_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(15),.INIT_FILE("deepfreeze_rom/deepfreeze_8_15.txt"))
    conv2_dw_O1_I1_R1_C141_rom_inst (.q(O1_I1_R1_C1_SM1 ),.address(input_fmap_1[39:32]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R1_C1_SM1  = 15'h1234;
//always@(posedge clk) begin 
//O1_I1_R1_C1_SM1  <= 15'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O1_I1_R1_C141_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(15))
//    conv2_dw_O1_I1_R1_C141_rom_inst (.q(O1_I1_R1_C1_SM1 ),.address(input_fmap_1[39:32]),.clock  (clk));
logic [13-1:0] O1_I1_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_dw_O1_I1_R1_C215_rom_inst (.q(O1_I1_R1_C2_SM1 ),.address(input_fmap_1[47:40]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R1_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O1_I1_R1_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O1_I1_R1_C215_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_dw_O1_I1_R1_C215_rom_inst (.q(O1_I1_R1_C2_SM1 ),.address(input_fmap_1[47:40]),.clock  (clk));
logic [13-1:0] O1_I1_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_dw_O1_I1_R2_C09_rom_inst (.q(O1_I1_R2_C0_SM1 ),.address(input_fmap_1[55:48]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R2_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O1_I1_R2_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O1_I1_R2_C09_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_dw_O1_I1_R2_C09_rom_inst (.q(O1_I1_R2_C0_SM1 ),.address(input_fmap_1[55:48]),.clock  (clk));
logic [13-1:0] O1_I1_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_dw_O1_I1_R2_C115_rom_inst (.q(O1_I1_R2_C1_SM1 ),.address(input_fmap_1[63:56]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R2_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O1_I1_R2_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O1_I1_R2_C115_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_dw_O1_I1_R2_C115_rom_inst (.q(O1_I1_R2_C1_SM1 ),.address(input_fmap_1[63:56]),.clock  (clk));
logic [13-1:0] O2_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_dw_O2_I2_R0_C012_rom_inst (.q(O2_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O2_I2_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O2_I2_R0_C012_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_dw_O2_I2_R0_C012_rom_inst (.q(O2_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [14-1:0] O2_I2_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv2_dw_O2_I2_R0_C119_rom_inst (.q(O2_I2_R0_C1_SM1 ),.address(input_fmap_2[15:8]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R0_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O2_I2_R0_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O2_I2_R0_C119_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv2_dw_O2_I2_R0_C119_rom_inst (.q(O2_I2_R0_C1_SM1 ),.address(input_fmap_2[15:8]),.clock  (clk));
logic [11-1:0] O2_I2_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_dw_O2_I2_R0_C22_rom_inst (.q(O2_I2_R0_C2_SM1 ),.address(input_fmap_2[23:16]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R0_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O2_I2_R0_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O2_I2_R0_C22_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_dw_O2_I2_R0_C22_rom_inst (.q(O2_I2_R0_C2_SM1 ),.address(input_fmap_2[23:16]),.clock  (clk));
logic [13-1:0] O2_I2_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_dw_O2_I2_R1_C014_rom_inst (.q(O2_I2_R1_C0_SM1 ),.address(input_fmap_2[31:24]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R1_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O2_I2_R1_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O2_I2_R1_C014_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_dw_O2_I2_R1_C014_rom_inst (.q(O2_I2_R1_C0_SM1 ),.address(input_fmap_2[31:24]),.clock  (clk));
logic [14-1:0] O2_I2_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv2_dw_O2_I2_R1_C120_rom_inst (.q(O2_I2_R1_C1_SM1 ),.address(input_fmap_2[39:32]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R1_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O2_I2_R1_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O2_I2_R1_C120_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv2_dw_O2_I2_R1_C120_rom_inst (.q(O2_I2_R1_C1_SM1 ),.address(input_fmap_2[39:32]),.clock  (clk));
logic [13-1:0] O2_I2_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_dw_O2_I2_R1_C210_rom_inst (.q(O2_I2_R1_C2_SM1 ),.address(input_fmap_2[47:40]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R1_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O2_I2_R1_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O2_I2_R1_C210_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_dw_O2_I2_R1_C210_rom_inst (.q(O2_I2_R1_C2_SM1 ),.address(input_fmap_2[47:40]),.clock  (clk));
logic [12-1:0] O2_I2_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv2_dw_O2_I2_R2_C07_rom_inst (.q(O2_I2_R2_C0_SM1 ),.address(input_fmap_2[55:48]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R2_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O2_I2_R2_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O2_I2_R2_C07_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv2_dw_O2_I2_R2_C07_rom_inst (.q(O2_I2_R2_C0_SM1 ),.address(input_fmap_2[55:48]),.clock  (clk));
logic [13-1:0] O2_I2_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_dw_O2_I2_R2_C115_rom_inst (.q(O2_I2_R2_C1_SM1 ),.address(input_fmap_2[63:56]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R2_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O2_I2_R2_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O2_I2_R2_C115_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_dw_O2_I2_R2_C115_rom_inst (.q(O2_I2_R2_C1_SM1 ),.address(input_fmap_2[63:56]),.clock  (clk));
logic [12-1:0] O2_I2_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv2_dw_O2_I2_R2_C27_rom_inst (.q(O2_I2_R2_C2_SM1 ),.address(input_fmap_2[71:64]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R2_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O2_I2_R2_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O2_I2_R2_C27_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv2_dw_O2_I2_R2_C27_rom_inst (.q(O2_I2_R2_C2_SM1 ),.address(input_fmap_2[71:64]),.clock  (clk));
logic [14-1:0] O3_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv2_dw_O3_I3_R0_C016_rom_inst (.q(O3_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R0_C0_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O3_I3_R0_C0_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O3_I3_R0_C016_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv2_dw_O3_I3_R0_C016_rom_inst (.q(O3_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [13-1:0] O3_I3_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_dw_O3_I3_R0_C19_rom_inst (.q(O3_I3_R0_C1_SM1 ),.address(input_fmap_3[15:8]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R0_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O3_I3_R0_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O3_I3_R0_C19_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_dw_O3_I3_R0_C19_rom_inst (.q(O3_I3_R0_C1_SM1 ),.address(input_fmap_3[15:8]),.clock  (clk));
logic [11-1:0] O3_I3_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_dw_O3_I3_R0_C23_rom_inst (.q(O3_I3_R0_C2_SM1 ),.address(input_fmap_3[23:16]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R0_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O3_I3_R0_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O3_I3_R0_C23_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_dw_O3_I3_R0_C23_rom_inst (.q(O3_I3_R0_C2_SM1 ),.address(input_fmap_3[23:16]),.clock  (clk));
logic [15-1:0] O3_I3_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(15),.INIT_FILE("deepfreeze_rom/deepfreeze_8_15.txt"))
    conv2_dw_O3_I3_R1_C037_rom_inst (.q(O3_I3_R1_C0_SM1 ),.address(input_fmap_3[31:24]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R1_C0_SM1  = 15'h1234;
//always@(posedge clk) begin 
//O3_I3_R1_C0_SM1  <= 15'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O3_I3_R1_C037_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(15))
//    conv2_dw_O3_I3_R1_C037_rom_inst (.q(O3_I3_R1_C0_SM1 ),.address(input_fmap_3[31:24]),.clock  (clk));
logic [14-1:0] O3_I3_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv2_dw_O3_I3_R1_C122_rom_inst (.q(O3_I3_R1_C1_SM1 ),.address(input_fmap_3[39:32]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R1_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O3_I3_R1_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O3_I3_R1_C122_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv2_dw_O3_I3_R1_C122_rom_inst (.q(O3_I3_R1_C1_SM1 ),.address(input_fmap_3[39:32]),.clock  (clk));
logic [11-1:0] O3_I3_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_dw_O3_I3_R1_C22_rom_inst (.q(O3_I3_R1_C2_SM1 ),.address(input_fmap_3[47:40]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R1_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O3_I3_R1_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O3_I3_R1_C22_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_dw_O3_I3_R1_C22_rom_inst (.q(O3_I3_R1_C2_SM1 ),.address(input_fmap_3[47:40]),.clock  (clk));
logic [13-1:0] O3_I3_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_dw_O3_I3_R2_C014_rom_inst (.q(O3_I3_R2_C0_SM1 ),.address(input_fmap_3[55:48]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R2_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O3_I3_R2_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O3_I3_R2_C014_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_dw_O3_I3_R2_C014_rom_inst (.q(O3_I3_R2_C0_SM1 ),.address(input_fmap_3[55:48]),.clock  (clk));
logic [13-1:0] O3_I3_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_dw_O3_I3_R2_C112_rom_inst (.q(O3_I3_R2_C1_SM1 ),.address(input_fmap_3[63:56]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R2_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O3_I3_R2_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O3_I3_R2_C112_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_dw_O3_I3_R2_C112_rom_inst (.q(O3_I3_R2_C1_SM1 ),.address(input_fmap_3[63:56]),.clock  (clk));
logic [11-1:0] O3_I3_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_dw_O3_I3_R2_C22_rom_inst (.q(O3_I3_R2_C2_SM1 ),.address(input_fmap_3[71:64]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R2_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O3_I3_R2_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O3_I3_R2_C22_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_dw_O3_I3_R2_C22_rom_inst (.q(O3_I3_R2_C2_SM1 ),.address(input_fmap_3[71:64]),.clock  (clk));
logic [13-1:0] O4_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_dw_O4_I4_R0_C08_rom_inst (.q(O4_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O4_I4_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O4_I4_R0_C08_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_dw_O4_I4_R0_C08_rom_inst (.q(O4_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [13-1:0] O4_I4_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_dw_O4_I4_R0_C112_rom_inst (.q(O4_I4_R0_C1_SM1 ),.address(input_fmap_4[15:8]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R0_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O4_I4_R0_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O4_I4_R0_C112_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_dw_O4_I4_R0_C112_rom_inst (.q(O4_I4_R0_C1_SM1 ),.address(input_fmap_4[15:8]),.clock  (clk));
logic [11-1:0] O4_I4_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_dw_O4_I4_R0_C22_rom_inst (.q(O4_I4_R0_C2_SM1 ),.address(input_fmap_4[23:16]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R0_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O4_I4_R0_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O4_I4_R0_C22_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_dw_O4_I4_R0_C22_rom_inst (.q(O4_I4_R0_C2_SM1 ),.address(input_fmap_4[23:16]),.clock  (clk));
logic [14-1:0] O4_I4_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv2_dw_O4_I4_R1_C019_rom_inst (.q(O4_I4_R1_C0_SM1 ),.address(input_fmap_4[31:24]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R1_C0_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O4_I4_R1_C0_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O4_I4_R1_C019_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv2_dw_O4_I4_R1_C019_rom_inst (.q(O4_I4_R1_C0_SM1 ),.address(input_fmap_4[31:24]),.clock  (clk));
logic [14-1:0] O4_I4_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv2_dw_O4_I4_R1_C123_rom_inst (.q(O4_I4_R1_C1_SM1 ),.address(input_fmap_4[39:32]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R1_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O4_I4_R1_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O4_I4_R1_C123_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv2_dw_O4_I4_R1_C123_rom_inst (.q(O4_I4_R1_C1_SM1 ),.address(input_fmap_4[39:32]),.clock  (clk));
logic [12-1:0] O4_I4_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv2_dw_O4_I4_R1_C26_rom_inst (.q(O4_I4_R1_C2_SM1 ),.address(input_fmap_4[47:40]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R1_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O4_I4_R1_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O4_I4_R1_C26_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv2_dw_O4_I4_R1_C26_rom_inst (.q(O4_I4_R1_C2_SM1 ),.address(input_fmap_4[47:40]),.clock  (clk));
logic [13-1:0] O4_I4_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_dw_O4_I4_R2_C011_rom_inst (.q(O4_I4_R2_C0_SM1 ),.address(input_fmap_4[55:48]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R2_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O4_I4_R2_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O4_I4_R2_C011_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_dw_O4_I4_R2_C011_rom_inst (.q(O4_I4_R2_C0_SM1 ),.address(input_fmap_4[55:48]),.clock  (clk));
logic [13-1:0] O4_I4_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_dw_O4_I4_R2_C114_rom_inst (.q(O4_I4_R2_C1_SM1 ),.address(input_fmap_4[63:56]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R2_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O4_I4_R2_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O4_I4_R2_C114_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_dw_O4_I4_R2_C114_rom_inst (.q(O4_I4_R2_C1_SM1 ),.address(input_fmap_4[63:56]),.clock  (clk));
logic [11-1:0] O4_I4_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_dw_O4_I4_R2_C23_rom_inst (.q(O4_I4_R2_C2_SM1 ),.address(input_fmap_4[71:64]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R2_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O4_I4_R2_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O4_I4_R2_C23_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_dw_O4_I4_R2_C23_rom_inst (.q(O4_I4_R2_C2_SM1 ),.address(input_fmap_4[71:64]),.clock  (clk));
logic [12-1:0] O5_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv2_dw_O5_I5_R0_C04_rom_inst (.q(O5_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O5_I5_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O5_I5_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv2_dw_O5_I5_R0_C04_rom_inst (.q(O5_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [10-1:0] O5_I5_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv2_dw_O5_I5_R0_C11_rom_inst (.q(O5_I5_R0_C1_SM1 ),.address(input_fmap_5[15:8]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R0_C1_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I5_R0_C1_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O5_I5_R0_C11_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv2_dw_O5_I5_R0_C11_rom_inst (.q(O5_I5_R0_C1_SM1 ),.address(input_fmap_5[15:8]),.clock  (clk));
logic [11-1:0] O5_I5_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_dw_O5_I5_R0_C22_rom_inst (.q(O5_I5_R0_C2_SM1 ),.address(input_fmap_5[23:16]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R0_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O5_I5_R0_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O5_I5_R0_C22_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_dw_O5_I5_R0_C22_rom_inst (.q(O5_I5_R0_C2_SM1 ),.address(input_fmap_5[23:16]),.clock  (clk));
logic [11-1:0] O5_I5_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_dw_O5_I5_R1_C03_rom_inst (.q(O5_I5_R1_C0_SM1 ),.address(input_fmap_5[31:24]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R1_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O5_I5_R1_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O5_I5_R1_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_dw_O5_I5_R1_C03_rom_inst (.q(O5_I5_R1_C0_SM1 ),.address(input_fmap_5[31:24]),.clock  (clk));
logic [12-1:0] O5_I5_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv2_dw_O5_I5_R1_C16_rom_inst (.q(O5_I5_R1_C1_SM1 ),.address(input_fmap_5[39:32]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R1_C1_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O5_I5_R1_C1_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O5_I5_R1_C16_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv2_dw_O5_I5_R1_C16_rom_inst (.q(O5_I5_R1_C1_SM1 ),.address(input_fmap_5[39:32]),.clock  (clk));
logic [12-1:0] O5_I5_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv2_dw_O5_I5_R1_C24_rom_inst (.q(O5_I5_R1_C2_SM1 ),.address(input_fmap_5[47:40]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R1_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O5_I5_R1_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O5_I5_R1_C24_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv2_dw_O5_I5_R1_C24_rom_inst (.q(O5_I5_R1_C2_SM1 ),.address(input_fmap_5[47:40]),.clock  (clk));
logic [13-1:0] O5_I5_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_dw_O5_I5_R2_C010_rom_inst (.q(O5_I5_R2_C0_SM1 ),.address(input_fmap_5[55:48]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R2_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O5_I5_R2_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O5_I5_R2_C010_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_dw_O5_I5_R2_C010_rom_inst (.q(O5_I5_R2_C0_SM1 ),.address(input_fmap_5[55:48]),.clock  (clk));
logic [14-1:0] O5_I5_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv2_dw_O5_I5_R2_C117_rom_inst (.q(O5_I5_R2_C1_SM1 ),.address(input_fmap_5[63:56]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R2_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O5_I5_R2_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O5_I5_R2_C117_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv2_dw_O5_I5_R2_C117_rom_inst (.q(O5_I5_R2_C1_SM1 ),.address(input_fmap_5[63:56]),.clock  (clk));
logic [12-1:0] O5_I5_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv2_dw_O5_I5_R2_C25_rom_inst (.q(O5_I5_R2_C2_SM1 ),.address(input_fmap_5[71:64]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R2_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O5_I5_R2_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O5_I5_R2_C25_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv2_dw_O5_I5_R2_C25_rom_inst (.q(O5_I5_R2_C2_SM1 ),.address(input_fmap_5[71:64]),.clock  (clk));
logic [14-1:0] O6_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv2_dw_O6_I6_R0_C016_rom_inst (.q(O6_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R0_C0_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O6_I6_R0_C0_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O6_I6_R0_C016_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv2_dw_O6_I6_R0_C016_rom_inst (.q(O6_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [12-1:0] O6_I6_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv2_dw_O6_I6_R0_C14_rom_inst (.q(O6_I6_R0_C1_SM1 ),.address(input_fmap_6[15:8]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R0_C1_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O6_I6_R0_C1_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O6_I6_R0_C14_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv2_dw_O6_I6_R0_C14_rom_inst (.q(O6_I6_R0_C1_SM1 ),.address(input_fmap_6[15:8]),.clock  (clk));
logic [12-1:0] O6_I6_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv2_dw_O6_I6_R0_C24_rom_inst (.q(O6_I6_R0_C2_SM1 ),.address(input_fmap_6[23:16]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R0_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O6_I6_R0_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O6_I6_R0_C24_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv2_dw_O6_I6_R0_C24_rom_inst (.q(O6_I6_R0_C2_SM1 ),.address(input_fmap_6[23:16]),.clock  (clk));
logic [15-1:0] O6_I6_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(15),.INIT_FILE("deepfreeze_rom/deepfreeze_8_15.txt"))
    conv2_dw_O6_I6_R1_C033_rom_inst (.q(O6_I6_R1_C0_SM1 ),.address(input_fmap_6[31:24]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R1_C0_SM1  = 15'h1234;
//always@(posedge clk) begin 
//O6_I6_R1_C0_SM1  <= 15'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O6_I6_R1_C033_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(15))
//    conv2_dw_O6_I6_R1_C033_rom_inst (.q(O6_I6_R1_C0_SM1 ),.address(input_fmap_6[31:24]),.clock  (clk));
logic [13-1:0] O6_I6_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_dw_O6_I6_R1_C115_rom_inst (.q(O6_I6_R1_C1_SM1 ),.address(input_fmap_6[39:32]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R1_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O6_I6_R1_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O6_I6_R1_C115_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_dw_O6_I6_R1_C115_rom_inst (.q(O6_I6_R1_C1_SM1 ),.address(input_fmap_6[39:32]),.clock  (clk));
logic [14-1:0] O6_I6_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv2_dw_O6_I6_R1_C221_rom_inst (.q(O6_I6_R1_C2_SM1 ),.address(input_fmap_6[47:40]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R1_C2_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O6_I6_R1_C2_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O6_I6_R1_C221_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv2_dw_O6_I6_R1_C221_rom_inst (.q(O6_I6_R1_C2_SM1 ),.address(input_fmap_6[47:40]),.clock  (clk));
logic [14-1:0] O6_I6_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv2_dw_O6_I6_R2_C031_rom_inst (.q(O6_I6_R2_C0_SM1 ),.address(input_fmap_6[55:48]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R2_C0_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O6_I6_R2_C0_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O6_I6_R2_C031_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv2_dw_O6_I6_R2_C031_rom_inst (.q(O6_I6_R2_C0_SM1 ),.address(input_fmap_6[55:48]),.clock  (clk));
logic [13-1:0] O6_I6_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_dw_O6_I6_R2_C110_rom_inst (.q(O6_I6_R2_C1_SM1 ),.address(input_fmap_6[63:56]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R2_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O6_I6_R2_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O6_I6_R2_C110_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_dw_O6_I6_R2_C110_rom_inst (.q(O6_I6_R2_C1_SM1 ),.address(input_fmap_6[63:56]),.clock  (clk));
logic [13-1:0] O6_I6_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_dw_O6_I6_R2_C212_rom_inst (.q(O6_I6_R2_C2_SM1 ),.address(input_fmap_6[71:64]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R2_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O6_I6_R2_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O6_I6_R2_C212_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_dw_O6_I6_R2_C212_rom_inst (.q(O6_I6_R2_C2_SM1 ),.address(input_fmap_6[71:64]),.clock  (clk));
logic [13-1:0] O7_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_dw_O7_I7_R0_C012_rom_inst (.q(O7_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O7_I7_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O7_I7_R0_C012_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_dw_O7_I7_R0_C012_rom_inst (.q(O7_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [13-1:0] O7_I7_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_dw_O7_I7_R0_C115_rom_inst (.q(O7_I7_R0_C1_SM1 ),.address(input_fmap_7[15:8]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R0_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O7_I7_R0_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O7_I7_R0_C115_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_dw_O7_I7_R0_C115_rom_inst (.q(O7_I7_R0_C1_SM1 ),.address(input_fmap_7[15:8]),.clock  (clk));
logic [13-1:0] O7_I7_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_dw_O7_I7_R0_C28_rom_inst (.q(O7_I7_R0_C2_SM1 ),.address(input_fmap_7[23:16]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R0_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O7_I7_R0_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O7_I7_R0_C28_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_dw_O7_I7_R0_C28_rom_inst (.q(O7_I7_R0_C2_SM1 ),.address(input_fmap_7[23:16]),.clock  (clk));
logic [14-1:0] O7_I7_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv2_dw_O7_I7_R1_C019_rom_inst (.q(O7_I7_R1_C0_SM1 ),.address(input_fmap_7[31:24]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R1_C0_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O7_I7_R1_C0_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O7_I7_R1_C019_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv2_dw_O7_I7_R1_C019_rom_inst (.q(O7_I7_R1_C0_SM1 ),.address(input_fmap_7[31:24]),.clock  (clk));
logic [14-1:0] O7_I7_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv2_dw_O7_I7_R1_C125_rom_inst (.q(O7_I7_R1_C1_SM1 ),.address(input_fmap_7[39:32]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R1_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O7_I7_R1_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O7_I7_R1_C125_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv2_dw_O7_I7_R1_C125_rom_inst (.q(O7_I7_R1_C1_SM1 ),.address(input_fmap_7[39:32]),.clock  (clk));
logic [13-1:0] O7_I7_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_dw_O7_I7_R1_C212_rom_inst (.q(O7_I7_R1_C2_SM1 ),.address(input_fmap_7[47:40]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R1_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O7_I7_R1_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O7_I7_R1_C212_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_dw_O7_I7_R1_C212_rom_inst (.q(O7_I7_R1_C2_SM1 ),.address(input_fmap_7[47:40]),.clock  (clk));
logic [13-1:0] O7_I7_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_dw_O7_I7_R2_C010_rom_inst (.q(O7_I7_R2_C0_SM1 ),.address(input_fmap_7[55:48]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R2_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O7_I7_R2_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O7_I7_R2_C010_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_dw_O7_I7_R2_C010_rom_inst (.q(O7_I7_R2_C0_SM1 ),.address(input_fmap_7[55:48]),.clock  (clk));
logic [13-1:0] O7_I7_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_dw_O7_I7_R2_C115_rom_inst (.q(O7_I7_R2_C1_SM1 ),.address(input_fmap_7[63:56]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R2_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O7_I7_R2_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O7_I7_R2_C115_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_dw_O7_I7_R2_C115_rom_inst (.q(O7_I7_R2_C1_SM1 ),.address(input_fmap_7[63:56]),.clock  (clk));
logic [13-1:0] O7_I7_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_dw_O7_I7_R2_C210_rom_inst (.q(O7_I7_R2_C2_SM1 ),.address(input_fmap_7[71:64]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R2_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O7_I7_R2_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_dw_O7_I7_R2_C210_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_dw_O7_I7_R2_C210_rom_inst (.q(O7_I7_R2_C2_SM1 ),.address(input_fmap_7[71:64]),.clock  (clk));
logic signed [31:0] conv_mac_0;
logic signed [31:0] O0_N0_S0;		always @(posedge clk) O0_N0_S0 <=     O0_I0_R0_C0_SM1   +  O0_I0_R0_C1_SM1  ;
 logic signed [31:0] O0_N2_S0;		always @(posedge clk) O0_N2_S0 <=     O0_I0_R0_C2_SM1   +  O0_I0_R1_C0_SM1  ;
 logic signed [31:0] O0_N4_S0;		always @(posedge clk) O0_N4_S0 <=     O0_I0_R1_C1_SM1   +  O0_I0_R1_C2_SM1  ;
 logic signed [31:0] O0_N6_S0;		always @(posedge clk) O0_N6_S0 <=     O0_I0_R2_C0_SM1   +  O0_I0_R2_C1_SM1  ;
 logic signed [31:0] O0_N8_S0;		always @(posedge clk) O0_N8_S0 <=     O0_I0_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O0_N0_S1;		always @(posedge clk) O0_N0_S1 <=     O0_N0_S0  +  O0_N2_S0 ;
 logic signed [31:0] O0_N2_S1;		always @(posedge clk) O0_N2_S1 <=     O0_N4_S0  +  O0_N6_S0 ;
 logic signed [31:0] O0_N4_S1;		always @(posedge clk) O0_N4_S1 <=     O0_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O0_N0_S2;		always @(posedge clk) O0_N0_S2 <=     O0_N0_S1  +  O0_N2_S1 ;
 logic signed [31:0] O0_N2_S2;		always @(posedge clk) O0_N2_S2 <=     O0_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O0_N0_S3;		always @(posedge clk) O0_N0_S3 <=     O0_N0_S2  +  O0_N2_S2 ;
 assign conv_mac_0 = O0_N0_S3;

logic signed [31:0] conv_mac_1;
logic signed [31:0] O1_N0_S0;		always @(posedge clk) O1_N0_S0 <=     O1_I1_R0_C0_SM1   +  O1_I1_R0_C1_SM1  ;
 logic signed [31:0] O1_N2_S0;		always @(posedge clk) O1_N2_S0 <=     O1_I1_R0_C2_SM1   +  O1_I1_R1_C0_SM1  ;
 logic signed [31:0] O1_N4_S0;		always @(posedge clk) O1_N4_S0 <=     O1_I1_R1_C1_SM1   +  O1_I1_R1_C2_SM1  ;
 logic signed [31:0] O1_N6_S0;		always @(posedge clk) O1_N6_S0 <=     O1_I1_R2_C0_SM1   +  O1_I1_R2_C1_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O1_N0_S1;		always @(posedge clk) O1_N0_S1 <=     O1_N0_S0  +  O1_N2_S0 ;
 logic signed [31:0] O1_N2_S1;		always @(posedge clk) O1_N2_S1 <=     O1_N4_S0  +  O1_N6_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O1_N0_S2;		always @(posedge clk) O1_N0_S2 <=     O1_N0_S1  +  O1_N2_S1 ;
 assign conv_mac_1 = O1_N0_S2;

logic signed [31:0] conv_mac_2;
logic signed [31:0] O2_N0_S0;		always @(posedge clk) O2_N0_S0 <=     O2_I2_R0_C0_SM1   +  O2_I2_R0_C1_SM1  ;
 logic signed [31:0] O2_N2_S0;		always @(posedge clk) O2_N2_S0 <=     O2_I2_R0_C2_SM1   +  O2_I2_R1_C0_SM1  ;
 logic signed [31:0] O2_N4_S0;		always @(posedge clk) O2_N4_S0 <=     O2_I2_R1_C1_SM1   +  O2_I2_R1_C2_SM1  ;
 logic signed [31:0] O2_N6_S0;		always @(posedge clk) O2_N6_S0 <=     O2_I2_R2_C0_SM1   +  O2_I2_R2_C1_SM1  ;
 logic signed [31:0] O2_N8_S0;		always @(posedge clk) O2_N8_S0 <=     O2_I2_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O2_N0_S1;		always @(posedge clk) O2_N0_S1 <=     O2_N0_S0  +  O2_N2_S0 ;
 logic signed [31:0] O2_N2_S1;		always @(posedge clk) O2_N2_S1 <=     O2_N4_S0  +  O2_N6_S0 ;
 logic signed [31:0] O2_N4_S1;		always @(posedge clk) O2_N4_S1 <=     O2_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O2_N0_S2;		always @(posedge clk) O2_N0_S2 <=     O2_N0_S1  +  O2_N2_S1 ;
 logic signed [31:0] O2_N2_S2;		always @(posedge clk) O2_N2_S2 <=     O2_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O2_N0_S3;		always @(posedge clk) O2_N0_S3 <=     O2_N0_S2  +  O2_N2_S2 ;
 assign conv_mac_2 = O2_N0_S3;

logic signed [31:0] conv_mac_3;
logic signed [31:0] O3_N0_S0;		always @(posedge clk) O3_N0_S0 <=     O3_I3_R0_C0_SM1   +  O3_I3_R0_C1_SM1  ;
 logic signed [31:0] O3_N2_S0;		always @(posedge clk) O3_N2_S0 <=     O3_I3_R0_C2_SM1   +  O3_I3_R1_C0_SM1  ;
 logic signed [31:0] O3_N4_S0;		always @(posedge clk) O3_N4_S0 <=     O3_I3_R1_C1_SM1   +  O3_I3_R1_C2_SM1  ;
 logic signed [31:0] O3_N6_S0;		always @(posedge clk) O3_N6_S0 <=     O3_I3_R2_C0_SM1   +  O3_I3_R2_C1_SM1  ;
 logic signed [31:0] O3_N8_S0;		always @(posedge clk) O3_N8_S0 <=     O3_I3_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O3_N0_S1;		always @(posedge clk) O3_N0_S1 <=     O3_N0_S0  +  O3_N2_S0 ;
 logic signed [31:0] O3_N2_S1;		always @(posedge clk) O3_N2_S1 <=     O3_N4_S0  +  O3_N6_S0 ;
 logic signed [31:0] O3_N4_S1;		always @(posedge clk) O3_N4_S1 <=     O3_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O3_N0_S2;		always @(posedge clk) O3_N0_S2 <=     O3_N0_S1  +  O3_N2_S1 ;
 logic signed [31:0] O3_N2_S2;		always @(posedge clk) O3_N2_S2 <=     O3_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O3_N0_S3;		always @(posedge clk) O3_N0_S3 <=     O3_N0_S2  +  O3_N2_S2 ;
 assign conv_mac_3 = O3_N0_S3;

logic signed [31:0] conv_mac_4;
logic signed [31:0] O4_N0_S0;		always @(posedge clk) O4_N0_S0 <=     O4_I4_R0_C0_SM1   +  O4_I4_R0_C1_SM1  ;
 logic signed [31:0] O4_N2_S0;		always @(posedge clk) O4_N2_S0 <=     O4_I4_R0_C2_SM1   +  O4_I4_R1_C0_SM1  ;
 logic signed [31:0] O4_N4_S0;		always @(posedge clk) O4_N4_S0 <=     O4_I4_R1_C1_SM1   +  O4_I4_R1_C2_SM1  ;
 logic signed [31:0] O4_N6_S0;		always @(posedge clk) O4_N6_S0 <=     O4_I4_R2_C0_SM1   +  O4_I4_R2_C1_SM1  ;
 logic signed [31:0] O4_N8_S0;		always @(posedge clk) O4_N8_S0 <=     O4_I4_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O4_N0_S1;		always @(posedge clk) O4_N0_S1 <=     O4_N0_S0  +  O4_N2_S0 ;
 logic signed [31:0] O4_N2_S1;		always @(posedge clk) O4_N2_S1 <=     O4_N4_S0  +  O4_N6_S0 ;
 logic signed [31:0] O4_N4_S1;		always @(posedge clk) O4_N4_S1 <=     O4_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O4_N0_S2;		always @(posedge clk) O4_N0_S2 <=     O4_N0_S1  +  O4_N2_S1 ;
 logic signed [31:0] O4_N2_S2;		always @(posedge clk) O4_N2_S2 <=     O4_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O4_N0_S3;		always @(posedge clk) O4_N0_S3 <=     O4_N0_S2  +  O4_N2_S2 ;
 assign conv_mac_4 = O4_N0_S3;

logic signed [31:0] conv_mac_5;
logic signed [31:0] O5_N0_S0;		always @(posedge clk) O5_N0_S0 <=     O5_I5_R0_C0_SM1   +  O5_I5_R0_C1_SM1  ;
 logic signed [31:0] O5_N2_S0;		always @(posedge clk) O5_N2_S0 <=     O5_I5_R0_C2_SM1   +  O5_I5_R1_C0_SM1  ;
 logic signed [31:0] O5_N4_S0;		always @(posedge clk) O5_N4_S0 <=     O5_I5_R1_C1_SM1   +  O5_I5_R1_C2_SM1  ;
 logic signed [31:0] O5_N6_S0;		always @(posedge clk) O5_N6_S0 <=     O5_I5_R2_C0_SM1   +  O5_I5_R2_C1_SM1  ;
 logic signed [31:0] O5_N8_S0;		always @(posedge clk) O5_N8_S0 <=     O5_I5_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O5_N0_S1;		always @(posedge clk) O5_N0_S1 <=     O5_N0_S0  +  O5_N2_S0 ;
 logic signed [31:0] O5_N2_S1;		always @(posedge clk) O5_N2_S1 <=     O5_N4_S0  +  O5_N6_S0 ;
 logic signed [31:0] O5_N4_S1;		always @(posedge clk) O5_N4_S1 <=     O5_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O5_N0_S2;		always @(posedge clk) O5_N0_S2 <=     O5_N0_S1  +  O5_N2_S1 ;
 logic signed [31:0] O5_N2_S2;		always @(posedge clk) O5_N2_S2 <=     O5_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O5_N0_S3;		always @(posedge clk) O5_N0_S3 <=     O5_N0_S2  +  O5_N2_S2 ;
 assign conv_mac_5 = O5_N0_S3;

logic signed [31:0] conv_mac_6;
logic signed [31:0] O6_N0_S0;		always @(posedge clk) O6_N0_S0 <=     O6_I6_R0_C0_SM1   +  O6_I6_R0_C1_SM1  ;
 logic signed [31:0] O6_N2_S0;		always @(posedge clk) O6_N2_S0 <=     O6_I6_R0_C2_SM1   +  O6_I6_R1_C0_SM1  ;
 logic signed [31:0] O6_N4_S0;		always @(posedge clk) O6_N4_S0 <=     O6_I6_R1_C1_SM1   +  O6_I6_R1_C2_SM1  ;
 logic signed [31:0] O6_N6_S0;		always @(posedge clk) O6_N6_S0 <=     O6_I6_R2_C0_SM1   +  O6_I6_R2_C1_SM1  ;
 logic signed [31:0] O6_N8_S0;		always @(posedge clk) O6_N8_S0 <=     O6_I6_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O6_N0_S1;		always @(posedge clk) O6_N0_S1 <=     O6_N0_S0  +  O6_N2_S0 ;
 logic signed [31:0] O6_N2_S1;		always @(posedge clk) O6_N2_S1 <=     O6_N4_S0  +  O6_N6_S0 ;
 logic signed [31:0] O6_N4_S1;		always @(posedge clk) O6_N4_S1 <=     O6_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O6_N0_S2;		always @(posedge clk) O6_N0_S2 <=     O6_N0_S1  +  O6_N2_S1 ;
 logic signed [31:0] O6_N2_S2;		always @(posedge clk) O6_N2_S2 <=     O6_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O6_N0_S3;		always @(posedge clk) O6_N0_S3 <=     O6_N0_S2  +  O6_N2_S2 ;
 assign conv_mac_6 = O6_N0_S3;

logic signed [31:0] conv_mac_7;
logic signed [31:0] O7_N0_S0;		always @(posedge clk) O7_N0_S0 <=     O7_I7_R0_C0_SM1   +  O7_I7_R0_C1_SM1  ;
 logic signed [31:0] O7_N2_S0;		always @(posedge clk) O7_N2_S0 <=     O7_I7_R0_C2_SM1   +  O7_I7_R1_C0_SM1  ;
 logic signed [31:0] O7_N4_S0;		always @(posedge clk) O7_N4_S0 <=     O7_I7_R1_C1_SM1   +  O7_I7_R1_C2_SM1  ;
 logic signed [31:0] O7_N6_S0;		always @(posedge clk) O7_N6_S0 <=     O7_I7_R2_C0_SM1   +  O7_I7_R2_C1_SM1  ;
 logic signed [31:0] O7_N8_S0;		always @(posedge clk) O7_N8_S0 <=     O7_I7_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O7_N0_S1;		always @(posedge clk) O7_N0_S1 <=     O7_N0_S0  +  O7_N2_S0 ;
 logic signed [31:0] O7_N2_S1;		always @(posedge clk) O7_N2_S1 <=     O7_N4_S0  +  O7_N6_S0 ;
 logic signed [31:0] O7_N4_S1;		always @(posedge clk) O7_N4_S1 <=     O7_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O7_N0_S2;		always @(posedge clk) O7_N0_S2 <=     O7_N0_S1  +  O7_N2_S1 ;
 logic signed [31:0] O7_N2_S2;		always @(posedge clk) O7_N2_S2 <=     O7_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O7_N0_S3;		always @(posedge clk) O7_N0_S3 <=     O7_N0_S2  +  O7_N2_S2 ;
 assign conv_mac_7 = O7_N0_S3;

logic valid_D1;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D1<= 0 ;
	else valid_D1<=valid;
end
logic valid_D2;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D2<= 0 ;
	else valid_D2<=valid_D1;
end
logic valid_D3;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D3<= 0 ;
	else valid_D3<=valid_D2;
end
logic valid_D4;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D4<= 0 ;
	else valid_D4<=valid_D3;
end
logic valid_D5;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D5<= 0 ;
	else valid_D5<=valid_D4;
end
always_ff @(posedge clk) begin
	if (rstn == 0) ready <= 0 ;
	else ready <=valid_D5;
end
logic [31:0] bias_add_0;
assign bias_add_0 = conv_mac_0 + 5'd8;
logic [31:0] bias_add_1;
assign bias_add_1 = conv_mac_1 + 7'd44;
logic [31:0] bias_add_2;
assign bias_add_2 = conv_mac_2 - 5'd9;
logic [31:0] bias_add_3;
assign bias_add_3 = conv_mac_3 + 6'd25;
logic [31:0] bias_add_4;
assign bias_add_4 = conv_mac_4 + 7'd56;
logic [31:0] bias_add_5;
assign bias_add_5 = conv_mac_5 + 7'd47;
logic [31:0] bias_add_6;
assign bias_add_6 = conv_mac_6 + 8'd64;
logic [31:0] bias_add_7;
assign bias_add_7 = conv_mac_7 + 7'd35;

logic [7:0] relu_0;
assign relu_0[7:0] = (bias_add_0[31]==0) ? ((bias_add_0<3'd6) ? {{bias_add_0[31],bias_add_0[10:4]}} :'d6) : '0;
logic [7:0] relu_1;
assign relu_1[7:0] = (bias_add_1[31]==0) ? ((bias_add_1<3'd6) ? {{bias_add_1[31],bias_add_1[10:4]}} :'d6) : '0;
logic [7:0] relu_2;
assign relu_2[7:0] = (bias_add_2[31]==0) ? ((bias_add_2<3'd6) ? {{bias_add_2[31],bias_add_2[10:4]}} :'d6) : '0;
logic [7:0] relu_3;
assign relu_3[7:0] = (bias_add_3[31]==0) ? ((bias_add_3<3'd6) ? {{bias_add_3[31],bias_add_3[10:4]}} :'d6) : '0;
logic [7:0] relu_4;
assign relu_4[7:0] = (bias_add_4[31]==0) ? ((bias_add_4<3'd6) ? {{bias_add_4[31],bias_add_4[10:4]}} :'d6) : '0;
logic [7:0] relu_5;
assign relu_5[7:0] = (bias_add_5[31]==0) ? ((bias_add_5<3'd6) ? {{bias_add_5[31],bias_add_5[10:4]}} :'d6) : '0;
logic [7:0] relu_6;
assign relu_6[7:0] = (bias_add_6[31]==0) ? ((bias_add_6<3'd6) ? {{bias_add_6[31],bias_add_6[10:4]}} :'d6) : '0;
logic [7:0] relu_7;
assign relu_7[7:0] = (bias_add_7[31]==0) ? ((bias_add_7<3'd6) ? {{bias_add_7[31],bias_add_7[10:4]}} :'d6) : '0;

assign output_act = {
	relu_7,
	relu_6,
	relu_5,
	relu_4,
	relu_3,
	relu_2,
	relu_1,
	relu_0
};

endmodule
module conv3_dw (
    input logic clk,
    input logic rstn,
    input logic valid,
    input logic [16*72-1:0] input_act,
    output logic [128-1:0] output_act,
    output logic ready
);
logic we;
logic [8:0] zero_number; 
assign zero_number = 9'd0; 
logic [16*72-1:0] input_act_ff;
genvar i;
generate
for (i=0;i<16;i++)
    begin: genblk_8
        always_ff @(posedge clk) begin
            if (rstn == 0) begin
                input_act_ff[(i+1)*72-1:i*72] <= '0;
            end
            else begin
                input_act_ff[(i+1)*72-1:i*72] <= input_act[(i+1)*72-1:i*72];
            end
        end
    end
endgenerate
logic [71:0] input_fmap_0;
assign input_fmap_0 = input_act_ff[71:0];
logic [71:0] input_fmap_1;
assign input_fmap_1 = input_act_ff[143:72];
logic [71:0] input_fmap_2;
assign input_fmap_2 = input_act_ff[215:144];
logic [71:0] input_fmap_3;
assign input_fmap_3 = input_act_ff[287:216];
logic [71:0] input_fmap_4;
assign input_fmap_4 = input_act_ff[359:288];
logic [71:0] input_fmap_5;
assign input_fmap_5 = input_act_ff[431:360];
logic [71:0] input_fmap_6;
assign input_fmap_6 = input_act_ff[503:432];
logic [71:0] input_fmap_7;
assign input_fmap_7 = input_act_ff[575:504];
logic [71:0] input_fmap_8;
assign input_fmap_8 = input_act_ff[647:576];
logic [71:0] input_fmap_9;
assign input_fmap_9 = input_act_ff[719:648];
logic [71:0] input_fmap_10;
assign input_fmap_10 = input_act_ff[791:720];
logic [71:0] input_fmap_11;
assign input_fmap_11 = input_act_ff[863:792];
logic [71:0] input_fmap_12;
assign input_fmap_12 = input_act_ff[935:864];
logic [71:0] input_fmap_13;
assign input_fmap_13 = input_act_ff[1007:936];
logic [71:0] input_fmap_14;
assign input_fmap_14 = input_act_ff[1079:1008];
logic [71:0] input_fmap_15;
assign input_fmap_15 = input_act_ff[1151:1080];

logic [12-1:0] O0_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_dw_O0_I0_R0_C07_rom_inst (.q(O0_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O0_I0_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O0_I0_R0_C07_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_dw_O0_I0_R0_C07_rom_inst (.q(O0_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [12-1:0] O0_I0_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_dw_O0_I0_R0_C14_rom_inst (.q(O0_I0_R0_C1_SM1 ),.address(input_fmap_0[15:8]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R0_C1_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O0_I0_R0_C1_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O0_I0_R0_C14_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_dw_O0_I0_R0_C14_rom_inst (.q(O0_I0_R0_C1_SM1 ),.address(input_fmap_0[15:8]),.clock  (clk));
logic [12-1:0] O0_I0_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_dw_O0_I0_R0_C25_rom_inst (.q(O0_I0_R0_C2_SM1 ),.address(input_fmap_0[23:16]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R0_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O0_I0_R0_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O0_I0_R0_C25_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_dw_O0_I0_R0_C25_rom_inst (.q(O0_I0_R0_C2_SM1 ),.address(input_fmap_0[23:16]),.clock  (clk));
logic [11-1:0] O0_I0_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_dw_O0_I0_R1_C02_rom_inst (.q(O0_I0_R1_C0_SM1 ),.address(input_fmap_0[31:24]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R1_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O0_I0_R1_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O0_I0_R1_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_dw_O0_I0_R1_C02_rom_inst (.q(O0_I0_R1_C0_SM1 ),.address(input_fmap_0[31:24]),.clock  (clk));
logic [11-1:0] O0_I0_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_dw_O0_I0_R1_C12_rom_inst (.q(O0_I0_R1_C1_SM1 ),.address(input_fmap_0[39:32]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R1_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O0_I0_R1_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O0_I0_R1_C12_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_dw_O0_I0_R1_C12_rom_inst (.q(O0_I0_R1_C1_SM1 ),.address(input_fmap_0[39:32]),.clock  (clk));
logic [13-1:0] O0_I0_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv3_dw_O0_I0_R1_C213_rom_inst (.q(O0_I0_R1_C2_SM1 ),.address(input_fmap_0[47:40]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R1_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O0_I0_R1_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O0_I0_R1_C213_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv3_dw_O0_I0_R1_C213_rom_inst (.q(O0_I0_R1_C2_SM1 ),.address(input_fmap_0[47:40]),.clock  (clk));
logic [13-1:0] O0_I0_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv3_dw_O0_I0_R2_C09_rom_inst (.q(O0_I0_R2_C0_SM1 ),.address(input_fmap_0[55:48]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R2_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O0_I0_R2_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O0_I0_R2_C09_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv3_dw_O0_I0_R2_C09_rom_inst (.q(O0_I0_R2_C0_SM1 ),.address(input_fmap_0[55:48]),.clock  (clk));
logic [12-1:0] O0_I0_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_dw_O0_I0_R2_C14_rom_inst (.q(O0_I0_R2_C1_SM1 ),.address(input_fmap_0[63:56]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R2_C1_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O0_I0_R2_C1_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O0_I0_R2_C14_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_dw_O0_I0_R2_C14_rom_inst (.q(O0_I0_R2_C1_SM1 ),.address(input_fmap_0[63:56]),.clock  (clk));
logic [13-1:0] O0_I0_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv3_dw_O0_I0_R2_C29_rom_inst (.q(O0_I0_R2_C2_SM1 ),.address(input_fmap_0[71:64]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R2_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O0_I0_R2_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O0_I0_R2_C29_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv3_dw_O0_I0_R2_C29_rom_inst (.q(O0_I0_R2_C2_SM1 ),.address(input_fmap_0[71:64]),.clock  (clk));
logic [14-1:0] O1_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv3_dw_O1_I1_R0_C016_rom_inst (.q(O1_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R0_C0_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O1_I1_R0_C0_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O1_I1_R0_C016_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv3_dw_O1_I1_R0_C016_rom_inst (.q(O1_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [13-1:0] O1_I1_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv3_dw_O1_I1_R0_C114_rom_inst (.q(O1_I1_R0_C1_SM1 ),.address(input_fmap_1[15:8]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R0_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O1_I1_R0_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O1_I1_R0_C114_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv3_dw_O1_I1_R0_C114_rom_inst (.q(O1_I1_R0_C1_SM1 ),.address(input_fmap_1[15:8]),.clock  (clk));
logic [12-1:0] O1_I1_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_dw_O1_I1_R0_C24_rom_inst (.q(O1_I1_R0_C2_SM1 ),.address(input_fmap_1[23:16]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R0_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O1_I1_R0_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O1_I1_R0_C24_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_dw_O1_I1_R0_C24_rom_inst (.q(O1_I1_R0_C2_SM1 ),.address(input_fmap_1[23:16]),.clock  (clk));
logic [15-1:0] O1_I1_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(15),.INIT_FILE("deepfreeze_rom/deepfreeze_8_15.txt"))
    conv3_dw_O1_I1_R1_C045_rom_inst (.q(O1_I1_R1_C0_SM1 ),.address(input_fmap_1[31:24]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R1_C0_SM1  = 15'h1234;
//always@(posedge clk) begin 
//O1_I1_R1_C0_SM1  <= 15'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O1_I1_R1_C045_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(15))
//    conv3_dw_O1_I1_R1_C045_rom_inst (.q(O1_I1_R1_C0_SM1 ),.address(input_fmap_1[31:24]),.clock  (clk));
logic [14-1:0] O1_I1_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv3_dw_O1_I1_R1_C129_rom_inst (.q(O1_I1_R1_C1_SM1 ),.address(input_fmap_1[39:32]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R1_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O1_I1_R1_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O1_I1_R1_C129_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv3_dw_O1_I1_R1_C129_rom_inst (.q(O1_I1_R1_C1_SM1 ),.address(input_fmap_1[39:32]),.clock  (clk));
logic [13-1:0] O1_I1_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv3_dw_O1_I1_R1_C210_rom_inst (.q(O1_I1_R1_C2_SM1 ),.address(input_fmap_1[47:40]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R1_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O1_I1_R1_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O1_I1_R1_C210_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv3_dw_O1_I1_R1_C210_rom_inst (.q(O1_I1_R1_C2_SM1 ),.address(input_fmap_1[47:40]),.clock  (clk));
logic [15-1:0] O1_I1_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(15),.INIT_FILE("deepfreeze_rom/deepfreeze_8_15.txt"))
    conv3_dw_O1_I1_R2_C052_rom_inst (.q(O1_I1_R2_C0_SM1 ),.address(input_fmap_1[55:48]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R2_C0_SM1  = 15'h1234;
//always@(posedge clk) begin 
//O1_I1_R2_C0_SM1  <= 15'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O1_I1_R2_C052_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(15))
//    conv3_dw_O1_I1_R2_C052_rom_inst (.q(O1_I1_R2_C0_SM1 ),.address(input_fmap_1[55:48]),.clock  (clk));
logic [15-1:0] O1_I1_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(15),.INIT_FILE("deepfreeze_rom/deepfreeze_8_15.txt"))
    conv3_dw_O1_I1_R2_C142_rom_inst (.q(O1_I1_R2_C1_SM1 ),.address(input_fmap_1[63:56]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R2_C1_SM1  = 15'h1234;
//always@(posedge clk) begin 
//O1_I1_R2_C1_SM1  <= 15'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O1_I1_R2_C142_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(15))
//    conv3_dw_O1_I1_R2_C142_rom_inst (.q(O1_I1_R2_C1_SM1 ),.address(input_fmap_1[63:56]),.clock  (clk));
logic [13-1:0] O1_I1_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv3_dw_O1_I1_R2_C211_rom_inst (.q(O1_I1_R2_C2_SM1 ),.address(input_fmap_1[71:64]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R2_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O1_I1_R2_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O1_I1_R2_C211_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv3_dw_O1_I1_R2_C211_rom_inst (.q(O1_I1_R2_C2_SM1 ),.address(input_fmap_1[71:64]),.clock  (clk));
logic [14-1:0] O2_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv3_dw_O2_I2_R0_C024_rom_inst (.q(O2_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R0_C0_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O2_I2_R0_C0_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O2_I2_R0_C024_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv3_dw_O2_I2_R0_C024_rom_inst (.q(O2_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [14-1:0] O2_I2_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv3_dw_O2_I2_R0_C127_rom_inst (.q(O2_I2_R0_C1_SM1 ),.address(input_fmap_2[15:8]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R0_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O2_I2_R0_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O2_I2_R0_C127_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv3_dw_O2_I2_R0_C127_rom_inst (.q(O2_I2_R0_C1_SM1 ),.address(input_fmap_2[15:8]),.clock  (clk));
logic [12-1:0] O2_I2_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_dw_O2_I2_R0_C25_rom_inst (.q(O2_I2_R0_C2_SM1 ),.address(input_fmap_2[23:16]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R0_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O2_I2_R0_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O2_I2_R0_C25_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_dw_O2_I2_R0_C25_rom_inst (.q(O2_I2_R0_C2_SM1 ),.address(input_fmap_2[23:16]),.clock  (clk));
logic [14-1:0] O2_I2_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv3_dw_O2_I2_R1_C026_rom_inst (.q(O2_I2_R1_C0_SM1 ),.address(input_fmap_2[31:24]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R1_C0_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O2_I2_R1_C0_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O2_I2_R1_C026_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv3_dw_O2_I2_R1_C026_rom_inst (.q(O2_I2_R1_C0_SM1 ),.address(input_fmap_2[31:24]),.clock  (clk));
logic [15-1:0] O2_I2_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(15),.INIT_FILE("deepfreeze_rom/deepfreeze_8_15.txt"))
    conv3_dw_O2_I2_R1_C132_rom_inst (.q(O2_I2_R1_C1_SM1 ),.address(input_fmap_2[39:32]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R1_C1_SM1  = 15'h1234;
//always@(posedge clk) begin 
//O2_I2_R1_C1_SM1  <= 15'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O2_I2_R1_C132_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(15))
//    conv3_dw_O2_I2_R1_C132_rom_inst (.q(O2_I2_R1_C1_SM1 ),.address(input_fmap_2[39:32]),.clock  (clk));
logic [13-1:0] O2_I2_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv3_dw_O2_I2_R1_C29_rom_inst (.q(O2_I2_R1_C2_SM1 ),.address(input_fmap_2[47:40]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R1_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O2_I2_R1_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O2_I2_R1_C29_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv3_dw_O2_I2_R1_C29_rom_inst (.q(O2_I2_R1_C2_SM1 ),.address(input_fmap_2[47:40]),.clock  (clk));
logic [11-1:0] O2_I2_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_dw_O2_I2_R2_C02_rom_inst (.q(O2_I2_R2_C0_SM1 ),.address(input_fmap_2[55:48]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R2_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O2_I2_R2_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O2_I2_R2_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_dw_O2_I2_R2_C02_rom_inst (.q(O2_I2_R2_C0_SM1 ),.address(input_fmap_2[55:48]),.clock  (clk));
logic [12-1:0] O2_I2_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_dw_O2_I2_R2_C16_rom_inst (.q(O2_I2_R2_C1_SM1 ),.address(input_fmap_2[63:56]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R2_C1_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O2_I2_R2_C1_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O2_I2_R2_C16_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_dw_O2_I2_R2_C16_rom_inst (.q(O2_I2_R2_C1_SM1 ),.address(input_fmap_2[63:56]),.clock  (clk));
logic [12-1:0] O2_I2_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_dw_O2_I2_R2_C25_rom_inst (.q(O2_I2_R2_C2_SM1 ),.address(input_fmap_2[71:64]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R2_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O2_I2_R2_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O2_I2_R2_C25_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_dw_O2_I2_R2_C25_rom_inst (.q(O2_I2_R2_C2_SM1 ),.address(input_fmap_2[71:64]),.clock  (clk));
logic [11-1:0] O3_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_dw_O3_I3_R0_C02_rom_inst (.q(O3_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O3_I3_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O3_I3_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_dw_O3_I3_R0_C02_rom_inst (.q(O3_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [14-1:0] O3_I3_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv3_dw_O3_I3_R0_C127_rom_inst (.q(O3_I3_R0_C1_SM1 ),.address(input_fmap_3[15:8]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R0_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O3_I3_R0_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O3_I3_R0_C127_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv3_dw_O3_I3_R0_C127_rom_inst (.q(O3_I3_R0_C1_SM1 ),.address(input_fmap_3[15:8]),.clock  (clk));
logic [12-1:0] O3_I3_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_dw_O3_I3_R1_C05_rom_inst (.q(O3_I3_R1_C0_SM1 ),.address(input_fmap_3[31:24]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R1_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O3_I3_R1_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O3_I3_R1_C05_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_dw_O3_I3_R1_C05_rom_inst (.q(O3_I3_R1_C0_SM1 ),.address(input_fmap_3[31:24]),.clock  (clk));
logic [14-1:0] O3_I3_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv3_dw_O3_I3_R1_C126_rom_inst (.q(O3_I3_R1_C1_SM1 ),.address(input_fmap_3[39:32]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R1_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O3_I3_R1_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O3_I3_R1_C126_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv3_dw_O3_I3_R1_C126_rom_inst (.q(O3_I3_R1_C1_SM1 ),.address(input_fmap_3[39:32]),.clock  (clk));
logic [13-1:0] O3_I3_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv3_dw_O3_I3_R1_C210_rom_inst (.q(O3_I3_R1_C2_SM1 ),.address(input_fmap_3[47:40]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R1_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O3_I3_R1_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O3_I3_R1_C210_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv3_dw_O3_I3_R1_C210_rom_inst (.q(O3_I3_R1_C2_SM1 ),.address(input_fmap_3[47:40]),.clock  (clk));
logic [11-1:0] O3_I3_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_dw_O3_I3_R2_C03_rom_inst (.q(O3_I3_R2_C0_SM1 ),.address(input_fmap_3[55:48]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R2_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O3_I3_R2_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O3_I3_R2_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_dw_O3_I3_R2_C03_rom_inst (.q(O3_I3_R2_C0_SM1 ),.address(input_fmap_3[55:48]),.clock  (clk));
logic [12-1:0] O3_I3_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_dw_O3_I3_R2_C16_rom_inst (.q(O3_I3_R2_C1_SM1 ),.address(input_fmap_3[63:56]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R2_C1_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O3_I3_R2_C1_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O3_I3_R2_C16_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_dw_O3_I3_R2_C16_rom_inst (.q(O3_I3_R2_C1_SM1 ),.address(input_fmap_3[63:56]),.clock  (clk));
logic [12-1:0] O3_I3_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_dw_O3_I3_R2_C24_rom_inst (.q(O3_I3_R2_C2_SM1 ),.address(input_fmap_3[71:64]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R2_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O3_I3_R2_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O3_I3_R2_C24_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_dw_O3_I3_R2_C24_rom_inst (.q(O3_I3_R2_C2_SM1 ),.address(input_fmap_3[71:64]),.clock  (clk));
logic [13-1:0] O4_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv3_dw_O4_I4_R0_C08_rom_inst (.q(O4_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O4_I4_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O4_I4_R0_C08_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv3_dw_O4_I4_R0_C08_rom_inst (.q(O4_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [13-1:0] O4_I4_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv3_dw_O4_I4_R0_C111_rom_inst (.q(O4_I4_R0_C1_SM1 ),.address(input_fmap_4[15:8]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R0_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O4_I4_R0_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O4_I4_R0_C111_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv3_dw_O4_I4_R0_C111_rom_inst (.q(O4_I4_R0_C1_SM1 ),.address(input_fmap_4[15:8]),.clock  (clk));
logic [14-1:0] O4_I4_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv3_dw_O4_I4_R0_C216_rom_inst (.q(O4_I4_R0_C2_SM1 ),.address(input_fmap_4[23:16]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R0_C2_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O4_I4_R0_C2_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O4_I4_R0_C216_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv3_dw_O4_I4_R0_C216_rom_inst (.q(O4_I4_R0_C2_SM1 ),.address(input_fmap_4[23:16]),.clock  (clk));
logic [13-1:0] O4_I4_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv3_dw_O4_I4_R1_C012_rom_inst (.q(O4_I4_R1_C0_SM1 ),.address(input_fmap_4[31:24]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R1_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O4_I4_R1_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O4_I4_R1_C012_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv3_dw_O4_I4_R1_C012_rom_inst (.q(O4_I4_R1_C0_SM1 ),.address(input_fmap_4[31:24]),.clock  (clk));
logic [14-1:0] O4_I4_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv3_dw_O4_I4_R1_C117_rom_inst (.q(O4_I4_R1_C1_SM1 ),.address(input_fmap_4[39:32]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R1_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O4_I4_R1_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O4_I4_R1_C117_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv3_dw_O4_I4_R1_C117_rom_inst (.q(O4_I4_R1_C1_SM1 ),.address(input_fmap_4[39:32]),.clock  (clk));
logic [14-1:0] O4_I4_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv3_dw_O4_I4_R1_C222_rom_inst (.q(O4_I4_R1_C2_SM1 ),.address(input_fmap_4[47:40]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R1_C2_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O4_I4_R1_C2_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O4_I4_R1_C222_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv3_dw_O4_I4_R1_C222_rom_inst (.q(O4_I4_R1_C2_SM1 ),.address(input_fmap_4[47:40]),.clock  (clk));
logic [12-1:0] O4_I4_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_dw_O4_I4_R2_C14_rom_inst (.q(O4_I4_R2_C1_SM1 ),.address(input_fmap_4[63:56]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R2_C1_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O4_I4_R2_C1_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O4_I4_R2_C14_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_dw_O4_I4_R2_C14_rom_inst (.q(O4_I4_R2_C1_SM1 ),.address(input_fmap_4[63:56]),.clock  (clk));
logic [14-1:0] O5_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv3_dw_O5_I5_R0_C031_rom_inst (.q(O5_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R0_C0_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O5_I5_R0_C0_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O5_I5_R0_C031_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv3_dw_O5_I5_R0_C031_rom_inst (.q(O5_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [15-1:0] O5_I5_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(15),.INIT_FILE("deepfreeze_rom/deepfreeze_8_15.txt"))
    conv3_dw_O5_I5_R0_C141_rom_inst (.q(O5_I5_R0_C1_SM1 ),.address(input_fmap_5[15:8]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R0_C1_SM1  = 15'h1234;
//always@(posedge clk) begin 
//O5_I5_R0_C1_SM1  <= 15'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O5_I5_R0_C141_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(15))
//    conv3_dw_O5_I5_R0_C141_rom_inst (.q(O5_I5_R0_C1_SM1 ),.address(input_fmap_5[15:8]),.clock  (clk));
logic [14-1:0] O5_I5_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv3_dw_O5_I5_R0_C231_rom_inst (.q(O5_I5_R0_C2_SM1 ),.address(input_fmap_5[23:16]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R0_C2_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O5_I5_R0_C2_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O5_I5_R0_C231_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv3_dw_O5_I5_R0_C231_rom_inst (.q(O5_I5_R0_C2_SM1 ),.address(input_fmap_5[23:16]),.clock  (clk));
logic [10-1:0] O5_I5_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_dw_O5_I5_R1_C01_rom_inst (.q(O5_I5_R1_C0_SM1 ),.address(input_fmap_5[31:24]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R1_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I5_R1_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O5_I5_R1_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_dw_O5_I5_R1_C01_rom_inst (.q(O5_I5_R1_C0_SM1 ),.address(input_fmap_5[31:24]),.clock  (clk));
logic [10-1:0] O5_I5_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_dw_O5_I5_R1_C21_rom_inst (.q(O5_I5_R1_C2_SM1 ),.address(input_fmap_5[47:40]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R1_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I5_R1_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O5_I5_R1_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_dw_O5_I5_R1_C21_rom_inst (.q(O5_I5_R1_C2_SM1 ),.address(input_fmap_5[47:40]),.clock  (clk));
logic [13-1:0] O5_I5_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv3_dw_O5_I5_R2_C012_rom_inst (.q(O5_I5_R2_C0_SM1 ),.address(input_fmap_5[55:48]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R2_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O5_I5_R2_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O5_I5_R2_C012_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv3_dw_O5_I5_R2_C012_rom_inst (.q(O5_I5_R2_C0_SM1 ),.address(input_fmap_5[55:48]),.clock  (clk));
logic [13-1:0] O5_I5_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv3_dw_O5_I5_R2_C19_rom_inst (.q(O5_I5_R2_C1_SM1 ),.address(input_fmap_5[63:56]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R2_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O5_I5_R2_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O5_I5_R2_C19_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv3_dw_O5_I5_R2_C19_rom_inst (.q(O5_I5_R2_C1_SM1 ),.address(input_fmap_5[63:56]),.clock  (clk));
logic [12-1:0] O5_I5_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_dw_O5_I5_R2_C26_rom_inst (.q(O5_I5_R2_C2_SM1 ),.address(input_fmap_5[71:64]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R2_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O5_I5_R2_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O5_I5_R2_C26_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_dw_O5_I5_R2_C26_rom_inst (.q(O5_I5_R2_C2_SM1 ),.address(input_fmap_5[71:64]),.clock  (clk));
logic [15-1:0] O6_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(15),.INIT_FILE("deepfreeze_rom/deepfreeze_8_15.txt"))
    conv3_dw_O6_I6_R0_C040_rom_inst (.q(O6_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R0_C0_SM1  = 15'h1234;
//always@(posedge clk) begin 
//O6_I6_R0_C0_SM1  <= 15'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O6_I6_R0_C040_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(15))
//    conv3_dw_O6_I6_R0_C040_rom_inst (.q(O6_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [16-1:0] O6_I6_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(16),.INIT_FILE("deepfreeze_rom/deepfreeze_8_16.txt"))
    conv3_dw_O6_I6_R0_C177_rom_inst (.q(O6_I6_R0_C1_SM1 ),.address(input_fmap_6[15:8]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R0_C1_SM1  = 16'h1234;
//always@(posedge clk) begin 
//O6_I6_R0_C1_SM1  <= 16'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O6_I6_R0_C177_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(16))
//    conv3_dw_O6_I6_R0_C177_rom_inst (.q(O6_I6_R0_C1_SM1 ),.address(input_fmap_6[15:8]),.clock  (clk));
logic [15-1:0] O6_I6_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(15),.INIT_FILE("deepfreeze_rom/deepfreeze_8_15.txt"))
    conv3_dw_O6_I6_R0_C236_rom_inst (.q(O6_I6_R0_C2_SM1 ),.address(input_fmap_6[23:16]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R0_C2_SM1  = 15'h1234;
//always@(posedge clk) begin 
//O6_I6_R0_C2_SM1  <= 15'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O6_I6_R0_C236_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(15))
//    conv3_dw_O6_I6_R0_C236_rom_inst (.q(O6_I6_R0_C2_SM1 ),.address(input_fmap_6[23:16]),.clock  (clk));
logic [11-1:0] O6_I6_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_dw_O6_I6_R1_C02_rom_inst (.q(O6_I6_R1_C0_SM1 ),.address(input_fmap_6[31:24]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R1_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O6_I6_R1_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O6_I6_R1_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_dw_O6_I6_R1_C02_rom_inst (.q(O6_I6_R1_C0_SM1 ),.address(input_fmap_6[31:24]),.clock  (clk));
logic [12-1:0] O6_I6_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_dw_O6_I6_R1_C15_rom_inst (.q(O6_I6_R1_C1_SM1 ),.address(input_fmap_6[39:32]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R1_C1_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O6_I6_R1_C1_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O6_I6_R1_C15_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_dw_O6_I6_R1_C15_rom_inst (.q(O6_I6_R1_C1_SM1 ),.address(input_fmap_6[39:32]),.clock  (clk));
logic [14-1:0] O6_I6_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv3_dw_O6_I6_R1_C231_rom_inst (.q(O6_I6_R1_C2_SM1 ),.address(input_fmap_6[47:40]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R1_C2_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O6_I6_R1_C2_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O6_I6_R1_C231_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv3_dw_O6_I6_R1_C231_rom_inst (.q(O6_I6_R1_C2_SM1 ),.address(input_fmap_6[47:40]),.clock  (clk));
logic [13-1:0] O6_I6_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv3_dw_O6_I6_R2_C09_rom_inst (.q(O6_I6_R2_C0_SM1 ),.address(input_fmap_6[55:48]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R2_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O6_I6_R2_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O6_I6_R2_C09_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv3_dw_O6_I6_R2_C09_rom_inst (.q(O6_I6_R2_C0_SM1 ),.address(input_fmap_6[55:48]),.clock  (clk));
logic [14-1:0] O6_I6_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv3_dw_O6_I6_R2_C116_rom_inst (.q(O6_I6_R2_C1_SM1 ),.address(input_fmap_6[63:56]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R2_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O6_I6_R2_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O6_I6_R2_C116_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv3_dw_O6_I6_R2_C116_rom_inst (.q(O6_I6_R2_C1_SM1 ),.address(input_fmap_6[63:56]),.clock  (clk));
logic [12-1:0] O6_I6_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_dw_O6_I6_R2_C25_rom_inst (.q(O6_I6_R2_C2_SM1 ),.address(input_fmap_6[71:64]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R2_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O6_I6_R2_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O6_I6_R2_C25_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_dw_O6_I6_R2_C25_rom_inst (.q(O6_I6_R2_C2_SM1 ),.address(input_fmap_6[71:64]),.clock  (clk));
logic [11-1:0] O7_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_dw_O7_I7_R0_C02_rom_inst (.q(O7_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O7_I7_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O7_I7_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_dw_O7_I7_R0_C02_rom_inst (.q(O7_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [11-1:0] O7_I7_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_dw_O7_I7_R0_C12_rom_inst (.q(O7_I7_R0_C1_SM1 ),.address(input_fmap_7[15:8]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R0_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O7_I7_R0_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O7_I7_R0_C12_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_dw_O7_I7_R0_C12_rom_inst (.q(O7_I7_R0_C1_SM1 ),.address(input_fmap_7[15:8]),.clock  (clk));
logic [12-1:0] O7_I7_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_dw_O7_I7_R0_C26_rom_inst (.q(O7_I7_R0_C2_SM1 ),.address(input_fmap_7[23:16]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R0_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O7_I7_R0_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O7_I7_R0_C26_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_dw_O7_I7_R0_C26_rom_inst (.q(O7_I7_R0_C2_SM1 ),.address(input_fmap_7[23:16]),.clock  (clk));
logic [12-1:0] O7_I7_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_dw_O7_I7_R1_C05_rom_inst (.q(O7_I7_R1_C0_SM1 ),.address(input_fmap_7[31:24]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R1_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O7_I7_R1_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O7_I7_R1_C05_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_dw_O7_I7_R1_C05_rom_inst (.q(O7_I7_R1_C0_SM1 ),.address(input_fmap_7[31:24]),.clock  (clk));
logic [14-1:0] O7_I7_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv3_dw_O7_I7_R1_C124_rom_inst (.q(O7_I7_R1_C1_SM1 ),.address(input_fmap_7[39:32]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R1_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O7_I7_R1_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O7_I7_R1_C124_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv3_dw_O7_I7_R1_C124_rom_inst (.q(O7_I7_R1_C1_SM1 ),.address(input_fmap_7[39:32]),.clock  (clk));
logic [13-1:0] O7_I7_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv3_dw_O7_I7_R1_C214_rom_inst (.q(O7_I7_R1_C2_SM1 ),.address(input_fmap_7[47:40]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R1_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O7_I7_R1_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O7_I7_R1_C214_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv3_dw_O7_I7_R1_C214_rom_inst (.q(O7_I7_R1_C2_SM1 ),.address(input_fmap_7[47:40]),.clock  (clk));
logic [10-1:0] O7_I7_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_dw_O7_I7_R2_C01_rom_inst (.q(O7_I7_R2_C0_SM1 ),.address(input_fmap_7[55:48]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R2_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O7_I7_R2_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O7_I7_R2_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_dw_O7_I7_R2_C01_rom_inst (.q(O7_I7_R2_C0_SM1 ),.address(input_fmap_7[55:48]),.clock  (clk));
logic [13-1:0] O7_I7_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv3_dw_O7_I7_R2_C19_rom_inst (.q(O7_I7_R2_C1_SM1 ),.address(input_fmap_7[63:56]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R2_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O7_I7_R2_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O7_I7_R2_C19_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv3_dw_O7_I7_R2_C19_rom_inst (.q(O7_I7_R2_C1_SM1 ),.address(input_fmap_7[63:56]),.clock  (clk));
logic [12-1:0] O7_I7_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_dw_O7_I7_R2_C25_rom_inst (.q(O7_I7_R2_C2_SM1 ),.address(input_fmap_7[71:64]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R2_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O7_I7_R2_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O7_I7_R2_C25_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_dw_O7_I7_R2_C25_rom_inst (.q(O7_I7_R2_C2_SM1 ),.address(input_fmap_7[71:64]),.clock  (clk));
logic [13-1:0] O8_I8_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv3_dw_O8_I8_R0_C112_rom_inst (.q(O8_I8_R0_C1_SM1 ),.address(input_fmap_8[15:8]),.clk(clk),.d(0),.we(0));
//assign O8_I8_R0_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O8_I8_R0_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O8_I8_R0_C112_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv3_dw_O8_I8_R0_C112_rom_inst (.q(O8_I8_R0_C1_SM1 ),.address(input_fmap_8[15:8]),.clock  (clk));
logic [13-1:0] O8_I8_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv3_dw_O8_I8_R0_C213_rom_inst (.q(O8_I8_R0_C2_SM1 ),.address(input_fmap_8[23:16]),.clk(clk),.d(0),.we(0));
//assign O8_I8_R0_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O8_I8_R0_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O8_I8_R0_C213_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv3_dw_O8_I8_R0_C213_rom_inst (.q(O8_I8_R0_C2_SM1 ),.address(input_fmap_8[23:16]),.clock  (clk));
logic [13-1:0] O8_I8_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv3_dw_O8_I8_R1_C013_rom_inst (.q(O8_I8_R1_C0_SM1 ),.address(input_fmap_8[31:24]),.clk(clk),.d(0),.we(0));
//assign O8_I8_R1_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O8_I8_R1_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O8_I8_R1_C013_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv3_dw_O8_I8_R1_C013_rom_inst (.q(O8_I8_R1_C0_SM1 ),.address(input_fmap_8[31:24]),.clock  (clk));
logic [15-1:0] O8_I8_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(15),.INIT_FILE("deepfreeze_rom/deepfreeze_8_15.txt"))
    conv3_dw_O8_I8_R1_C133_rom_inst (.q(O8_I8_R1_C1_SM1 ),.address(input_fmap_8[39:32]),.clk(clk),.d(0),.we(0));
//assign O8_I8_R1_C1_SM1  = 15'h1234;
//always@(posedge clk) begin 
//O8_I8_R1_C1_SM1  <= 15'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O8_I8_R1_C133_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(15))
//    conv3_dw_O8_I8_R1_C133_rom_inst (.q(O8_I8_R1_C1_SM1 ),.address(input_fmap_8[39:32]),.clock  (clk));
logic [14-1:0] O8_I8_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv3_dw_O8_I8_R1_C226_rom_inst (.q(O8_I8_R1_C2_SM1 ),.address(input_fmap_8[47:40]),.clk(clk),.d(0),.we(0));
//assign O8_I8_R1_C2_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O8_I8_R1_C2_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O8_I8_R1_C226_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv3_dw_O8_I8_R1_C226_rom_inst (.q(O8_I8_R1_C2_SM1 ),.address(input_fmap_8[47:40]),.clock  (clk));
logic [12-1:0] O8_I8_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_dw_O8_I8_R2_C06_rom_inst (.q(O8_I8_R2_C0_SM1 ),.address(input_fmap_8[55:48]),.clk(clk),.d(0),.we(0));
//assign O8_I8_R2_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O8_I8_R2_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O8_I8_R2_C06_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_dw_O8_I8_R2_C06_rom_inst (.q(O8_I8_R2_C0_SM1 ),.address(input_fmap_8[55:48]),.clock  (clk));
logic [10-1:0] O8_I8_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_dw_O8_I8_R2_C11_rom_inst (.q(O8_I8_R2_C1_SM1 ),.address(input_fmap_8[63:56]),.clk(clk),.d(0),.we(0));
//assign O8_I8_R2_C1_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O8_I8_R2_C1_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O8_I8_R2_C11_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_dw_O8_I8_R2_C11_rom_inst (.q(O8_I8_R2_C1_SM1 ),.address(input_fmap_8[63:56]),.clock  (clk));
logic [10-1:0] O8_I8_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_dw_O8_I8_R2_C21_rom_inst (.q(O8_I8_R2_C2_SM1 ),.address(input_fmap_8[71:64]),.clk(clk),.d(0),.we(0));
//assign O8_I8_R2_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O8_I8_R2_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O8_I8_R2_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_dw_O8_I8_R2_C21_rom_inst (.q(O8_I8_R2_C2_SM1 ),.address(input_fmap_8[71:64]),.clock  (clk));
logic [11-1:0] O9_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_dw_O9_I9_R0_C03_rom_inst (.q(O9_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O9_I9_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O9_I9_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O9_I9_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_dw_O9_I9_R0_C03_rom_inst (.q(O9_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [13-1:0] O9_I9_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv3_dw_O9_I9_R0_C214_rom_inst (.q(O9_I9_R0_C2_SM1 ),.address(input_fmap_9[23:16]),.clk(clk),.d(0),.we(0));
//assign O9_I9_R0_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O9_I9_R0_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O9_I9_R0_C214_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv3_dw_O9_I9_R0_C214_rom_inst (.q(O9_I9_R0_C2_SM1 ),.address(input_fmap_9[23:16]),.clock  (clk));
logic [13-1:0] O9_I9_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv3_dw_O9_I9_R1_C09_rom_inst (.q(O9_I9_R1_C0_SM1 ),.address(input_fmap_9[31:24]),.clk(clk),.d(0),.we(0));
//assign O9_I9_R1_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O9_I9_R1_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O9_I9_R1_C09_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv3_dw_O9_I9_R1_C09_rom_inst (.q(O9_I9_R1_C0_SM1 ),.address(input_fmap_9[31:24]),.clock  (clk));
logic [15-1:0] O9_I9_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(15),.INIT_FILE("deepfreeze_rom/deepfreeze_8_15.txt"))
    conv3_dw_O9_I9_R1_C147_rom_inst (.q(O9_I9_R1_C1_SM1 ),.address(input_fmap_9[39:32]),.clk(clk),.d(0),.we(0));
//assign O9_I9_R1_C1_SM1  = 15'h1234;
//always@(posedge clk) begin 
//O9_I9_R1_C1_SM1  <= 15'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O9_I9_R1_C147_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(15))
//    conv3_dw_O9_I9_R1_C147_rom_inst (.q(O9_I9_R1_C1_SM1 ),.address(input_fmap_9[39:32]),.clock  (clk));
logic [13-1:0] O9_I9_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv3_dw_O9_I9_R1_C211_rom_inst (.q(O9_I9_R1_C2_SM1 ),.address(input_fmap_9[47:40]),.clk(clk),.d(0),.we(0));
//assign O9_I9_R1_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O9_I9_R1_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O9_I9_R1_C211_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv3_dw_O9_I9_R1_C211_rom_inst (.q(O9_I9_R1_C2_SM1 ),.address(input_fmap_9[47:40]),.clock  (clk));
logic [10-1:0] O9_I9_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_dw_O9_I9_R2_C01_rom_inst (.q(O9_I9_R2_C0_SM1 ),.address(input_fmap_9[55:48]),.clk(clk),.d(0),.we(0));
//assign O9_I9_R2_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O9_I9_R2_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O9_I9_R2_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_dw_O9_I9_R2_C01_rom_inst (.q(O9_I9_R2_C0_SM1 ),.address(input_fmap_9[55:48]),.clock  (clk));
logic [14-1:0] O9_I9_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv3_dw_O9_I9_R2_C117_rom_inst (.q(O9_I9_R2_C1_SM1 ),.address(input_fmap_9[63:56]),.clk(clk),.d(0),.we(0));
//assign O9_I9_R2_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O9_I9_R2_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O9_I9_R2_C117_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv3_dw_O9_I9_R2_C117_rom_inst (.q(O9_I9_R2_C1_SM1 ),.address(input_fmap_9[63:56]),.clock  (clk));
logic [11-1:0] O9_I9_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_dw_O9_I9_R2_C22_rom_inst (.q(O9_I9_R2_C2_SM1 ),.address(input_fmap_9[71:64]),.clk(clk),.d(0),.we(0));
//assign O9_I9_R2_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O9_I9_R2_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O9_I9_R2_C22_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_dw_O9_I9_R2_C22_rom_inst (.q(O9_I9_R2_C2_SM1 ),.address(input_fmap_9[71:64]),.clock  (clk));
logic [16-1:0] O10_I10_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(16),.INIT_FILE("deepfreeze_rom/deepfreeze_8_16.txt"))
    conv3_dw_O10_I10_R0_C067_rom_inst (.q(O10_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clk(clk),.d(0),.we(0));
//assign O10_I10_R0_C0_SM1  = 16'h1234;
//always@(posedge clk) begin 
//O10_I10_R0_C0_SM1  <= 16'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O10_I10_R0_C067_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(16))
//    conv3_dw_O10_I10_R0_C067_rom_inst (.q(O10_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clock  (clk));
logic [12-1:0] O10_I10_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_dw_O10_I10_R0_C15_rom_inst (.q(O10_I10_R0_C1_SM1 ),.address(input_fmap_10[15:8]),.clk(clk),.d(0),.we(0));
//assign O10_I10_R0_C1_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O10_I10_R0_C1_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O10_I10_R0_C15_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_dw_O10_I10_R0_C15_rom_inst (.q(O10_I10_R0_C1_SM1 ),.address(input_fmap_10[15:8]),.clock  (clk));
logic [14-1:0] O10_I10_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv3_dw_O10_I10_R0_C224_rom_inst (.q(O10_I10_R0_C2_SM1 ),.address(input_fmap_10[23:16]),.clk(clk),.d(0),.we(0));
//assign O10_I10_R0_C2_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O10_I10_R0_C2_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O10_I10_R0_C224_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv3_dw_O10_I10_R0_C224_rom_inst (.q(O10_I10_R0_C2_SM1 ),.address(input_fmap_10[23:16]),.clock  (clk));
logic [11-1:0] O10_I10_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_dw_O10_I10_R1_C02_rom_inst (.q(O10_I10_R1_C0_SM1 ),.address(input_fmap_10[31:24]),.clk(clk),.d(0),.we(0));
//assign O10_I10_R1_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O10_I10_R1_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O10_I10_R1_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_dw_O10_I10_R1_C02_rom_inst (.q(O10_I10_R1_C0_SM1 ),.address(input_fmap_10[31:24]),.clock  (clk));
logic [12-1:0] O10_I10_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_dw_O10_I10_R1_C14_rom_inst (.q(O10_I10_R1_C1_SM1 ),.address(input_fmap_10[39:32]),.clk(clk),.d(0),.we(0));
//assign O10_I10_R1_C1_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O10_I10_R1_C1_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O10_I10_R1_C14_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_dw_O10_I10_R1_C14_rom_inst (.q(O10_I10_R1_C1_SM1 ),.address(input_fmap_10[39:32]),.clock  (clk));
logic [11-1:0] O10_I10_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_dw_O10_I10_R1_C23_rom_inst (.q(O10_I10_R1_C2_SM1 ),.address(input_fmap_10[47:40]),.clk(clk),.d(0),.we(0));
//assign O10_I10_R1_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O10_I10_R1_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O10_I10_R1_C23_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_dw_O10_I10_R1_C23_rom_inst (.q(O10_I10_R1_C2_SM1 ),.address(input_fmap_10[47:40]),.clock  (clk));
logic [13-1:0] O10_I10_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv3_dw_O10_I10_R2_C08_rom_inst (.q(O10_I10_R2_C0_SM1 ),.address(input_fmap_10[55:48]),.clk(clk),.d(0),.we(0));
//assign O10_I10_R2_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O10_I10_R2_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O10_I10_R2_C08_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv3_dw_O10_I10_R2_C08_rom_inst (.q(O10_I10_R2_C0_SM1 ),.address(input_fmap_10[55:48]),.clock  (clk));
logic [10-1:0] O10_I10_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_dw_O10_I10_R2_C11_rom_inst (.q(O10_I10_R2_C1_SM1 ),.address(input_fmap_10[63:56]),.clk(clk),.d(0),.we(0));
//assign O10_I10_R2_C1_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O10_I10_R2_C1_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O10_I10_R2_C11_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_dw_O10_I10_R2_C11_rom_inst (.q(O10_I10_R2_C1_SM1 ),.address(input_fmap_10[63:56]),.clock  (clk));
logic [12-1:0] O10_I10_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_dw_O10_I10_R2_C26_rom_inst (.q(O10_I10_R2_C2_SM1 ),.address(input_fmap_10[71:64]),.clk(clk),.d(0),.we(0));
//assign O10_I10_R2_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O10_I10_R2_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O10_I10_R2_C26_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_dw_O10_I10_R2_C26_rom_inst (.q(O10_I10_R2_C2_SM1 ),.address(input_fmap_10[71:64]),.clock  (clk));
logic [12-1:0] O11_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_dw_O11_I11_R0_C05_rom_inst (.q(O11_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I11_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O11_I11_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O11_I11_R0_C05_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_dw_O11_I11_R0_C05_rom_inst (.q(O11_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [14-1:0] O11_I11_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv3_dw_O11_I11_R0_C124_rom_inst (.q(O11_I11_R0_C1_SM1 ),.address(input_fmap_11[15:8]),.clk(clk),.d(0),.we(0));
//assign O11_I11_R0_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O11_I11_R0_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O11_I11_R0_C124_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv3_dw_O11_I11_R0_C124_rom_inst (.q(O11_I11_R0_C1_SM1 ),.address(input_fmap_11[15:8]),.clock  (clk));
logic [14-1:0] O11_I11_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv3_dw_O11_I11_R0_C223_rom_inst (.q(O11_I11_R0_C2_SM1 ),.address(input_fmap_11[23:16]),.clk(clk),.d(0),.we(0));
//assign O11_I11_R0_C2_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O11_I11_R0_C2_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O11_I11_R0_C223_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv3_dw_O11_I11_R0_C223_rom_inst (.q(O11_I11_R0_C2_SM1 ),.address(input_fmap_11[23:16]),.clock  (clk));
logic [13-1:0] O11_I11_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv3_dw_O11_I11_R1_C08_rom_inst (.q(O11_I11_R1_C0_SM1 ),.address(input_fmap_11[31:24]),.clk(clk),.d(0),.we(0));
//assign O11_I11_R1_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O11_I11_R1_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O11_I11_R1_C08_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv3_dw_O11_I11_R1_C08_rom_inst (.q(O11_I11_R1_C0_SM1 ),.address(input_fmap_11[31:24]),.clock  (clk));
logic [14-1:0] O11_I11_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv3_dw_O11_I11_R1_C126_rom_inst (.q(O11_I11_R1_C1_SM1 ),.address(input_fmap_11[39:32]),.clk(clk),.d(0),.we(0));
//assign O11_I11_R1_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O11_I11_R1_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O11_I11_R1_C126_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv3_dw_O11_I11_R1_C126_rom_inst (.q(O11_I11_R1_C1_SM1 ),.address(input_fmap_11[39:32]),.clock  (clk));
logic [14-1:0] O11_I11_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv3_dw_O11_I11_R1_C227_rom_inst (.q(O11_I11_R1_C2_SM1 ),.address(input_fmap_11[47:40]),.clk(clk),.d(0),.we(0));
//assign O11_I11_R1_C2_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O11_I11_R1_C2_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O11_I11_R1_C227_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv3_dw_O11_I11_R1_C227_rom_inst (.q(O11_I11_R1_C2_SM1 ),.address(input_fmap_11[47:40]),.clock  (clk));
logic [10-1:0] O11_I11_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_dw_O11_I11_R2_C01_rom_inst (.q(O11_I11_R2_C0_SM1 ),.address(input_fmap_11[55:48]),.clk(clk),.d(0),.we(0));
//assign O11_I11_R2_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O11_I11_R2_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O11_I11_R2_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_dw_O11_I11_R2_C01_rom_inst (.q(O11_I11_R2_C0_SM1 ),.address(input_fmap_11[55:48]),.clock  (clk));
logic [10-1:0] O11_I11_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_dw_O11_I11_R2_C11_rom_inst (.q(O11_I11_R2_C1_SM1 ),.address(input_fmap_11[63:56]),.clk(clk),.d(0),.we(0));
//assign O11_I11_R2_C1_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O11_I11_R2_C1_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O11_I11_R2_C11_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_dw_O11_I11_R2_C11_rom_inst (.q(O11_I11_R2_C1_SM1 ),.address(input_fmap_11[63:56]),.clock  (clk));
logic [10-1:0] O11_I11_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_dw_O11_I11_R2_C21_rom_inst (.q(O11_I11_R2_C2_SM1 ),.address(input_fmap_11[71:64]),.clk(clk),.d(0),.we(0));
//assign O11_I11_R2_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O11_I11_R2_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O11_I11_R2_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_dw_O11_I11_R2_C21_rom_inst (.q(O11_I11_R2_C2_SM1 ),.address(input_fmap_11[71:64]),.clock  (clk));
logic [12-1:0] O12_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_dw_O12_I12_R0_C04_rom_inst (.q(O12_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I12_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O12_I12_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O12_I12_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_dw_O12_I12_R0_C04_rom_inst (.q(O12_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [14-1:0] O12_I12_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv3_dw_O12_I12_R0_C123_rom_inst (.q(O12_I12_R0_C1_SM1 ),.address(input_fmap_12[15:8]),.clk(clk),.d(0),.we(0));
//assign O12_I12_R0_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O12_I12_R0_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O12_I12_R0_C123_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv3_dw_O12_I12_R0_C123_rom_inst (.q(O12_I12_R0_C1_SM1 ),.address(input_fmap_12[15:8]),.clock  (clk));
logic [14-1:0] O12_I12_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv3_dw_O12_I12_R0_C216_rom_inst (.q(O12_I12_R0_C2_SM1 ),.address(input_fmap_12[23:16]),.clk(clk),.d(0),.we(0));
//assign O12_I12_R0_C2_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O12_I12_R0_C2_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O12_I12_R0_C216_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv3_dw_O12_I12_R0_C216_rom_inst (.q(O12_I12_R0_C2_SM1 ),.address(input_fmap_12[23:16]),.clock  (clk));
logic [13-1:0] O12_I12_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv3_dw_O12_I12_R1_C010_rom_inst (.q(O12_I12_R1_C0_SM1 ),.address(input_fmap_12[31:24]),.clk(clk),.d(0),.we(0));
//assign O12_I12_R1_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O12_I12_R1_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O12_I12_R1_C010_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv3_dw_O12_I12_R1_C010_rom_inst (.q(O12_I12_R1_C0_SM1 ),.address(input_fmap_12[31:24]),.clock  (clk));
logic [15-1:0] O12_I12_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(15),.INIT_FILE("deepfreeze_rom/deepfreeze_8_15.txt"))
    conv3_dw_O12_I12_R1_C133_rom_inst (.q(O12_I12_R1_C1_SM1 ),.address(input_fmap_12[39:32]),.clk(clk),.d(0),.we(0));
//assign O12_I12_R1_C1_SM1  = 15'h1234;
//always@(posedge clk) begin 
//O12_I12_R1_C1_SM1  <= 15'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O12_I12_R1_C133_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(15))
//    conv3_dw_O12_I12_R1_C133_rom_inst (.q(O12_I12_R1_C1_SM1 ),.address(input_fmap_12[39:32]),.clock  (clk));
logic [14-1:0] O12_I12_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv3_dw_O12_I12_R1_C227_rom_inst (.q(O12_I12_R1_C2_SM1 ),.address(input_fmap_12[47:40]),.clk(clk),.d(0),.we(0));
//assign O12_I12_R1_C2_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O12_I12_R1_C2_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O12_I12_R1_C227_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv3_dw_O12_I12_R1_C227_rom_inst (.q(O12_I12_R1_C2_SM1 ),.address(input_fmap_12[47:40]),.clock  (clk));
logic [13-1:0] O12_I12_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv3_dw_O12_I12_R2_C09_rom_inst (.q(O12_I12_R2_C0_SM1 ),.address(input_fmap_12[55:48]),.clk(clk),.d(0),.we(0));
//assign O12_I12_R2_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O12_I12_R2_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O12_I12_R2_C09_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv3_dw_O12_I12_R2_C09_rom_inst (.q(O12_I12_R2_C0_SM1 ),.address(input_fmap_12[55:48]),.clock  (clk));
logic [11-1:0] O12_I12_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_dw_O12_I12_R2_C12_rom_inst (.q(O12_I12_R2_C1_SM1 ),.address(input_fmap_12[63:56]),.clk(clk),.d(0),.we(0));
//assign O12_I12_R2_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O12_I12_R2_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O12_I12_R2_C12_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_dw_O12_I12_R2_C12_rom_inst (.q(O12_I12_R2_C1_SM1 ),.address(input_fmap_12[63:56]),.clock  (clk));
logic [13-1:0] O12_I12_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv3_dw_O12_I12_R2_C28_rom_inst (.q(O12_I12_R2_C2_SM1 ),.address(input_fmap_12[71:64]),.clk(clk),.d(0),.we(0));
//assign O12_I12_R2_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O12_I12_R2_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O12_I12_R2_C28_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv3_dw_O12_I12_R2_C28_rom_inst (.q(O12_I12_R2_C2_SM1 ),.address(input_fmap_12[71:64]),.clock  (clk));
logic [12-1:0] O13_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_dw_O13_I13_R0_C05_rom_inst (.q(O13_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O13_I13_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O13_I13_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O13_I13_R0_C05_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_dw_O13_I13_R0_C05_rom_inst (.q(O13_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [13-1:0] O13_I13_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv3_dw_O13_I13_R0_C113_rom_inst (.q(O13_I13_R0_C1_SM1 ),.address(input_fmap_13[15:8]),.clk(clk),.d(0),.we(0));
//assign O13_I13_R0_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O13_I13_R0_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O13_I13_R0_C113_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv3_dw_O13_I13_R0_C113_rom_inst (.q(O13_I13_R0_C1_SM1 ),.address(input_fmap_13[15:8]),.clock  (clk));
logic [11-1:0] O13_I13_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_dw_O13_I13_R0_C23_rom_inst (.q(O13_I13_R0_C2_SM1 ),.address(input_fmap_13[23:16]),.clk(clk),.d(0),.we(0));
//assign O13_I13_R0_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O13_I13_R0_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O13_I13_R0_C23_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_dw_O13_I13_R0_C23_rom_inst (.q(O13_I13_R0_C2_SM1 ),.address(input_fmap_13[23:16]),.clock  (clk));
logic [12-1:0] O13_I13_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_dw_O13_I13_R1_C04_rom_inst (.q(O13_I13_R1_C0_SM1 ),.address(input_fmap_13[31:24]),.clk(clk),.d(0),.we(0));
//assign O13_I13_R1_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O13_I13_R1_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O13_I13_R1_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_dw_O13_I13_R1_C04_rom_inst (.q(O13_I13_R1_C0_SM1 ),.address(input_fmap_13[31:24]),.clock  (clk));
logic [14-1:0] O13_I13_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv3_dw_O13_I13_R1_C125_rom_inst (.q(O13_I13_R1_C1_SM1 ),.address(input_fmap_13[39:32]),.clk(clk),.d(0),.we(0));
//assign O13_I13_R1_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O13_I13_R1_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O13_I13_R1_C125_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv3_dw_O13_I13_R1_C125_rom_inst (.q(O13_I13_R1_C1_SM1 ),.address(input_fmap_13[39:32]),.clock  (clk));
logic [13-1:0] O13_I13_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv3_dw_O13_I13_R1_C214_rom_inst (.q(O13_I13_R1_C2_SM1 ),.address(input_fmap_13[47:40]),.clk(clk),.d(0),.we(0));
//assign O13_I13_R1_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O13_I13_R1_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O13_I13_R1_C214_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv3_dw_O13_I13_R1_C214_rom_inst (.q(O13_I13_R1_C2_SM1 ),.address(input_fmap_13[47:40]),.clock  (clk));
logic [10-1:0] O13_I13_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_dw_O13_I13_R2_C01_rom_inst (.q(O13_I13_R2_C0_SM1 ),.address(input_fmap_13[55:48]),.clk(clk),.d(0),.we(0));
//assign O13_I13_R2_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O13_I13_R2_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O13_I13_R2_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_dw_O13_I13_R2_C01_rom_inst (.q(O13_I13_R2_C0_SM1 ),.address(input_fmap_13[55:48]),.clock  (clk));
logic [13-1:0] O13_I13_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv3_dw_O13_I13_R2_C115_rom_inst (.q(O13_I13_R2_C1_SM1 ),.address(input_fmap_13[63:56]),.clk(clk),.d(0),.we(0));
//assign O13_I13_R2_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O13_I13_R2_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O13_I13_R2_C115_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv3_dw_O13_I13_R2_C115_rom_inst (.q(O13_I13_R2_C1_SM1 ),.address(input_fmap_13[63:56]),.clock  (clk));
logic [12-1:0] O13_I13_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_dw_O13_I13_R2_C24_rom_inst (.q(O13_I13_R2_C2_SM1 ),.address(input_fmap_13[71:64]),.clk(clk),.d(0),.we(0));
//assign O13_I13_R2_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O13_I13_R2_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O13_I13_R2_C24_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_dw_O13_I13_R2_C24_rom_inst (.q(O13_I13_R2_C2_SM1 ),.address(input_fmap_13[71:64]),.clock  (clk));
logic [11-1:0] O14_I14_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_dw_O14_I14_R0_C02_rom_inst (.q(O14_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I14_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O14_I14_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O14_I14_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_dw_O14_I14_R0_C02_rom_inst (.q(O14_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clock  (clk));
logic [10-1:0] O14_I14_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_dw_O14_I14_R0_C11_rom_inst (.q(O14_I14_R0_C1_SM1 ),.address(input_fmap_14[15:8]),.clk(clk),.d(0),.we(0));
//assign O14_I14_R0_C1_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O14_I14_R0_C1_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O14_I14_R0_C11_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_dw_O14_I14_R0_C11_rom_inst (.q(O14_I14_R0_C1_SM1 ),.address(input_fmap_14[15:8]),.clock  (clk));
logic [12-1:0] O14_I14_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_dw_O14_I14_R0_C24_rom_inst (.q(O14_I14_R0_C2_SM1 ),.address(input_fmap_14[23:16]),.clk(clk),.d(0),.we(0));
//assign O14_I14_R0_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O14_I14_R0_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O14_I14_R0_C24_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_dw_O14_I14_R0_C24_rom_inst (.q(O14_I14_R0_C2_SM1 ),.address(input_fmap_14[23:16]),.clock  (clk));
logic [15-1:0] O14_I14_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(15),.INIT_FILE("deepfreeze_rom/deepfreeze_8_15.txt"))
    conv3_dw_O14_I14_R1_C134_rom_inst (.q(O14_I14_R1_C1_SM1 ),.address(input_fmap_14[39:32]),.clk(clk),.d(0),.we(0));
//assign O14_I14_R1_C1_SM1  = 15'h1234;
//always@(posedge clk) begin 
//O14_I14_R1_C1_SM1  <= 15'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O14_I14_R1_C134_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(15))
//    conv3_dw_O14_I14_R1_C134_rom_inst (.q(O14_I14_R1_C1_SM1 ),.address(input_fmap_14[39:32]),.clock  (clk));
logic [14-1:0] O14_I14_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv3_dw_O14_I14_R1_C220_rom_inst (.q(O14_I14_R1_C2_SM1 ),.address(input_fmap_14[47:40]),.clk(clk),.d(0),.we(0));
//assign O14_I14_R1_C2_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O14_I14_R1_C2_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O14_I14_R1_C220_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv3_dw_O14_I14_R1_C220_rom_inst (.q(O14_I14_R1_C2_SM1 ),.address(input_fmap_14[47:40]),.clock  (clk));
logic [11-1:0] O14_I14_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_dw_O14_I14_R2_C02_rom_inst (.q(O14_I14_R2_C0_SM1 ),.address(input_fmap_14[55:48]),.clk(clk),.d(0),.we(0));
//assign O14_I14_R2_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O14_I14_R2_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O14_I14_R2_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_dw_O14_I14_R2_C02_rom_inst (.q(O14_I14_R2_C0_SM1 ),.address(input_fmap_14[55:48]),.clock  (clk));
logic [13-1:0] O14_I14_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv3_dw_O14_I14_R2_C115_rom_inst (.q(O14_I14_R2_C1_SM1 ),.address(input_fmap_14[63:56]),.clk(clk),.d(0),.we(0));
//assign O14_I14_R2_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O14_I14_R2_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O14_I14_R2_C115_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv3_dw_O14_I14_R2_C115_rom_inst (.q(O14_I14_R2_C1_SM1 ),.address(input_fmap_14[63:56]),.clock  (clk));
logic [13-1:0] O14_I14_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv3_dw_O14_I14_R2_C28_rom_inst (.q(O14_I14_R2_C2_SM1 ),.address(input_fmap_14[71:64]),.clk(clk),.d(0),.we(0));
//assign O14_I14_R2_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O14_I14_R2_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O14_I14_R2_C28_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv3_dw_O14_I14_R2_C28_rom_inst (.q(O14_I14_R2_C2_SM1 ),.address(input_fmap_14[71:64]),.clock  (clk));
logic [13-1:0] O15_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv3_dw_O15_I15_R0_C013_rom_inst (.q(O15_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I15_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O15_I15_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O15_I15_R0_C013_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv3_dw_O15_I15_R0_C013_rom_inst (.q(O15_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [15-1:0] O15_I15_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(15),.INIT_FILE("deepfreeze_rom/deepfreeze_8_15.txt"))
    conv3_dw_O15_I15_R0_C132_rom_inst (.q(O15_I15_R0_C1_SM1 ),.address(input_fmap_15[15:8]),.clk(clk),.d(0),.we(0));
//assign O15_I15_R0_C1_SM1  = 15'h1234;
//always@(posedge clk) begin 
//O15_I15_R0_C1_SM1  <= 15'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O15_I15_R0_C132_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(15))
//    conv3_dw_O15_I15_R0_C132_rom_inst (.q(O15_I15_R0_C1_SM1 ),.address(input_fmap_15[15:8]),.clock  (clk));
logic [14-1:0] O15_I15_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv3_dw_O15_I15_R0_C222_rom_inst (.q(O15_I15_R0_C2_SM1 ),.address(input_fmap_15[23:16]),.clk(clk),.d(0),.we(0));
//assign O15_I15_R0_C2_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O15_I15_R0_C2_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O15_I15_R0_C222_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv3_dw_O15_I15_R0_C222_rom_inst (.q(O15_I15_R0_C2_SM1 ),.address(input_fmap_15[23:16]),.clock  (clk));
logic [13-1:0] O15_I15_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv3_dw_O15_I15_R1_C09_rom_inst (.q(O15_I15_R1_C0_SM1 ),.address(input_fmap_15[31:24]),.clk(clk),.d(0),.we(0));
//assign O15_I15_R1_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O15_I15_R1_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O15_I15_R1_C09_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv3_dw_O15_I15_R1_C09_rom_inst (.q(O15_I15_R1_C0_SM1 ),.address(input_fmap_15[31:24]),.clock  (clk));
logic [10-1:0] O15_I15_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_dw_O15_I15_R1_C11_rom_inst (.q(O15_I15_R1_C1_SM1 ),.address(input_fmap_15[39:32]),.clk(clk),.d(0),.we(0));
//assign O15_I15_R1_C1_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O15_I15_R1_C1_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O15_I15_R1_C11_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_dw_O15_I15_R1_C11_rom_inst (.q(O15_I15_R1_C1_SM1 ),.address(input_fmap_15[39:32]),.clock  (clk));
logic [15-1:0] O15_I15_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(15),.INIT_FILE("deepfreeze_rom/deepfreeze_8_15.txt"))
    conv3_dw_O15_I15_R1_C233_rom_inst (.q(O15_I15_R1_C2_SM1 ),.address(input_fmap_15[47:40]),.clk(clk),.d(0),.we(0));
//assign O15_I15_R1_C2_SM1  = 15'h1234;
//always@(posedge clk) begin 
//O15_I15_R1_C2_SM1  <= 15'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O15_I15_R1_C233_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(15))
//    conv3_dw_O15_I15_R1_C233_rom_inst (.q(O15_I15_R1_C2_SM1 ),.address(input_fmap_15[47:40]),.clock  (clk));
logic [10-1:0] O15_I15_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_dw_O15_I15_R2_C01_rom_inst (.q(O15_I15_R2_C0_SM1 ),.address(input_fmap_15[55:48]),.clk(clk),.d(0),.we(0));
//assign O15_I15_R2_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O15_I15_R2_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O15_I15_R2_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_dw_O15_I15_R2_C01_rom_inst (.q(O15_I15_R2_C0_SM1 ),.address(input_fmap_15[55:48]),.clock  (clk));
logic [10-1:0] O15_I15_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_dw_O15_I15_R2_C11_rom_inst (.q(O15_I15_R2_C1_SM1 ),.address(input_fmap_15[63:56]),.clk(clk),.d(0),.we(0));
//assign O15_I15_R2_C1_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O15_I15_R2_C1_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O15_I15_R2_C11_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_dw_O15_I15_R2_C11_rom_inst (.q(O15_I15_R2_C1_SM1 ),.address(input_fmap_15[63:56]),.clock  (clk));
logic [12-1:0] O15_I15_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_dw_O15_I15_R2_C25_rom_inst (.q(O15_I15_R2_C2_SM1 ),.address(input_fmap_15[71:64]),.clk(clk),.d(0),.we(0));
//assign O15_I15_R2_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O15_I15_R2_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_dw_O15_I15_R2_C25_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_dw_O15_I15_R2_C25_rom_inst (.q(O15_I15_R2_C2_SM1 ),.address(input_fmap_15[71:64]),.clock  (clk));
logic signed [31:0] conv_mac_0;
logic signed [31:0] O0_N0_S0;		always @(posedge clk) O0_N0_S0 <=     O0_I0_R0_C0_SM1   +  O0_I0_R0_C1_SM1  ;
 logic signed [31:0] O0_N2_S0;		always @(posedge clk) O0_N2_S0 <=     O0_I0_R0_C2_SM1   +  O0_I0_R1_C0_SM1  ;
 logic signed [31:0] O0_N4_S0;		always @(posedge clk) O0_N4_S0 <=     O0_I0_R1_C1_SM1   +  O0_I0_R1_C2_SM1  ;
 logic signed [31:0] O0_N6_S0;		always @(posedge clk) O0_N6_S0 <=     O0_I0_R2_C0_SM1   +  O0_I0_R2_C1_SM1  ;
 logic signed [31:0] O0_N8_S0;		always @(posedge clk) O0_N8_S0 <=     O0_I0_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O0_N0_S1;		always @(posedge clk) O0_N0_S1 <=     O0_N0_S0  +  O0_N2_S0 ;
 logic signed [31:0] O0_N2_S1;		always @(posedge clk) O0_N2_S1 <=     O0_N4_S0  +  O0_N6_S0 ;
 logic signed [31:0] O0_N4_S1;		always @(posedge clk) O0_N4_S1 <=     O0_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O0_N0_S2;		always @(posedge clk) O0_N0_S2 <=     O0_N0_S1  +  O0_N2_S1 ;
 logic signed [31:0] O0_N2_S2;		always @(posedge clk) O0_N2_S2 <=     O0_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O0_N0_S3;		always @(posedge clk) O0_N0_S3 <=     O0_N0_S2  +  O0_N2_S2 ;
 assign conv_mac_0 = O0_N0_S3;

logic signed [31:0] conv_mac_1;
logic signed [31:0] O1_N0_S0;		always @(posedge clk) O1_N0_S0 <=     O1_I1_R0_C0_SM1   +  O1_I1_R0_C1_SM1  ;
 logic signed [31:0] O1_N2_S0;		always @(posedge clk) O1_N2_S0 <=     O1_I1_R0_C2_SM1   +  O1_I1_R1_C0_SM1  ;
 logic signed [31:0] O1_N4_S0;		always @(posedge clk) O1_N4_S0 <=     O1_I1_R1_C1_SM1   +  O1_I1_R1_C2_SM1  ;
 logic signed [31:0] O1_N6_S0;		always @(posedge clk) O1_N6_S0 <=     O1_I1_R2_C0_SM1   +  O1_I1_R2_C1_SM1  ;
 logic signed [31:0] O1_N8_S0;		always @(posedge clk) O1_N8_S0 <=     O1_I1_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O1_N0_S1;		always @(posedge clk) O1_N0_S1 <=     O1_N0_S0  +  O1_N2_S0 ;
 logic signed [31:0] O1_N2_S1;		always @(posedge clk) O1_N2_S1 <=     O1_N4_S0  +  O1_N6_S0 ;
 logic signed [31:0] O1_N4_S1;		always @(posedge clk) O1_N4_S1 <=     O1_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O1_N0_S2;		always @(posedge clk) O1_N0_S2 <=     O1_N0_S1  +  O1_N2_S1 ;
 logic signed [31:0] O1_N2_S2;		always @(posedge clk) O1_N2_S2 <=     O1_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O1_N0_S3;		always @(posedge clk) O1_N0_S3 <=     O1_N0_S2  +  O1_N2_S2 ;
 assign conv_mac_1 = O1_N0_S3;

logic signed [31:0] conv_mac_2;
logic signed [31:0] O2_N0_S0;		always @(posedge clk) O2_N0_S0 <=     O2_I2_R0_C0_SM1   +  O2_I2_R0_C1_SM1  ;
 logic signed [31:0] O2_N2_S0;		always @(posedge clk) O2_N2_S0 <=     O2_I2_R0_C2_SM1   +  O2_I2_R1_C0_SM1  ;
 logic signed [31:0] O2_N4_S0;		always @(posedge clk) O2_N4_S0 <=     O2_I2_R1_C1_SM1   +  O2_I2_R1_C2_SM1  ;
 logic signed [31:0] O2_N6_S0;		always @(posedge clk) O2_N6_S0 <=     O2_I2_R2_C0_SM1   +  O2_I2_R2_C1_SM1  ;
 logic signed [31:0] O2_N8_S0;		always @(posedge clk) O2_N8_S0 <=     O2_I2_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O2_N0_S1;		always @(posedge clk) O2_N0_S1 <=     O2_N0_S0  +  O2_N2_S0 ;
 logic signed [31:0] O2_N2_S1;		always @(posedge clk) O2_N2_S1 <=     O2_N4_S0  +  O2_N6_S0 ;
 logic signed [31:0] O2_N4_S1;		always @(posedge clk) O2_N4_S1 <=     O2_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O2_N0_S2;		always @(posedge clk) O2_N0_S2 <=     O2_N0_S1  +  O2_N2_S1 ;
 logic signed [31:0] O2_N2_S2;		always @(posedge clk) O2_N2_S2 <=     O2_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O2_N0_S3;		always @(posedge clk) O2_N0_S3 <=     O2_N0_S2  +  O2_N2_S2 ;
 assign conv_mac_2 = O2_N0_S3;

logic signed [31:0] conv_mac_3;
logic signed [31:0] O3_N0_S0;		always @(posedge clk) O3_N0_S0 <=     O3_I3_R0_C0_SM1   +  O3_I3_R0_C1_SM1  ;
 logic signed [31:0] O3_N2_S0;		always @(posedge clk) O3_N2_S0 <=     O3_I3_R1_C0_SM1   +  O3_I3_R1_C1_SM1  ;
 logic signed [31:0] O3_N4_S0;		always @(posedge clk) O3_N4_S0 <=     O3_I3_R1_C2_SM1   +  O3_I3_R2_C0_SM1  ;
 logic signed [31:0] O3_N6_S0;		always @(posedge clk) O3_N6_S0 <=     O3_I3_R2_C1_SM1   +  O3_I3_R2_C2_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O3_N0_S1;		always @(posedge clk) O3_N0_S1 <=     O3_N0_S0  +  O3_N2_S0 ;
 logic signed [31:0] O3_N2_S1;		always @(posedge clk) O3_N2_S1 <=     O3_N4_S0  +  O3_N6_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O3_N0_S2;		always @(posedge clk) O3_N0_S2 <=     O3_N0_S1  +  O3_N2_S1 ;
 assign conv_mac_3 = O3_N0_S2;

logic signed [31:0] conv_mac_4;
logic signed [31:0] O4_N0_S0;		always @(posedge clk) O4_N0_S0 <=     O4_I4_R0_C0_SM1   +  O4_I4_R0_C1_SM1  ;
 logic signed [31:0] O4_N2_S0;		always @(posedge clk) O4_N2_S0 <=     O4_I4_R0_C2_SM1   +  O4_I4_R1_C0_SM1  ;
 logic signed [31:0] O4_N4_S0;		always @(posedge clk) O4_N4_S0 <=     O4_I4_R1_C1_SM1   +  O4_I4_R1_C2_SM1  ;
 logic signed [31:0] O4_N6_S0;		always @(posedge clk) O4_N6_S0 <=     O4_I4_R2_C1_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O4_N0_S1;		always @(posedge clk) O4_N0_S1 <=     O4_N0_S0  +  O4_N2_S0 ;
 logic signed [31:0] O4_N2_S1;		always @(posedge clk) O4_N2_S1 <=     O4_N4_S0  +  O4_N6_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O4_N0_S2;		always @(posedge clk) O4_N0_S2 <=     O4_N0_S1  +  O4_N2_S1 ;
 assign conv_mac_4 = O4_N0_S2;

logic signed [31:0] conv_mac_5;
logic signed [31:0] O5_N0_S0;		always @(posedge clk) O5_N0_S0 <=     O5_I5_R0_C0_SM1   +  O5_I5_R0_C1_SM1  ;
 logic signed [31:0] O5_N2_S0;		always @(posedge clk) O5_N2_S0 <=     O5_I5_R0_C2_SM1   +  O5_I5_R1_C0_SM1  ;
 logic signed [31:0] O5_N4_S0;		always @(posedge clk) O5_N4_S0 <=     O5_I5_R1_C2_SM1   +  O5_I5_R2_C0_SM1  ;
 logic signed [31:0] O5_N6_S0;		always @(posedge clk) O5_N6_S0 <=     O5_I5_R2_C1_SM1   +  O5_I5_R2_C2_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O5_N0_S1;		always @(posedge clk) O5_N0_S1 <=     O5_N0_S0  +  O5_N2_S0 ;
 logic signed [31:0] O5_N2_S1;		always @(posedge clk) O5_N2_S1 <=     O5_N4_S0  +  O5_N6_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O5_N0_S2;		always @(posedge clk) O5_N0_S2 <=     O5_N0_S1  +  O5_N2_S1 ;
 assign conv_mac_5 = O5_N0_S2;

logic signed [31:0] conv_mac_6;
logic signed [31:0] O6_N0_S0;		always @(posedge clk) O6_N0_S0 <=     O6_I6_R0_C0_SM1   +  O6_I6_R0_C1_SM1  ;
 logic signed [31:0] O6_N2_S0;		always @(posedge clk) O6_N2_S0 <=     O6_I6_R0_C2_SM1   +  O6_I6_R1_C0_SM1  ;
 logic signed [31:0] O6_N4_S0;		always @(posedge clk) O6_N4_S0 <=     O6_I6_R1_C1_SM1   +  O6_I6_R1_C2_SM1  ;
 logic signed [31:0] O6_N6_S0;		always @(posedge clk) O6_N6_S0 <=     O6_I6_R2_C0_SM1   +  O6_I6_R2_C1_SM1  ;
 logic signed [31:0] O6_N8_S0;		always @(posedge clk) O6_N8_S0 <=     O6_I6_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O6_N0_S1;		always @(posedge clk) O6_N0_S1 <=     O6_N0_S0  +  O6_N2_S0 ;
 logic signed [31:0] O6_N2_S1;		always @(posedge clk) O6_N2_S1 <=     O6_N4_S0  +  O6_N6_S0 ;
 logic signed [31:0] O6_N4_S1;		always @(posedge clk) O6_N4_S1 <=     O6_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O6_N0_S2;		always @(posedge clk) O6_N0_S2 <=     O6_N0_S1  +  O6_N2_S1 ;
 logic signed [31:0] O6_N2_S2;		always @(posedge clk) O6_N2_S2 <=     O6_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O6_N0_S3;		always @(posedge clk) O6_N0_S3 <=     O6_N0_S2  +  O6_N2_S2 ;
 assign conv_mac_6 = O6_N0_S3;

logic signed [31:0] conv_mac_7;
logic signed [31:0] O7_N0_S0;		always @(posedge clk) O7_N0_S0 <=     O7_I7_R0_C0_SM1   +  O7_I7_R0_C1_SM1  ;
 logic signed [31:0] O7_N2_S0;		always @(posedge clk) O7_N2_S0 <=     O7_I7_R0_C2_SM1   +  O7_I7_R1_C0_SM1  ;
 logic signed [31:0] O7_N4_S0;		always @(posedge clk) O7_N4_S0 <=     O7_I7_R1_C1_SM1   +  O7_I7_R1_C2_SM1  ;
 logic signed [31:0] O7_N6_S0;		always @(posedge clk) O7_N6_S0 <=     O7_I7_R2_C0_SM1   +  O7_I7_R2_C1_SM1  ;
 logic signed [31:0] O7_N8_S0;		always @(posedge clk) O7_N8_S0 <=     O7_I7_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O7_N0_S1;		always @(posedge clk) O7_N0_S1 <=     O7_N0_S0  +  O7_N2_S0 ;
 logic signed [31:0] O7_N2_S1;		always @(posedge clk) O7_N2_S1 <=     O7_N4_S0  +  O7_N6_S0 ;
 logic signed [31:0] O7_N4_S1;		always @(posedge clk) O7_N4_S1 <=     O7_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O7_N0_S2;		always @(posedge clk) O7_N0_S2 <=     O7_N0_S1  +  O7_N2_S1 ;
 logic signed [31:0] O7_N2_S2;		always @(posedge clk) O7_N2_S2 <=     O7_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O7_N0_S3;		always @(posedge clk) O7_N0_S3 <=     O7_N0_S2  +  O7_N2_S2 ;
 assign conv_mac_7 = O7_N0_S3;

logic signed [31:0] conv_mac_8;
logic signed [31:0] O8_N0_S0;		always @(posedge clk) O8_N0_S0 <=     O8_I8_R0_C1_SM1   +  O8_I8_R0_C2_SM1  ;
 logic signed [31:0] O8_N2_S0;		always @(posedge clk) O8_N2_S0 <=     O8_I8_R1_C0_SM1   +  O8_I8_R1_C1_SM1  ;
 logic signed [31:0] O8_N4_S0;		always @(posedge clk) O8_N4_S0 <=     O8_I8_R1_C2_SM1   +  O8_I8_R2_C0_SM1  ;
 logic signed [31:0] O8_N6_S0;		always @(posedge clk) O8_N6_S0 <=     O8_I8_R2_C1_SM1   +  O8_I8_R2_C2_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O8_N0_S1;		always @(posedge clk) O8_N0_S1 <=     O8_N0_S0  +  O8_N2_S0 ;
 logic signed [31:0] O8_N2_S1;		always @(posedge clk) O8_N2_S1 <=     O8_N4_S0  +  O8_N6_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O8_N0_S2;		always @(posedge clk) O8_N0_S2 <=     O8_N0_S1  +  O8_N2_S1 ;
 assign conv_mac_8 = O8_N0_S2;

logic signed [31:0] conv_mac_9;
logic signed [31:0] O9_N0_S0;		always @(posedge clk) O9_N0_S0 <=     O9_I9_R0_C0_SM1   +  O9_I9_R0_C2_SM1  ;
 logic signed [31:0] O9_N2_S0;		always @(posedge clk) O9_N2_S0 <=     O9_I9_R1_C0_SM1   +  O9_I9_R1_C1_SM1  ;
 logic signed [31:0] O9_N4_S0;		always @(posedge clk) O9_N4_S0 <=     O9_I9_R1_C2_SM1   +  O9_I9_R2_C0_SM1  ;
 logic signed [31:0] O9_N6_S0;		always @(posedge clk) O9_N6_S0 <=     O9_I9_R2_C1_SM1   +  O9_I9_R2_C2_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O9_N0_S1;		always @(posedge clk) O9_N0_S1 <=     O9_N0_S0  +  O9_N2_S0 ;
 logic signed [31:0] O9_N2_S1;		always @(posedge clk) O9_N2_S1 <=     O9_N4_S0  +  O9_N6_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O9_N0_S2;		always @(posedge clk) O9_N0_S2 <=     O9_N0_S1  +  O9_N2_S1 ;
 assign conv_mac_9 = O9_N0_S2;

logic signed [31:0] conv_mac_10;
logic signed [31:0] O10_N0_S0;		always @(posedge clk) O10_N0_S0 <=     O10_I10_R0_C0_SM1   +  O10_I10_R0_C1_SM1  ;
 logic signed [31:0] O10_N2_S0;		always @(posedge clk) O10_N2_S0 <=     O10_I10_R0_C2_SM1   +  O10_I10_R1_C0_SM1  ;
 logic signed [31:0] O10_N4_S0;		always @(posedge clk) O10_N4_S0 <=     O10_I10_R1_C1_SM1   +  O10_I10_R1_C2_SM1  ;
 logic signed [31:0] O10_N6_S0;		always @(posedge clk) O10_N6_S0 <=     O10_I10_R2_C0_SM1   +  O10_I10_R2_C1_SM1  ;
 logic signed [31:0] O10_N8_S0;		always @(posedge clk) O10_N8_S0 <=     O10_I10_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O10_N0_S1;		always @(posedge clk) O10_N0_S1 <=     O10_N0_S0  +  O10_N2_S0 ;
 logic signed [31:0] O10_N2_S1;		always @(posedge clk) O10_N2_S1 <=     O10_N4_S0  +  O10_N6_S0 ;
 logic signed [31:0] O10_N4_S1;		always @(posedge clk) O10_N4_S1 <=     O10_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O10_N0_S2;		always @(posedge clk) O10_N0_S2 <=     O10_N0_S1  +  O10_N2_S1 ;
 logic signed [31:0] O10_N2_S2;		always @(posedge clk) O10_N2_S2 <=     O10_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O10_N0_S3;		always @(posedge clk) O10_N0_S3 <=     O10_N0_S2  +  O10_N2_S2 ;
 assign conv_mac_10 = O10_N0_S3;

logic signed [31:0] conv_mac_11;
logic signed [31:0] O11_N0_S0;		always @(posedge clk) O11_N0_S0 <=     O11_I11_R0_C0_SM1   +  O11_I11_R0_C1_SM1  ;
 logic signed [31:0] O11_N2_S0;		always @(posedge clk) O11_N2_S0 <=     O11_I11_R0_C2_SM1   +  O11_I11_R1_C0_SM1  ;
 logic signed [31:0] O11_N4_S0;		always @(posedge clk) O11_N4_S0 <=     O11_I11_R1_C1_SM1   +  O11_I11_R1_C2_SM1  ;
 logic signed [31:0] O11_N6_S0;		always @(posedge clk) O11_N6_S0 <=     O11_I11_R2_C0_SM1   +  O11_I11_R2_C1_SM1  ;
 logic signed [31:0] O11_N8_S0;		always @(posedge clk) O11_N8_S0 <=     O11_I11_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O11_N0_S1;		always @(posedge clk) O11_N0_S1 <=     O11_N0_S0  +  O11_N2_S0 ;
 logic signed [31:0] O11_N2_S1;		always @(posedge clk) O11_N2_S1 <=     O11_N4_S0  +  O11_N6_S0 ;
 logic signed [31:0] O11_N4_S1;		always @(posedge clk) O11_N4_S1 <=     O11_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O11_N0_S2;		always @(posedge clk) O11_N0_S2 <=     O11_N0_S1  +  O11_N2_S1 ;
 logic signed [31:0] O11_N2_S2;		always @(posedge clk) O11_N2_S2 <=     O11_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O11_N0_S3;		always @(posedge clk) O11_N0_S3 <=     O11_N0_S2  +  O11_N2_S2 ;
 assign conv_mac_11 = O11_N0_S3;

logic signed [31:0] conv_mac_12;
logic signed [31:0] O12_N0_S0;		always @(posedge clk) O12_N0_S0 <=     O12_I12_R0_C0_SM1   +  O12_I12_R0_C1_SM1  ;
 logic signed [31:0] O12_N2_S0;		always @(posedge clk) O12_N2_S0 <=     O12_I12_R0_C2_SM1   +  O12_I12_R1_C0_SM1  ;
 logic signed [31:0] O12_N4_S0;		always @(posedge clk) O12_N4_S0 <=     O12_I12_R1_C1_SM1   +  O12_I12_R1_C2_SM1  ;
 logic signed [31:0] O12_N6_S0;		always @(posedge clk) O12_N6_S0 <=     O12_I12_R2_C0_SM1   +  O12_I12_R2_C1_SM1  ;
 logic signed [31:0] O12_N8_S0;		always @(posedge clk) O12_N8_S0 <=     O12_I12_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O12_N0_S1;		always @(posedge clk) O12_N0_S1 <=     O12_N0_S0  +  O12_N2_S0 ;
 logic signed [31:0] O12_N2_S1;		always @(posedge clk) O12_N2_S1 <=     O12_N4_S0  +  O12_N6_S0 ;
 logic signed [31:0] O12_N4_S1;		always @(posedge clk) O12_N4_S1 <=     O12_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O12_N0_S2;		always @(posedge clk) O12_N0_S2 <=     O12_N0_S1  +  O12_N2_S1 ;
 logic signed [31:0] O12_N2_S2;		always @(posedge clk) O12_N2_S2 <=     O12_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O12_N0_S3;		always @(posedge clk) O12_N0_S3 <=     O12_N0_S2  +  O12_N2_S2 ;
 assign conv_mac_12 = O12_N0_S3;

logic signed [31:0] conv_mac_13;
logic signed [31:0] O13_N0_S0;		always @(posedge clk) O13_N0_S0 <=     O13_I13_R0_C0_SM1   +  O13_I13_R0_C1_SM1  ;
 logic signed [31:0] O13_N2_S0;		always @(posedge clk) O13_N2_S0 <=     O13_I13_R0_C2_SM1   +  O13_I13_R1_C0_SM1  ;
 logic signed [31:0] O13_N4_S0;		always @(posedge clk) O13_N4_S0 <=     O13_I13_R1_C1_SM1   +  O13_I13_R1_C2_SM1  ;
 logic signed [31:0] O13_N6_S0;		always @(posedge clk) O13_N6_S0 <=     O13_I13_R2_C0_SM1   +  O13_I13_R2_C1_SM1  ;
 logic signed [31:0] O13_N8_S0;		always @(posedge clk) O13_N8_S0 <=     O13_I13_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O13_N0_S1;		always @(posedge clk) O13_N0_S1 <=     O13_N0_S0  +  O13_N2_S0 ;
 logic signed [31:0] O13_N2_S1;		always @(posedge clk) O13_N2_S1 <=     O13_N4_S0  +  O13_N6_S0 ;
 logic signed [31:0] O13_N4_S1;		always @(posedge clk) O13_N4_S1 <=     O13_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O13_N0_S2;		always @(posedge clk) O13_N0_S2 <=     O13_N0_S1  +  O13_N2_S1 ;
 logic signed [31:0] O13_N2_S2;		always @(posedge clk) O13_N2_S2 <=     O13_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O13_N0_S3;		always @(posedge clk) O13_N0_S3 <=     O13_N0_S2  +  O13_N2_S2 ;
 assign conv_mac_13 = O13_N0_S3;

logic signed [31:0] conv_mac_14;
logic signed [31:0] O14_N0_S0;		always @(posedge clk) O14_N0_S0 <=     O14_I14_R0_C0_SM1   +  O14_I14_R0_C1_SM1  ;
 logic signed [31:0] O14_N2_S0;		always @(posedge clk) O14_N2_S0 <=     O14_I14_R0_C2_SM1   +  O14_I14_R1_C1_SM1  ;
 logic signed [31:0] O14_N4_S0;		always @(posedge clk) O14_N4_S0 <=     O14_I14_R1_C2_SM1   +  O14_I14_R2_C0_SM1  ;
 logic signed [31:0] O14_N6_S0;		always @(posedge clk) O14_N6_S0 <=     O14_I14_R2_C1_SM1   +  O14_I14_R2_C2_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O14_N0_S1;		always @(posedge clk) O14_N0_S1 <=     O14_N0_S0  +  O14_N2_S0 ;
 logic signed [31:0] O14_N2_S1;		always @(posedge clk) O14_N2_S1 <=     O14_N4_S0  +  O14_N6_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O14_N0_S2;		always @(posedge clk) O14_N0_S2 <=     O14_N0_S1  +  O14_N2_S1 ;
 assign conv_mac_14 = O14_N0_S2;

logic signed [31:0] conv_mac_15;
logic signed [31:0] O15_N0_S0;		always @(posedge clk) O15_N0_S0 <=     O15_I15_R0_C0_SM1   +  O15_I15_R0_C1_SM1  ;
 logic signed [31:0] O15_N2_S0;		always @(posedge clk) O15_N2_S0 <=     O15_I15_R0_C2_SM1   +  O15_I15_R1_C0_SM1  ;
 logic signed [31:0] O15_N4_S0;		always @(posedge clk) O15_N4_S0 <=     O15_I15_R1_C1_SM1   +  O15_I15_R1_C2_SM1  ;
 logic signed [31:0] O15_N6_S0;		always @(posedge clk) O15_N6_S0 <=     O15_I15_R2_C0_SM1   +  O15_I15_R2_C1_SM1  ;
 logic signed [31:0] O15_N8_S0;		always @(posedge clk) O15_N8_S0 <=     O15_I15_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O15_N0_S1;		always @(posedge clk) O15_N0_S1 <=     O15_N0_S0  +  O15_N2_S0 ;
 logic signed [31:0] O15_N2_S1;		always @(posedge clk) O15_N2_S1 <=     O15_N4_S0  +  O15_N6_S0 ;
 logic signed [31:0] O15_N4_S1;		always @(posedge clk) O15_N4_S1 <=     O15_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O15_N0_S2;		always @(posedge clk) O15_N0_S2 <=     O15_N0_S1  +  O15_N2_S1 ;
 logic signed [31:0] O15_N2_S2;		always @(posedge clk) O15_N2_S2 <=     O15_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O15_N0_S3;		always @(posedge clk) O15_N0_S3 <=     O15_N0_S2  +  O15_N2_S2 ;
 assign conv_mac_15 = O15_N0_S3;

logic valid_D1;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D1<= 0 ;
	else valid_D1<=valid;
end
logic valid_D2;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D2<= 0 ;
	else valid_D2<=valid_D1;
end
logic valid_D3;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D3<= 0 ;
	else valid_D3<=valid_D2;
end
logic valid_D4;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D4<= 0 ;
	else valid_D4<=valid_D3;
end
logic valid_D5;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D5<= 0 ;
	else valid_D5<=valid_D4;
end
always_ff @(posedge clk) begin
	if (rstn == 0) ready <= 0 ;
	else ready <=valid_D5;
end
logic [31:0] bias_add_0;
assign bias_add_0 = conv_mac_0 + 6'd28;
logic [31:0] bias_add_1;
assign bias_add_1 = conv_mac_1 + 2'd1;
logic [31:0] bias_add_2;
assign bias_add_2 = conv_mac_2 + 3'd2;
logic [31:0] bias_add_3;
assign bias_add_3 = conv_mac_3 + 8'd67;
logic [31:0] bias_add_4;
assign bias_add_4 = conv_mac_4 + 6'd21;
logic [31:0] bias_add_5;
assign bias_add_5 = conv_mac_5 + 2'd1;
logic [31:0] bias_add_6;
assign bias_add_6 = conv_mac_6 + 7'd36;
logic [31:0] bias_add_7;
assign bias_add_7 = conv_mac_7 - 4'd4;
logic [31:0] bias_add_8;
assign bias_add_8 = conv_mac_8 + 6'd19;
logic [31:0] bias_add_9;
assign bias_add_9 = conv_mac_9 + 7'd58;
logic [31:0] bias_add_10;
assign bias_add_10 = conv_mac_10 + 5'd12;
logic [31:0] bias_add_11;
assign bias_add_11 = conv_mac_11 - 4'd4;
logic [31:0] bias_add_12;
assign bias_add_12 = conv_mac_12 - 2'd1;
logic [31:0] bias_add_13;
assign bias_add_13 = conv_mac_13 + 7'd32;
logic [31:0] bias_add_14;
assign bias_add_14 = conv_mac_14 + 6'd26;
logic [31:0] bias_add_15;
assign bias_add_15 = conv_mac_15 + 7'd52;

logic [7:0] relu_0;
assign relu_0[7:0] = (bias_add_0[31]==0) ? ((bias_add_0<3'd6) ? {{bias_add_0[31],bias_add_0[10:4]}} :'d6) : '0;
logic [7:0] relu_1;
assign relu_1[7:0] = (bias_add_1[31]==0) ? ((bias_add_1<3'd6) ? {{bias_add_1[31],bias_add_1[10:4]}} :'d6) : '0;
logic [7:0] relu_2;
assign relu_2[7:0] = (bias_add_2[31]==0) ? ((bias_add_2<3'd6) ? {{bias_add_2[31],bias_add_2[10:4]}} :'d6) : '0;
logic [7:0] relu_3;
assign relu_3[7:0] = (bias_add_3[31]==0) ? ((bias_add_3<3'd6) ? {{bias_add_3[31],bias_add_3[10:4]}} :'d6) : '0;
logic [7:0] relu_4;
assign relu_4[7:0] = (bias_add_4[31]==0) ? ((bias_add_4<3'd6) ? {{bias_add_4[31],bias_add_4[10:4]}} :'d6) : '0;
logic [7:0] relu_5;
assign relu_5[7:0] = (bias_add_5[31]==0) ? ((bias_add_5<3'd6) ? {{bias_add_5[31],bias_add_5[10:4]}} :'d6) : '0;
logic [7:0] relu_6;
assign relu_6[7:0] = (bias_add_6[31]==0) ? ((bias_add_6<3'd6) ? {{bias_add_6[31],bias_add_6[10:4]}} :'d6) : '0;
logic [7:0] relu_7;
assign relu_7[7:0] = (bias_add_7[31]==0) ? ((bias_add_7<3'd6) ? {{bias_add_7[31],bias_add_7[10:4]}} :'d6) : '0;
logic [7:0] relu_8;
assign relu_8[7:0] = (bias_add_8[31]==0) ? ((bias_add_8<3'd6) ? {{bias_add_8[31],bias_add_8[10:4]}} :'d6) : '0;
logic [7:0] relu_9;
assign relu_9[7:0] = (bias_add_9[31]==0) ? ((bias_add_9<3'd6) ? {{bias_add_9[31],bias_add_9[10:4]}} :'d6) : '0;
logic [7:0] relu_10;
assign relu_10[7:0] = (bias_add_10[31]==0) ? ((bias_add_10<3'd6) ? {{bias_add_10[31],bias_add_10[10:4]}} :'d6) : '0;
logic [7:0] relu_11;
assign relu_11[7:0] = (bias_add_11[31]==0) ? ((bias_add_11<3'd6) ? {{bias_add_11[31],bias_add_11[10:4]}} :'d6) : '0;
logic [7:0] relu_12;
assign relu_12[7:0] = (bias_add_12[31]==0) ? ((bias_add_12<3'd6) ? {{bias_add_12[31],bias_add_12[10:4]}} :'d6) : '0;
logic [7:0] relu_13;
assign relu_13[7:0] = (bias_add_13[31]==0) ? ((bias_add_13<3'd6) ? {{bias_add_13[31],bias_add_13[10:4]}} :'d6) : '0;
logic [7:0] relu_14;
assign relu_14[7:0] = (bias_add_14[31]==0) ? ((bias_add_14<3'd6) ? {{bias_add_14[31],bias_add_14[10:4]}} :'d6) : '0;
logic [7:0] relu_15;
assign relu_15[7:0] = (bias_add_15[31]==0) ? ((bias_add_15<3'd6) ? {{bias_add_15[31],bias_add_15[10:4]}} :'d6) : '0;

assign output_act = {
	relu_15,
	relu_14,
	relu_13,
	relu_12,
	relu_11,
	relu_10,
	relu_9,
	relu_8,
	relu_7,
	relu_6,
	relu_5,
	relu_4,
	relu_3,
	relu_2,
	relu_1,
	relu_0
};

endmodule
module conv4_dw (
    input logic clk,
    input logic rstn,
    input logic valid,
    input logic [16*72-1:0] input_act,
    output logic [128-1:0] output_act,
    output logic ready
);
logic we;
logic [8:0] zero_number; 
assign zero_number = 9'd0; 
logic [16*72-1:0] input_act_ff;
genvar i;
generate
for (i=0;i<16;i++)
    begin: genblk_9
        always_ff @(posedge clk) begin
            if (rstn == 0) begin
                input_act_ff[(i+1)*72-1:i*72] <= '0;
            end
            else begin
                input_act_ff[(i+1)*72-1:i*72] <= input_act[(i+1)*72-1:i*72];
            end
        end
    end
endgenerate
logic [71:0] input_fmap_0;
assign input_fmap_0 = input_act_ff[71:0];
logic [71:0] input_fmap_1;
assign input_fmap_1 = input_act_ff[143:72];
logic [71:0] input_fmap_2;
assign input_fmap_2 = input_act_ff[215:144];
logic [71:0] input_fmap_3;
assign input_fmap_3 = input_act_ff[287:216];
logic [71:0] input_fmap_4;
assign input_fmap_4 = input_act_ff[359:288];
logic [71:0] input_fmap_5;
assign input_fmap_5 = input_act_ff[431:360];
logic [71:0] input_fmap_6;
assign input_fmap_6 = input_act_ff[503:432];
logic [71:0] input_fmap_7;
assign input_fmap_7 = input_act_ff[575:504];
logic [71:0] input_fmap_8;
assign input_fmap_8 = input_act_ff[647:576];
logic [71:0] input_fmap_9;
assign input_fmap_9 = input_act_ff[719:648];
logic [71:0] input_fmap_10;
assign input_fmap_10 = input_act_ff[791:720];
logic [71:0] input_fmap_11;
assign input_fmap_11 = input_act_ff[863:792];
logic [71:0] input_fmap_12;
assign input_fmap_12 = input_act_ff[935:864];
logic [71:0] input_fmap_13;
assign input_fmap_13 = input_act_ff[1007:936];
logic [71:0] input_fmap_14;
assign input_fmap_14 = input_act_ff[1079:1008];
logic [71:0] input_fmap_15;
assign input_fmap_15 = input_act_ff[1151:1080];

logic [13-1:0] O0_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O0_I0_R0_C010_rom_inst (.q(O0_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O0_I0_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O0_I0_R0_C010_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O0_I0_R0_C010_rom_inst (.q(O0_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [13-1:0] O0_I0_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O0_I0_R0_C110_rom_inst (.q(O0_I0_R0_C1_SM1 ),.address(input_fmap_0[15:8]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R0_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O0_I0_R0_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O0_I0_R0_C110_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O0_I0_R0_C110_rom_inst (.q(O0_I0_R0_C1_SM1 ),.address(input_fmap_0[15:8]),.clock  (clk));
logic [11-1:0] O0_I0_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_dw_O0_I0_R0_C22_rom_inst (.q(O0_I0_R0_C2_SM1 ),.address(input_fmap_0[23:16]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R0_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O0_I0_R0_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O0_I0_R0_C22_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_dw_O0_I0_R0_C22_rom_inst (.q(O0_I0_R0_C2_SM1 ),.address(input_fmap_0[23:16]),.clock  (clk));
logic [14-1:0] O0_I0_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv4_dw_O0_I0_R1_C016_rom_inst (.q(O0_I0_R1_C0_SM1 ),.address(input_fmap_0[31:24]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R1_C0_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O0_I0_R1_C0_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O0_I0_R1_C016_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv4_dw_O0_I0_R1_C016_rom_inst (.q(O0_I0_R1_C0_SM1 ),.address(input_fmap_0[31:24]),.clock  (clk));
logic [14-1:0] O0_I0_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv4_dw_O0_I0_R1_C119_rom_inst (.q(O0_I0_R1_C1_SM1 ),.address(input_fmap_0[39:32]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R1_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O0_I0_R1_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O0_I0_R1_C119_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv4_dw_O0_I0_R1_C119_rom_inst (.q(O0_I0_R1_C1_SM1 ),.address(input_fmap_0[39:32]),.clock  (clk));
logic [13-1:0] O0_I0_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O0_I0_R1_C28_rom_inst (.q(O0_I0_R1_C2_SM1 ),.address(input_fmap_0[47:40]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R1_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O0_I0_R1_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O0_I0_R1_C28_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O0_I0_R1_C28_rom_inst (.q(O0_I0_R1_C2_SM1 ),.address(input_fmap_0[47:40]),.clock  (clk));
logic [12-1:0] O0_I0_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_dw_O0_I0_R2_C07_rom_inst (.q(O0_I0_R2_C0_SM1 ),.address(input_fmap_0[55:48]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R2_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O0_I0_R2_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O0_I0_R2_C07_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_dw_O0_I0_R2_C07_rom_inst (.q(O0_I0_R2_C0_SM1 ),.address(input_fmap_0[55:48]),.clock  (clk));
logic [13-1:0] O0_I0_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O0_I0_R2_C110_rom_inst (.q(O0_I0_R2_C1_SM1 ),.address(input_fmap_0[63:56]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R2_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O0_I0_R2_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O0_I0_R2_C110_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O0_I0_R2_C110_rom_inst (.q(O0_I0_R2_C1_SM1 ),.address(input_fmap_0[63:56]),.clock  (clk));
logic [12-1:0] O0_I0_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_dw_O0_I0_R2_C25_rom_inst (.q(O0_I0_R2_C2_SM1 ),.address(input_fmap_0[71:64]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R2_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O0_I0_R2_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O0_I0_R2_C25_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_dw_O0_I0_R2_C25_rom_inst (.q(O0_I0_R2_C2_SM1 ),.address(input_fmap_0[71:64]),.clock  (clk));
logic [12-1:0] O1_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_dw_O1_I1_R0_C06_rom_inst (.q(O1_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O1_I1_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O1_I1_R0_C06_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_dw_O1_I1_R0_C06_rom_inst (.q(O1_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [13-1:0] O1_I1_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O1_I1_R0_C114_rom_inst (.q(O1_I1_R0_C1_SM1 ),.address(input_fmap_1[15:8]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R0_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O1_I1_R0_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O1_I1_R0_C114_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O1_I1_R0_C114_rom_inst (.q(O1_I1_R0_C1_SM1 ),.address(input_fmap_1[15:8]),.clock  (clk));
logic [13-1:0] O1_I1_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O1_I1_R0_C28_rom_inst (.q(O1_I1_R0_C2_SM1 ),.address(input_fmap_1[23:16]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R0_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O1_I1_R0_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O1_I1_R0_C28_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O1_I1_R0_C28_rom_inst (.q(O1_I1_R0_C2_SM1 ),.address(input_fmap_1[23:16]),.clock  (clk));
logic [13-1:0] O1_I1_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O1_I1_R1_C08_rom_inst (.q(O1_I1_R1_C0_SM1 ),.address(input_fmap_1[31:24]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R1_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O1_I1_R1_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O1_I1_R1_C08_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O1_I1_R1_C08_rom_inst (.q(O1_I1_R1_C0_SM1 ),.address(input_fmap_1[31:24]),.clock  (clk));
logic [14-1:0] O1_I1_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv4_dw_O1_I1_R1_C121_rom_inst (.q(O1_I1_R1_C1_SM1 ),.address(input_fmap_1[39:32]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R1_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O1_I1_R1_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O1_I1_R1_C121_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv4_dw_O1_I1_R1_C121_rom_inst (.q(O1_I1_R1_C1_SM1 ),.address(input_fmap_1[39:32]),.clock  (clk));
logic [13-1:0] O1_I1_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O1_I1_R1_C213_rom_inst (.q(O1_I1_R1_C2_SM1 ),.address(input_fmap_1[47:40]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R1_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O1_I1_R1_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O1_I1_R1_C213_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O1_I1_R1_C213_rom_inst (.q(O1_I1_R1_C2_SM1 ),.address(input_fmap_1[47:40]),.clock  (clk));
logic [12-1:0] O1_I1_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_dw_O1_I1_R2_C04_rom_inst (.q(O1_I1_R2_C0_SM1 ),.address(input_fmap_1[55:48]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R2_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O1_I1_R2_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O1_I1_R2_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_dw_O1_I1_R2_C04_rom_inst (.q(O1_I1_R2_C0_SM1 ),.address(input_fmap_1[55:48]),.clock  (clk));
logic [13-1:0] O1_I1_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O1_I1_R2_C19_rom_inst (.q(O1_I1_R2_C1_SM1 ),.address(input_fmap_1[63:56]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R2_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O1_I1_R2_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O1_I1_R2_C19_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O1_I1_R2_C19_rom_inst (.q(O1_I1_R2_C1_SM1 ),.address(input_fmap_1[63:56]),.clock  (clk));
logic [12-1:0] O1_I1_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_dw_O1_I1_R2_C26_rom_inst (.q(O1_I1_R2_C2_SM1 ),.address(input_fmap_1[71:64]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R2_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O1_I1_R2_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O1_I1_R2_C26_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_dw_O1_I1_R2_C26_rom_inst (.q(O1_I1_R2_C2_SM1 ),.address(input_fmap_1[71:64]),.clock  (clk));
logic [13-1:0] O2_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O2_I2_R0_C011_rom_inst (.q(O2_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O2_I2_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O2_I2_R0_C011_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O2_I2_R0_C011_rom_inst (.q(O2_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [13-1:0] O2_I2_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O2_I2_R0_C115_rom_inst (.q(O2_I2_R0_C1_SM1 ),.address(input_fmap_2[15:8]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R0_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O2_I2_R0_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O2_I2_R0_C115_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O2_I2_R0_C115_rom_inst (.q(O2_I2_R0_C1_SM1 ),.address(input_fmap_2[15:8]),.clock  (clk));
logic [12-1:0] O2_I2_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_dw_O2_I2_R0_C26_rom_inst (.q(O2_I2_R0_C2_SM1 ),.address(input_fmap_2[23:16]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R0_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O2_I2_R0_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O2_I2_R0_C26_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_dw_O2_I2_R0_C26_rom_inst (.q(O2_I2_R0_C2_SM1 ),.address(input_fmap_2[23:16]),.clock  (clk));
logic [13-1:0] O2_I2_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O2_I2_R1_C010_rom_inst (.q(O2_I2_R1_C0_SM1 ),.address(input_fmap_2[31:24]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R1_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O2_I2_R1_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O2_I2_R1_C010_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O2_I2_R1_C010_rom_inst (.q(O2_I2_R1_C0_SM1 ),.address(input_fmap_2[31:24]),.clock  (clk));
logic [14-1:0] O2_I2_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv4_dw_O2_I2_R1_C119_rom_inst (.q(O2_I2_R1_C1_SM1 ),.address(input_fmap_2[39:32]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R1_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O2_I2_R1_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O2_I2_R1_C119_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv4_dw_O2_I2_R1_C119_rom_inst (.q(O2_I2_R1_C1_SM1 ),.address(input_fmap_2[39:32]),.clock  (clk));
logic [13-1:0] O2_I2_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O2_I2_R1_C210_rom_inst (.q(O2_I2_R1_C2_SM1 ),.address(input_fmap_2[47:40]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R1_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O2_I2_R1_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O2_I2_R1_C210_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O2_I2_R1_C210_rom_inst (.q(O2_I2_R1_C2_SM1 ),.address(input_fmap_2[47:40]),.clock  (clk));
logic [11-1:0] O2_I2_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_dw_O2_I2_R2_C03_rom_inst (.q(O2_I2_R2_C0_SM1 ),.address(input_fmap_2[55:48]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R2_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O2_I2_R2_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O2_I2_R2_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_dw_O2_I2_R2_C03_rom_inst (.q(O2_I2_R2_C0_SM1 ),.address(input_fmap_2[55:48]),.clock  (clk));
logic [12-1:0] O2_I2_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_dw_O2_I2_R2_C17_rom_inst (.q(O2_I2_R2_C1_SM1 ),.address(input_fmap_2[63:56]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R2_C1_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O2_I2_R2_C1_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O2_I2_R2_C17_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_dw_O2_I2_R2_C17_rom_inst (.q(O2_I2_R2_C1_SM1 ),.address(input_fmap_2[63:56]),.clock  (clk));
logic [12-1:0] O2_I2_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_dw_O2_I2_R2_C25_rom_inst (.q(O2_I2_R2_C2_SM1 ),.address(input_fmap_2[71:64]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R2_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O2_I2_R2_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O2_I2_R2_C25_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_dw_O2_I2_R2_C25_rom_inst (.q(O2_I2_R2_C2_SM1 ),.address(input_fmap_2[71:64]),.clock  (clk));
logic [13-1:0] O3_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O3_I3_R0_C08_rom_inst (.q(O3_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O3_I3_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O3_I3_R0_C08_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O3_I3_R0_C08_rom_inst (.q(O3_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [13-1:0] O3_I3_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O3_I3_R0_C111_rom_inst (.q(O3_I3_R0_C1_SM1 ),.address(input_fmap_3[15:8]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R0_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O3_I3_R0_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O3_I3_R0_C111_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O3_I3_R0_C111_rom_inst (.q(O3_I3_R0_C1_SM1 ),.address(input_fmap_3[15:8]),.clock  (clk));
logic [12-1:0] O3_I3_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_dw_O3_I3_R0_C24_rom_inst (.q(O3_I3_R0_C2_SM1 ),.address(input_fmap_3[23:16]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R0_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O3_I3_R0_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O3_I3_R0_C24_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_dw_O3_I3_R0_C24_rom_inst (.q(O3_I3_R0_C2_SM1 ),.address(input_fmap_3[23:16]),.clock  (clk));
logic [13-1:0] O3_I3_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O3_I3_R1_C08_rom_inst (.q(O3_I3_R1_C0_SM1 ),.address(input_fmap_3[31:24]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R1_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O3_I3_R1_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O3_I3_R1_C08_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O3_I3_R1_C08_rom_inst (.q(O3_I3_R1_C0_SM1 ),.address(input_fmap_3[31:24]),.clock  (clk));
logic [14-1:0] O3_I3_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv4_dw_O3_I3_R1_C118_rom_inst (.q(O3_I3_R1_C1_SM1 ),.address(input_fmap_3[39:32]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R1_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O3_I3_R1_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O3_I3_R1_C118_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv4_dw_O3_I3_R1_C118_rom_inst (.q(O3_I3_R1_C1_SM1 ),.address(input_fmap_3[39:32]),.clock  (clk));
logic [13-1:0] O3_I3_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O3_I3_R1_C212_rom_inst (.q(O3_I3_R1_C2_SM1 ),.address(input_fmap_3[47:40]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R1_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O3_I3_R1_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O3_I3_R1_C212_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O3_I3_R1_C212_rom_inst (.q(O3_I3_R1_C2_SM1 ),.address(input_fmap_3[47:40]),.clock  (clk));
logic [11-1:0] O3_I3_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_dw_O3_I3_R2_C02_rom_inst (.q(O3_I3_R2_C0_SM1 ),.address(input_fmap_3[55:48]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R2_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O3_I3_R2_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O3_I3_R2_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_dw_O3_I3_R2_C02_rom_inst (.q(O3_I3_R2_C0_SM1 ),.address(input_fmap_3[55:48]),.clock  (clk));
logic [13-1:0] O3_I3_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O3_I3_R2_C19_rom_inst (.q(O3_I3_R2_C1_SM1 ),.address(input_fmap_3[63:56]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R2_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O3_I3_R2_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O3_I3_R2_C19_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O3_I3_R2_C19_rom_inst (.q(O3_I3_R2_C1_SM1 ),.address(input_fmap_3[63:56]),.clock  (clk));
logic [13-1:0] O3_I3_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O3_I3_R2_C212_rom_inst (.q(O3_I3_R2_C2_SM1 ),.address(input_fmap_3[71:64]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R2_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O3_I3_R2_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O3_I3_R2_C212_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O3_I3_R2_C212_rom_inst (.q(O3_I3_R2_C2_SM1 ),.address(input_fmap_3[71:64]),.clock  (clk));
logic [13-1:0] O4_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O4_I4_R0_C09_rom_inst (.q(O4_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O4_I4_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O4_I4_R0_C09_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O4_I4_R0_C09_rom_inst (.q(O4_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [13-1:0] O4_I4_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O4_I4_R0_C19_rom_inst (.q(O4_I4_R0_C1_SM1 ),.address(input_fmap_4[15:8]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R0_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O4_I4_R0_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O4_I4_R0_C19_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O4_I4_R0_C19_rom_inst (.q(O4_I4_R0_C1_SM1 ),.address(input_fmap_4[15:8]),.clock  (clk));
logic [11-1:0] O4_I4_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_dw_O4_I4_R0_C23_rom_inst (.q(O4_I4_R0_C2_SM1 ),.address(input_fmap_4[23:16]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R0_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O4_I4_R0_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O4_I4_R0_C23_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_dw_O4_I4_R0_C23_rom_inst (.q(O4_I4_R0_C2_SM1 ),.address(input_fmap_4[23:16]),.clock  (clk));
logic [13-1:0] O4_I4_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O4_I4_R1_C015_rom_inst (.q(O4_I4_R1_C0_SM1 ),.address(input_fmap_4[31:24]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R1_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O4_I4_R1_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O4_I4_R1_C015_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O4_I4_R1_C015_rom_inst (.q(O4_I4_R1_C0_SM1 ),.address(input_fmap_4[31:24]),.clock  (clk));
logic [14-1:0] O4_I4_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv4_dw_O4_I4_R1_C118_rom_inst (.q(O4_I4_R1_C1_SM1 ),.address(input_fmap_4[39:32]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R1_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O4_I4_R1_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O4_I4_R1_C118_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv4_dw_O4_I4_R1_C118_rom_inst (.q(O4_I4_R1_C1_SM1 ),.address(input_fmap_4[39:32]),.clock  (clk));
logic [12-1:0] O4_I4_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_dw_O4_I4_R1_C27_rom_inst (.q(O4_I4_R1_C2_SM1 ),.address(input_fmap_4[47:40]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R1_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O4_I4_R1_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O4_I4_R1_C27_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_dw_O4_I4_R1_C27_rom_inst (.q(O4_I4_R1_C2_SM1 ),.address(input_fmap_4[47:40]),.clock  (clk));
logic [12-1:0] O4_I4_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_dw_O4_I4_R2_C07_rom_inst (.q(O4_I4_R2_C0_SM1 ),.address(input_fmap_4[55:48]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R2_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O4_I4_R2_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O4_I4_R2_C07_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_dw_O4_I4_R2_C07_rom_inst (.q(O4_I4_R2_C0_SM1 ),.address(input_fmap_4[55:48]),.clock  (clk));
logic [13-1:0] O4_I4_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O4_I4_R2_C110_rom_inst (.q(O4_I4_R2_C1_SM1 ),.address(input_fmap_4[63:56]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R2_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O4_I4_R2_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O4_I4_R2_C110_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O4_I4_R2_C110_rom_inst (.q(O4_I4_R2_C1_SM1 ),.address(input_fmap_4[63:56]),.clock  (clk));
logic [11-1:0] O4_I4_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_dw_O4_I4_R2_C23_rom_inst (.q(O4_I4_R2_C2_SM1 ),.address(input_fmap_4[71:64]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R2_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O4_I4_R2_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O4_I4_R2_C23_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_dw_O4_I4_R2_C23_rom_inst (.q(O4_I4_R2_C2_SM1 ),.address(input_fmap_4[71:64]),.clock  (clk));
logic [13-1:0] O5_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O5_I5_R0_C012_rom_inst (.q(O5_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O5_I5_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O5_I5_R0_C012_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O5_I5_R0_C012_rom_inst (.q(O5_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [13-1:0] O5_I5_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O5_I5_R0_C113_rom_inst (.q(O5_I5_R0_C1_SM1 ),.address(input_fmap_5[15:8]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R0_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O5_I5_R0_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O5_I5_R0_C113_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O5_I5_R0_C113_rom_inst (.q(O5_I5_R0_C1_SM1 ),.address(input_fmap_5[15:8]),.clock  (clk));
logic [10-1:0] O5_I5_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_dw_O5_I5_R0_C21_rom_inst (.q(O5_I5_R0_C2_SM1 ),.address(input_fmap_5[23:16]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R0_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I5_R0_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O5_I5_R0_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_dw_O5_I5_R0_C21_rom_inst (.q(O5_I5_R0_C2_SM1 ),.address(input_fmap_5[23:16]),.clock  (clk));
logic [13-1:0] O5_I5_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O5_I5_R1_C014_rom_inst (.q(O5_I5_R1_C0_SM1 ),.address(input_fmap_5[31:24]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R1_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O5_I5_R1_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O5_I5_R1_C014_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O5_I5_R1_C014_rom_inst (.q(O5_I5_R1_C0_SM1 ),.address(input_fmap_5[31:24]),.clock  (clk));
logic [14-1:0] O5_I5_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv4_dw_O5_I5_R1_C120_rom_inst (.q(O5_I5_R1_C1_SM1 ),.address(input_fmap_5[39:32]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R1_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O5_I5_R1_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O5_I5_R1_C120_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv4_dw_O5_I5_R1_C120_rom_inst (.q(O5_I5_R1_C1_SM1 ),.address(input_fmap_5[39:32]),.clock  (clk));
logic [12-1:0] O5_I5_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_dw_O5_I5_R1_C25_rom_inst (.q(O5_I5_R1_C2_SM1 ),.address(input_fmap_5[47:40]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R1_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O5_I5_R1_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O5_I5_R1_C25_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_dw_O5_I5_R1_C25_rom_inst (.q(O5_I5_R1_C2_SM1 ),.address(input_fmap_5[47:40]),.clock  (clk));
logic [12-1:0] O5_I5_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_dw_O5_I5_R2_C04_rom_inst (.q(O5_I5_R2_C0_SM1 ),.address(input_fmap_5[55:48]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R2_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O5_I5_R2_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O5_I5_R2_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_dw_O5_I5_R2_C04_rom_inst (.q(O5_I5_R2_C0_SM1 ),.address(input_fmap_5[55:48]),.clock  (clk));
logic [13-1:0] O5_I5_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O5_I5_R2_C110_rom_inst (.q(O5_I5_R2_C1_SM1 ),.address(input_fmap_5[63:56]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R2_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O5_I5_R2_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O5_I5_R2_C110_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O5_I5_R2_C110_rom_inst (.q(O5_I5_R2_C1_SM1 ),.address(input_fmap_5[63:56]),.clock  (clk));
logic [11-1:0] O5_I5_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_dw_O5_I5_R2_C23_rom_inst (.q(O5_I5_R2_C2_SM1 ),.address(input_fmap_5[71:64]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R2_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O5_I5_R2_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O5_I5_R2_C23_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_dw_O5_I5_R2_C23_rom_inst (.q(O5_I5_R2_C2_SM1 ),.address(input_fmap_5[71:64]),.clock  (clk));
logic [12-1:0] O6_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_dw_O6_I6_R0_C06_rom_inst (.q(O6_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O6_I6_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O6_I6_R0_C06_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_dw_O6_I6_R0_C06_rom_inst (.q(O6_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [13-1:0] O6_I6_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O6_I6_R0_C112_rom_inst (.q(O6_I6_R0_C1_SM1 ),.address(input_fmap_6[15:8]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R0_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O6_I6_R0_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O6_I6_R0_C112_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O6_I6_R0_C112_rom_inst (.q(O6_I6_R0_C1_SM1 ),.address(input_fmap_6[15:8]),.clock  (clk));
logic [13-1:0] O6_I6_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O6_I6_R0_C210_rom_inst (.q(O6_I6_R0_C2_SM1 ),.address(input_fmap_6[23:16]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R0_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O6_I6_R0_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O6_I6_R0_C210_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O6_I6_R0_C210_rom_inst (.q(O6_I6_R0_C2_SM1 ),.address(input_fmap_6[23:16]),.clock  (clk));
logic [13-1:0] O6_I6_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O6_I6_R1_C011_rom_inst (.q(O6_I6_R1_C0_SM1 ),.address(input_fmap_6[31:24]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R1_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O6_I6_R1_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O6_I6_R1_C011_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O6_I6_R1_C011_rom_inst (.q(O6_I6_R1_C0_SM1 ),.address(input_fmap_6[31:24]),.clock  (clk));
logic [14-1:0] O6_I6_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv4_dw_O6_I6_R1_C123_rom_inst (.q(O6_I6_R1_C1_SM1 ),.address(input_fmap_6[39:32]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R1_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O6_I6_R1_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O6_I6_R1_C123_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv4_dw_O6_I6_R1_C123_rom_inst (.q(O6_I6_R1_C1_SM1 ),.address(input_fmap_6[39:32]),.clock  (clk));
logic [13-1:0] O6_I6_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O6_I6_R1_C211_rom_inst (.q(O6_I6_R1_C2_SM1 ),.address(input_fmap_6[47:40]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R1_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O6_I6_R1_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O6_I6_R1_C211_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O6_I6_R1_C211_rom_inst (.q(O6_I6_R1_C2_SM1 ),.address(input_fmap_6[47:40]),.clock  (clk));
logic [12-1:0] O6_I6_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_dw_O6_I6_R2_C06_rom_inst (.q(O6_I6_R2_C0_SM1 ),.address(input_fmap_6[55:48]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R2_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O6_I6_R2_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O6_I6_R2_C06_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_dw_O6_I6_R2_C06_rom_inst (.q(O6_I6_R2_C0_SM1 ),.address(input_fmap_6[55:48]),.clock  (clk));
logic [13-1:0] O6_I6_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O6_I6_R2_C19_rom_inst (.q(O6_I6_R2_C1_SM1 ),.address(input_fmap_6[63:56]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R2_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O6_I6_R2_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O6_I6_R2_C19_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O6_I6_R2_C19_rom_inst (.q(O6_I6_R2_C1_SM1 ),.address(input_fmap_6[63:56]),.clock  (clk));
logic [11-1:0] O6_I6_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_dw_O6_I6_R2_C23_rom_inst (.q(O6_I6_R2_C2_SM1 ),.address(input_fmap_6[71:64]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R2_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O6_I6_R2_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O6_I6_R2_C23_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_dw_O6_I6_R2_C23_rom_inst (.q(O6_I6_R2_C2_SM1 ),.address(input_fmap_6[71:64]),.clock  (clk));
logic [12-1:0] O7_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_dw_O7_I7_R0_C07_rom_inst (.q(O7_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O7_I7_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O7_I7_R0_C07_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_dw_O7_I7_R0_C07_rom_inst (.q(O7_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [13-1:0] O7_I7_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O7_I7_R0_C111_rom_inst (.q(O7_I7_R0_C1_SM1 ),.address(input_fmap_7[15:8]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R0_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O7_I7_R0_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O7_I7_R0_C111_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O7_I7_R0_C111_rom_inst (.q(O7_I7_R0_C1_SM1 ),.address(input_fmap_7[15:8]),.clock  (clk));
logic [12-1:0] O7_I7_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_dw_O7_I7_R0_C27_rom_inst (.q(O7_I7_R0_C2_SM1 ),.address(input_fmap_7[23:16]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R0_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O7_I7_R0_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O7_I7_R0_C27_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_dw_O7_I7_R0_C27_rom_inst (.q(O7_I7_R0_C2_SM1 ),.address(input_fmap_7[23:16]),.clock  (clk));
logic [13-1:0] O7_I7_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O7_I7_R1_C08_rom_inst (.q(O7_I7_R1_C0_SM1 ),.address(input_fmap_7[31:24]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R1_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O7_I7_R1_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O7_I7_R1_C08_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O7_I7_R1_C08_rom_inst (.q(O7_I7_R1_C0_SM1 ),.address(input_fmap_7[31:24]),.clock  (clk));
logic [14-1:0] O7_I7_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv4_dw_O7_I7_R1_C119_rom_inst (.q(O7_I7_R1_C1_SM1 ),.address(input_fmap_7[39:32]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R1_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O7_I7_R1_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O7_I7_R1_C119_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv4_dw_O7_I7_R1_C119_rom_inst (.q(O7_I7_R1_C1_SM1 ),.address(input_fmap_7[39:32]),.clock  (clk));
logic [13-1:0] O7_I7_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O7_I7_R1_C214_rom_inst (.q(O7_I7_R1_C2_SM1 ),.address(input_fmap_7[47:40]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R1_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O7_I7_R1_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O7_I7_R1_C214_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O7_I7_R1_C214_rom_inst (.q(O7_I7_R1_C2_SM1 ),.address(input_fmap_7[47:40]),.clock  (clk));
logic [12-1:0] O7_I7_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_dw_O7_I7_R2_C04_rom_inst (.q(O7_I7_R2_C0_SM1 ),.address(input_fmap_7[55:48]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R2_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O7_I7_R2_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O7_I7_R2_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_dw_O7_I7_R2_C04_rom_inst (.q(O7_I7_R2_C0_SM1 ),.address(input_fmap_7[55:48]),.clock  (clk));
logic [13-1:0] O7_I7_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O7_I7_R2_C19_rom_inst (.q(O7_I7_R2_C1_SM1 ),.address(input_fmap_7[63:56]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R2_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O7_I7_R2_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O7_I7_R2_C19_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O7_I7_R2_C19_rom_inst (.q(O7_I7_R2_C1_SM1 ),.address(input_fmap_7[63:56]),.clock  (clk));
logic [12-1:0] O7_I7_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_dw_O7_I7_R2_C25_rom_inst (.q(O7_I7_R2_C2_SM1 ),.address(input_fmap_7[71:64]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R2_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O7_I7_R2_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O7_I7_R2_C25_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_dw_O7_I7_R2_C25_rom_inst (.q(O7_I7_R2_C2_SM1 ),.address(input_fmap_7[71:64]),.clock  (clk));
logic [13-1:0] O8_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O8_I8_R0_C08_rom_inst (.q(O8_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O8_I8_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O8_I8_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O8_I8_R0_C08_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O8_I8_R0_C08_rom_inst (.q(O8_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [13-1:0] O8_I8_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O8_I8_R0_C110_rom_inst (.q(O8_I8_R0_C1_SM1 ),.address(input_fmap_8[15:8]),.clk(clk),.d(0),.we(0));
//assign O8_I8_R0_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O8_I8_R0_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O8_I8_R0_C110_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O8_I8_R0_C110_rom_inst (.q(O8_I8_R0_C1_SM1 ),.address(input_fmap_8[15:8]),.clock  (clk));
logic [13-1:0] O8_I8_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O8_I8_R1_C015_rom_inst (.q(O8_I8_R1_C0_SM1 ),.address(input_fmap_8[31:24]),.clk(clk),.d(0),.we(0));
//assign O8_I8_R1_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O8_I8_R1_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O8_I8_R1_C015_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O8_I8_R1_C015_rom_inst (.q(O8_I8_R1_C0_SM1 ),.address(input_fmap_8[31:24]),.clock  (clk));
logic [13-1:0] O8_I8_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O8_I8_R1_C111_rom_inst (.q(O8_I8_R1_C1_SM1 ),.address(input_fmap_8[39:32]),.clk(clk),.d(0),.we(0));
//assign O8_I8_R1_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O8_I8_R1_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O8_I8_R1_C111_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O8_I8_R1_C111_rom_inst (.q(O8_I8_R1_C1_SM1 ),.address(input_fmap_8[39:32]),.clock  (clk));
logic [14-1:0] O8_I8_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv4_dw_O8_I8_R2_C022_rom_inst (.q(O8_I8_R2_C0_SM1 ),.address(input_fmap_8[55:48]),.clk(clk),.d(0),.we(0));
//assign O8_I8_R2_C0_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O8_I8_R2_C0_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O8_I8_R2_C022_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv4_dw_O8_I8_R2_C022_rom_inst (.q(O8_I8_R2_C0_SM1 ),.address(input_fmap_8[55:48]),.clock  (clk));
logic [14-1:0] O8_I8_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv4_dw_O8_I8_R2_C121_rom_inst (.q(O8_I8_R2_C1_SM1 ),.address(input_fmap_8[63:56]),.clk(clk),.d(0),.we(0));
//assign O8_I8_R2_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O8_I8_R2_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O8_I8_R2_C121_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv4_dw_O8_I8_R2_C121_rom_inst (.q(O8_I8_R2_C1_SM1 ),.address(input_fmap_8[63:56]),.clock  (clk));
logic [13-1:0] O9_I9_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O9_I9_R0_C110_rom_inst (.q(O9_I9_R0_C1_SM1 ),.address(input_fmap_9[15:8]),.clk(clk),.d(0),.we(0));
//assign O9_I9_R0_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O9_I9_R0_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O9_I9_R0_C110_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O9_I9_R0_C110_rom_inst (.q(O9_I9_R0_C1_SM1 ),.address(input_fmap_9[15:8]),.clock  (clk));
logic [13-1:0] O9_I9_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O9_I9_R0_C28_rom_inst (.q(O9_I9_R0_C2_SM1 ),.address(input_fmap_9[23:16]),.clk(clk),.d(0),.we(0));
//assign O9_I9_R0_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O9_I9_R0_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O9_I9_R0_C28_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O9_I9_R0_C28_rom_inst (.q(O9_I9_R0_C2_SM1 ),.address(input_fmap_9[23:16]),.clock  (clk));
logic [11-1:0] O9_I9_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_dw_O9_I9_R1_C02_rom_inst (.q(O9_I9_R1_C0_SM1 ),.address(input_fmap_9[31:24]),.clk(clk),.d(0),.we(0));
//assign O9_I9_R1_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O9_I9_R1_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O9_I9_R1_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_dw_O9_I9_R1_C02_rom_inst (.q(O9_I9_R1_C0_SM1 ),.address(input_fmap_9[31:24]),.clock  (clk));
logic [14-1:0] O9_I9_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv4_dw_O9_I9_R1_C118_rom_inst (.q(O9_I9_R1_C1_SM1 ),.address(input_fmap_9[39:32]),.clk(clk),.d(0),.we(0));
//assign O9_I9_R1_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O9_I9_R1_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O9_I9_R1_C118_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv4_dw_O9_I9_R1_C118_rom_inst (.q(O9_I9_R1_C1_SM1 ),.address(input_fmap_9[39:32]),.clock  (clk));
logic [14-1:0] O9_I9_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv4_dw_O9_I9_R1_C219_rom_inst (.q(O9_I9_R1_C2_SM1 ),.address(input_fmap_9[47:40]),.clk(clk),.d(0),.we(0));
//assign O9_I9_R1_C2_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O9_I9_R1_C2_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O9_I9_R1_C219_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv4_dw_O9_I9_R1_C219_rom_inst (.q(O9_I9_R1_C2_SM1 ),.address(input_fmap_9[47:40]),.clock  (clk));
logic [10-1:0] O9_I9_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_dw_O9_I9_R2_C01_rom_inst (.q(O9_I9_R2_C0_SM1 ),.address(input_fmap_9[55:48]),.clk(clk),.d(0),.we(0));
//assign O9_I9_R2_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O9_I9_R2_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O9_I9_R2_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_dw_O9_I9_R2_C01_rom_inst (.q(O9_I9_R2_C0_SM1 ),.address(input_fmap_9[55:48]),.clock  (clk));
logic [13-1:0] O9_I9_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O9_I9_R2_C110_rom_inst (.q(O9_I9_R2_C1_SM1 ),.address(input_fmap_9[63:56]),.clk(clk),.d(0),.we(0));
//assign O9_I9_R2_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O9_I9_R2_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O9_I9_R2_C110_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O9_I9_R2_C110_rom_inst (.q(O9_I9_R2_C1_SM1 ),.address(input_fmap_9[63:56]),.clock  (clk));
logic [13-1:0] O9_I9_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O9_I9_R2_C212_rom_inst (.q(O9_I9_R2_C2_SM1 ),.address(input_fmap_9[71:64]),.clk(clk),.d(0),.we(0));
//assign O9_I9_R2_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O9_I9_R2_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O9_I9_R2_C212_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O9_I9_R2_C212_rom_inst (.q(O9_I9_R2_C2_SM1 ),.address(input_fmap_9[71:64]),.clock  (clk));
logic [12-1:0] O10_I10_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_dw_O10_I10_R0_C04_rom_inst (.q(O10_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clk(clk),.d(0),.we(0));
//assign O10_I10_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O10_I10_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O10_I10_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_dw_O10_I10_R0_C04_rom_inst (.q(O10_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clock  (clk));
logic [11-1:0] O10_I10_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_dw_O10_I10_R0_C13_rom_inst (.q(O10_I10_R0_C1_SM1 ),.address(input_fmap_10[15:8]),.clk(clk),.d(0),.we(0));
//assign O10_I10_R0_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O10_I10_R0_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O10_I10_R0_C13_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_dw_O10_I10_R0_C13_rom_inst (.q(O10_I10_R0_C1_SM1 ),.address(input_fmap_10[15:8]),.clock  (clk));
logic [12-1:0] O10_I10_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_dw_O10_I10_R0_C24_rom_inst (.q(O10_I10_R0_C2_SM1 ),.address(input_fmap_10[23:16]),.clk(clk),.d(0),.we(0));
//assign O10_I10_R0_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O10_I10_R0_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O10_I10_R0_C24_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_dw_O10_I10_R0_C24_rom_inst (.q(O10_I10_R0_C2_SM1 ),.address(input_fmap_10[23:16]),.clock  (clk));
logic [12-1:0] O10_I10_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_dw_O10_I10_R1_C05_rom_inst (.q(O10_I10_R1_C0_SM1 ),.address(input_fmap_10[31:24]),.clk(clk),.d(0),.we(0));
//assign O10_I10_R1_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O10_I10_R1_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O10_I10_R1_C05_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_dw_O10_I10_R1_C05_rom_inst (.q(O10_I10_R1_C0_SM1 ),.address(input_fmap_10[31:24]),.clock  (clk));
logic [13-1:0] O10_I10_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O10_I10_R1_C111_rom_inst (.q(O10_I10_R1_C1_SM1 ),.address(input_fmap_10[39:32]),.clk(clk),.d(0),.we(0));
//assign O10_I10_R1_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O10_I10_R1_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O10_I10_R1_C111_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O10_I10_R1_C111_rom_inst (.q(O10_I10_R1_C1_SM1 ),.address(input_fmap_10[39:32]),.clock  (clk));
logic [13-1:0] O10_I10_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O10_I10_R1_C215_rom_inst (.q(O10_I10_R1_C2_SM1 ),.address(input_fmap_10[47:40]),.clk(clk),.d(0),.we(0));
//assign O10_I10_R1_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O10_I10_R1_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O10_I10_R1_C215_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O10_I10_R1_C215_rom_inst (.q(O10_I10_R1_C2_SM1 ),.address(input_fmap_10[47:40]),.clock  (clk));
logic [11-1:0] O10_I10_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_dw_O10_I10_R2_C03_rom_inst (.q(O10_I10_R2_C0_SM1 ),.address(input_fmap_10[55:48]),.clk(clk),.d(0),.we(0));
//assign O10_I10_R2_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O10_I10_R2_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O10_I10_R2_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_dw_O10_I10_R2_C03_rom_inst (.q(O10_I10_R2_C0_SM1 ),.address(input_fmap_10[55:48]),.clock  (clk));
logic [12-1:0] O10_I10_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_dw_O10_I10_R2_C17_rom_inst (.q(O10_I10_R2_C1_SM1 ),.address(input_fmap_10[63:56]),.clk(clk),.d(0),.we(0));
//assign O10_I10_R2_C1_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O10_I10_R2_C1_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O10_I10_R2_C17_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_dw_O10_I10_R2_C17_rom_inst (.q(O10_I10_R2_C1_SM1 ),.address(input_fmap_10[63:56]),.clock  (clk));
logic [13-1:0] O10_I10_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O10_I10_R2_C210_rom_inst (.q(O10_I10_R2_C2_SM1 ),.address(input_fmap_10[71:64]),.clk(clk),.d(0),.we(0));
//assign O10_I10_R2_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O10_I10_R2_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O10_I10_R2_C210_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O10_I10_R2_C210_rom_inst (.q(O10_I10_R2_C2_SM1 ),.address(input_fmap_10[71:64]),.clock  (clk));
logic [13-1:0] O11_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O11_I11_R0_C011_rom_inst (.q(O11_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I11_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O11_I11_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O11_I11_R0_C011_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O11_I11_R0_C011_rom_inst (.q(O11_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [13-1:0] O11_I11_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O11_I11_R0_C115_rom_inst (.q(O11_I11_R0_C1_SM1 ),.address(input_fmap_11[15:8]),.clk(clk),.d(0),.we(0));
//assign O11_I11_R0_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O11_I11_R0_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O11_I11_R0_C115_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O11_I11_R0_C115_rom_inst (.q(O11_I11_R0_C1_SM1 ),.address(input_fmap_11[15:8]),.clock  (clk));
logic [12-1:0] O11_I11_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_dw_O11_I11_R0_C26_rom_inst (.q(O11_I11_R0_C2_SM1 ),.address(input_fmap_11[23:16]),.clk(clk),.d(0),.we(0));
//assign O11_I11_R0_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O11_I11_R0_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O11_I11_R0_C26_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_dw_O11_I11_R0_C26_rom_inst (.q(O11_I11_R0_C2_SM1 ),.address(input_fmap_11[23:16]),.clock  (clk));
logic [13-1:0] O11_I11_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O11_I11_R1_C013_rom_inst (.q(O11_I11_R1_C0_SM1 ),.address(input_fmap_11[31:24]),.clk(clk),.d(0),.we(0));
//assign O11_I11_R1_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O11_I11_R1_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O11_I11_R1_C013_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O11_I11_R1_C013_rom_inst (.q(O11_I11_R1_C0_SM1 ),.address(input_fmap_11[31:24]),.clock  (clk));
logic [14-1:0] O11_I11_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv4_dw_O11_I11_R1_C124_rom_inst (.q(O11_I11_R1_C1_SM1 ),.address(input_fmap_11[39:32]),.clk(clk),.d(0),.we(0));
//assign O11_I11_R1_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O11_I11_R1_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O11_I11_R1_C124_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv4_dw_O11_I11_R1_C124_rom_inst (.q(O11_I11_R1_C1_SM1 ),.address(input_fmap_11[39:32]),.clock  (clk));
logic [13-1:0] O11_I11_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O11_I11_R1_C210_rom_inst (.q(O11_I11_R1_C2_SM1 ),.address(input_fmap_11[47:40]),.clk(clk),.d(0),.we(0));
//assign O11_I11_R1_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O11_I11_R1_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O11_I11_R1_C210_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O11_I11_R1_C210_rom_inst (.q(O11_I11_R1_C2_SM1 ),.address(input_fmap_11[47:40]),.clock  (clk));
logic [12-1:0] O11_I11_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_dw_O11_I11_R2_C05_rom_inst (.q(O11_I11_R2_C0_SM1 ),.address(input_fmap_11[55:48]),.clk(clk),.d(0),.we(0));
//assign O11_I11_R2_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O11_I11_R2_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O11_I11_R2_C05_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_dw_O11_I11_R2_C05_rom_inst (.q(O11_I11_R2_C0_SM1 ),.address(input_fmap_11[55:48]),.clock  (clk));
logic [13-1:0] O11_I11_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O11_I11_R2_C18_rom_inst (.q(O11_I11_R2_C1_SM1 ),.address(input_fmap_11[63:56]),.clk(clk),.d(0),.we(0));
//assign O11_I11_R2_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O11_I11_R2_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O11_I11_R2_C18_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O11_I11_R2_C18_rom_inst (.q(O11_I11_R2_C1_SM1 ),.address(input_fmap_11[63:56]),.clock  (clk));
logic [12-1:0] O11_I11_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_dw_O11_I11_R2_C24_rom_inst (.q(O11_I11_R2_C2_SM1 ),.address(input_fmap_11[71:64]),.clk(clk),.d(0),.we(0));
//assign O11_I11_R2_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O11_I11_R2_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O11_I11_R2_C24_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_dw_O11_I11_R2_C24_rom_inst (.q(O11_I11_R2_C2_SM1 ),.address(input_fmap_11[71:64]),.clock  (clk));
logic [11-1:0] O12_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_dw_O12_I12_R0_C03_rom_inst (.q(O12_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I12_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O12_I12_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O12_I12_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_dw_O12_I12_R0_C03_rom_inst (.q(O12_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [12-1:0] O12_I12_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_dw_O12_I12_R0_C17_rom_inst (.q(O12_I12_R0_C1_SM1 ),.address(input_fmap_12[15:8]),.clk(clk),.d(0),.we(0));
//assign O12_I12_R0_C1_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O12_I12_R0_C1_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O12_I12_R0_C17_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_dw_O12_I12_R0_C17_rom_inst (.q(O12_I12_R0_C1_SM1 ),.address(input_fmap_12[15:8]),.clock  (clk));
logic [12-1:0] O12_I12_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_dw_O12_I12_R0_C25_rom_inst (.q(O12_I12_R0_C2_SM1 ),.address(input_fmap_12[23:16]),.clk(clk),.d(0),.we(0));
//assign O12_I12_R0_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O12_I12_R0_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O12_I12_R0_C25_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_dw_O12_I12_R0_C25_rom_inst (.q(O12_I12_R0_C2_SM1 ),.address(input_fmap_12[23:16]),.clock  (clk));
logic [12-1:0] O12_I12_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_dw_O12_I12_R1_C05_rom_inst (.q(O12_I12_R1_C0_SM1 ),.address(input_fmap_12[31:24]),.clk(clk),.d(0),.we(0));
//assign O12_I12_R1_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O12_I12_R1_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O12_I12_R1_C05_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_dw_O12_I12_R1_C05_rom_inst (.q(O12_I12_R1_C0_SM1 ),.address(input_fmap_12[31:24]),.clock  (clk));
logic [14-1:0] O12_I12_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv4_dw_O12_I12_R1_C119_rom_inst (.q(O12_I12_R1_C1_SM1 ),.address(input_fmap_12[39:32]),.clk(clk),.d(0),.we(0));
//assign O12_I12_R1_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O12_I12_R1_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O12_I12_R1_C119_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv4_dw_O12_I12_R1_C119_rom_inst (.q(O12_I12_R1_C1_SM1 ),.address(input_fmap_12[39:32]),.clock  (clk));
logic [13-1:0] O12_I12_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O12_I12_R1_C212_rom_inst (.q(O12_I12_R1_C2_SM1 ),.address(input_fmap_12[47:40]),.clk(clk),.d(0),.we(0));
//assign O12_I12_R1_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O12_I12_R1_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O12_I12_R1_C212_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O12_I12_R1_C212_rom_inst (.q(O12_I12_R1_C2_SM1 ),.address(input_fmap_12[47:40]),.clock  (clk));
logic [13-1:0] O12_I12_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O12_I12_R2_C111_rom_inst (.q(O12_I12_R2_C1_SM1 ),.address(input_fmap_12[63:56]),.clk(clk),.d(0),.we(0));
//assign O12_I12_R2_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O12_I12_R2_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O12_I12_R2_C111_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O12_I12_R2_C111_rom_inst (.q(O12_I12_R2_C1_SM1 ),.address(input_fmap_12[63:56]),.clock  (clk));
logic [13-1:0] O12_I12_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O12_I12_R2_C28_rom_inst (.q(O12_I12_R2_C2_SM1 ),.address(input_fmap_12[71:64]),.clk(clk),.d(0),.we(0));
//assign O12_I12_R2_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O12_I12_R2_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O12_I12_R2_C28_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O12_I12_R2_C28_rom_inst (.q(O12_I12_R2_C2_SM1 ),.address(input_fmap_12[71:64]),.clock  (clk));
logic [10-1:0] O13_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_dw_O13_I13_R0_C01_rom_inst (.q(O13_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O13_I13_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O13_I13_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O13_I13_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_dw_O13_I13_R0_C01_rom_inst (.q(O13_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [13-1:0] O13_I13_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O13_I13_R0_C112_rom_inst (.q(O13_I13_R0_C1_SM1 ),.address(input_fmap_13[15:8]),.clk(clk),.d(0),.we(0));
//assign O13_I13_R0_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O13_I13_R0_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O13_I13_R0_C112_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O13_I13_R0_C112_rom_inst (.q(O13_I13_R0_C1_SM1 ),.address(input_fmap_13[15:8]),.clock  (clk));
logic [13-1:0] O13_I13_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O13_I13_R0_C211_rom_inst (.q(O13_I13_R0_C2_SM1 ),.address(input_fmap_13[23:16]),.clk(clk),.d(0),.we(0));
//assign O13_I13_R0_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O13_I13_R0_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O13_I13_R0_C211_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O13_I13_R0_C211_rom_inst (.q(O13_I13_R0_C2_SM1 ),.address(input_fmap_13[23:16]),.clock  (clk));
logic [10-1:0] O13_I13_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_dw_O13_I13_R1_C01_rom_inst (.q(O13_I13_R1_C0_SM1 ),.address(input_fmap_13[31:24]),.clk(clk),.d(0),.we(0));
//assign O13_I13_R1_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O13_I13_R1_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O13_I13_R1_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_dw_O13_I13_R1_C01_rom_inst (.q(O13_I13_R1_C0_SM1 ),.address(input_fmap_13[31:24]),.clock  (clk));
logic [13-1:0] O13_I13_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O13_I13_R1_C113_rom_inst (.q(O13_I13_R1_C1_SM1 ),.address(input_fmap_13[39:32]),.clk(clk),.d(0),.we(0));
//assign O13_I13_R1_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O13_I13_R1_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O13_I13_R1_C113_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O13_I13_R1_C113_rom_inst (.q(O13_I13_R1_C1_SM1 ),.address(input_fmap_13[39:32]),.clock  (clk));
logic [13-1:0] O13_I13_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O13_I13_R1_C214_rom_inst (.q(O13_I13_R1_C2_SM1 ),.address(input_fmap_13[47:40]),.clk(clk),.d(0),.we(0));
//assign O13_I13_R1_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O13_I13_R1_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O13_I13_R1_C214_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O13_I13_R1_C214_rom_inst (.q(O13_I13_R1_C2_SM1 ),.address(input_fmap_13[47:40]),.clock  (clk));
logic [12-1:0] O13_I13_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_dw_O13_I13_R2_C05_rom_inst (.q(O13_I13_R2_C0_SM1 ),.address(input_fmap_13[55:48]),.clk(clk),.d(0),.we(0));
//assign O13_I13_R2_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O13_I13_R2_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O13_I13_R2_C05_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_dw_O13_I13_R2_C05_rom_inst (.q(O13_I13_R2_C0_SM1 ),.address(input_fmap_13[55:48]),.clock  (clk));
logic [12-1:0] O13_I13_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_dw_O13_I13_R2_C15_rom_inst (.q(O13_I13_R2_C1_SM1 ),.address(input_fmap_13[63:56]),.clk(clk),.d(0),.we(0));
//assign O13_I13_R2_C1_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O13_I13_R2_C1_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O13_I13_R2_C15_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_dw_O13_I13_R2_C15_rom_inst (.q(O13_I13_R2_C1_SM1 ),.address(input_fmap_13[63:56]),.clock  (clk));
logic [13-1:0] O13_I13_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O13_I13_R2_C28_rom_inst (.q(O13_I13_R2_C2_SM1 ),.address(input_fmap_13[71:64]),.clk(clk),.d(0),.we(0));
//assign O13_I13_R2_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O13_I13_R2_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O13_I13_R2_C28_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O13_I13_R2_C28_rom_inst (.q(O13_I13_R2_C2_SM1 ),.address(input_fmap_13[71:64]),.clock  (clk));
logic [13-1:0] O14_I14_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O14_I14_R0_C011_rom_inst (.q(O14_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I14_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O14_I14_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O14_I14_R0_C011_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O14_I14_R0_C011_rom_inst (.q(O14_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clock  (clk));
logic [14-1:0] O14_I14_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv4_dw_O14_I14_R0_C117_rom_inst (.q(O14_I14_R0_C1_SM1 ),.address(input_fmap_14[15:8]),.clk(clk),.d(0),.we(0));
//assign O14_I14_R0_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O14_I14_R0_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O14_I14_R0_C117_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv4_dw_O14_I14_R0_C117_rom_inst (.q(O14_I14_R0_C1_SM1 ),.address(input_fmap_14[15:8]),.clock  (clk));
logic [12-1:0] O14_I14_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_dw_O14_I14_R0_C25_rom_inst (.q(O14_I14_R0_C2_SM1 ),.address(input_fmap_14[23:16]),.clk(clk),.d(0),.we(0));
//assign O14_I14_R0_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O14_I14_R0_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O14_I14_R0_C25_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_dw_O14_I14_R0_C25_rom_inst (.q(O14_I14_R0_C2_SM1 ),.address(input_fmap_14[23:16]),.clock  (clk));
logic [12-1:0] O14_I14_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_dw_O14_I14_R1_C07_rom_inst (.q(O14_I14_R1_C0_SM1 ),.address(input_fmap_14[31:24]),.clk(clk),.d(0),.we(0));
//assign O14_I14_R1_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O14_I14_R1_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O14_I14_R1_C07_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_dw_O14_I14_R1_C07_rom_inst (.q(O14_I14_R1_C0_SM1 ),.address(input_fmap_14[31:24]),.clock  (clk));
logic [14-1:0] O14_I14_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv4_dw_O14_I14_R1_C121_rom_inst (.q(O14_I14_R1_C1_SM1 ),.address(input_fmap_14[39:32]),.clk(clk),.d(0),.we(0));
//assign O14_I14_R1_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O14_I14_R1_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O14_I14_R1_C121_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv4_dw_O14_I14_R1_C121_rom_inst (.q(O14_I14_R1_C1_SM1 ),.address(input_fmap_14[39:32]),.clock  (clk));
logic [13-1:0] O14_I14_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O14_I14_R1_C212_rom_inst (.q(O14_I14_R1_C2_SM1 ),.address(input_fmap_14[47:40]),.clk(clk),.d(0),.we(0));
//assign O14_I14_R1_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O14_I14_R1_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O14_I14_R1_C212_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O14_I14_R1_C212_rom_inst (.q(O14_I14_R1_C2_SM1 ),.address(input_fmap_14[47:40]),.clock  (clk));
logic [10-1:0] O14_I14_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_dw_O14_I14_R2_C01_rom_inst (.q(O14_I14_R2_C0_SM1 ),.address(input_fmap_14[55:48]),.clk(clk),.d(0),.we(0));
//assign O14_I14_R2_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O14_I14_R2_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O14_I14_R2_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_dw_O14_I14_R2_C01_rom_inst (.q(O14_I14_R2_C0_SM1 ),.address(input_fmap_14[55:48]),.clock  (clk));
logic [12-1:0] O14_I14_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_dw_O14_I14_R2_C16_rom_inst (.q(O14_I14_R2_C1_SM1 ),.address(input_fmap_14[63:56]),.clk(clk),.d(0),.we(0));
//assign O14_I14_R2_C1_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O14_I14_R2_C1_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O14_I14_R2_C16_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_dw_O14_I14_R2_C16_rom_inst (.q(O14_I14_R2_C1_SM1 ),.address(input_fmap_14[63:56]),.clock  (clk));
logic [13-1:0] O14_I14_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O14_I14_R2_C28_rom_inst (.q(O14_I14_R2_C2_SM1 ),.address(input_fmap_14[71:64]),.clk(clk),.d(0),.we(0));
//assign O14_I14_R2_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O14_I14_R2_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O14_I14_R2_C28_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O14_I14_R2_C28_rom_inst (.q(O14_I14_R2_C2_SM1 ),.address(input_fmap_14[71:64]),.clock  (clk));
logic [13-1:0] O15_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O15_I15_R0_C010_rom_inst (.q(O15_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I15_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O15_I15_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O15_I15_R0_C010_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O15_I15_R0_C010_rom_inst (.q(O15_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [13-1:0] O15_I15_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O15_I15_R0_C110_rom_inst (.q(O15_I15_R0_C1_SM1 ),.address(input_fmap_15[15:8]),.clk(clk),.d(0),.we(0));
//assign O15_I15_R0_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O15_I15_R0_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O15_I15_R0_C110_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O15_I15_R0_C110_rom_inst (.q(O15_I15_R0_C1_SM1 ),.address(input_fmap_15[15:8]),.clock  (clk));
logic [12-1:0] O15_I15_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_dw_O15_I15_R0_C24_rom_inst (.q(O15_I15_R0_C2_SM1 ),.address(input_fmap_15[23:16]),.clk(clk),.d(0),.we(0));
//assign O15_I15_R0_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O15_I15_R0_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O15_I15_R0_C24_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_dw_O15_I15_R0_C24_rom_inst (.q(O15_I15_R0_C2_SM1 ),.address(input_fmap_15[23:16]),.clock  (clk));
logic [13-1:0] O15_I15_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O15_I15_R1_C012_rom_inst (.q(O15_I15_R1_C0_SM1 ),.address(input_fmap_15[31:24]),.clk(clk),.d(0),.we(0));
//assign O15_I15_R1_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O15_I15_R1_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O15_I15_R1_C012_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O15_I15_R1_C012_rom_inst (.q(O15_I15_R1_C0_SM1 ),.address(input_fmap_15[31:24]),.clock  (clk));
logic [13-1:0] O15_I15_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O15_I15_R1_C115_rom_inst (.q(O15_I15_R1_C1_SM1 ),.address(input_fmap_15[39:32]),.clk(clk),.d(0),.we(0));
//assign O15_I15_R1_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O15_I15_R1_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O15_I15_R1_C115_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O15_I15_R1_C115_rom_inst (.q(O15_I15_R1_C1_SM1 ),.address(input_fmap_15[39:32]),.clock  (clk));
logic [13-1:0] O15_I15_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_dw_O15_I15_R1_C28_rom_inst (.q(O15_I15_R1_C2_SM1 ),.address(input_fmap_15[47:40]),.clk(clk),.d(0),.we(0));
//assign O15_I15_R1_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O15_I15_R1_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O15_I15_R1_C28_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_dw_O15_I15_R1_C28_rom_inst (.q(O15_I15_R1_C2_SM1 ),.address(input_fmap_15[47:40]),.clock  (clk));
logic [11-1:0] O15_I15_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_dw_O15_I15_R2_C03_rom_inst (.q(O15_I15_R2_C0_SM1 ),.address(input_fmap_15[55:48]),.clk(clk),.d(0),.we(0));
//assign O15_I15_R2_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O15_I15_R2_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O15_I15_R2_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_dw_O15_I15_R2_C03_rom_inst (.q(O15_I15_R2_C0_SM1 ),.address(input_fmap_15[55:48]),.clock  (clk));
logic [12-1:0] O15_I15_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_dw_O15_I15_R2_C15_rom_inst (.q(O15_I15_R2_C1_SM1 ),.address(input_fmap_15[63:56]),.clk(clk),.d(0),.we(0));
//assign O15_I15_R2_C1_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O15_I15_R2_C1_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O15_I15_R2_C15_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_dw_O15_I15_R2_C15_rom_inst (.q(O15_I15_R2_C1_SM1 ),.address(input_fmap_15[63:56]),.clock  (clk));
logic [12-1:0] O15_I15_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_dw_O15_I15_R2_C27_rom_inst (.q(O15_I15_R2_C2_SM1 ),.address(input_fmap_15[71:64]),.clk(clk),.d(0),.we(0));
//assign O15_I15_R2_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O15_I15_R2_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_dw_O15_I15_R2_C27_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_dw_O15_I15_R2_C27_rom_inst (.q(O15_I15_R2_C2_SM1 ),.address(input_fmap_15[71:64]),.clock  (clk));
logic signed [31:0] conv_mac_0;
logic signed [31:0] O0_N0_S0;		always @(posedge clk) O0_N0_S0 <=     O0_I0_R0_C0_SM1   +  O0_I0_R0_C1_SM1  ;
 logic signed [31:0] O0_N2_S0;		always @(posedge clk) O0_N2_S0 <=     O0_I0_R0_C2_SM1   +  O0_I0_R1_C0_SM1  ;
 logic signed [31:0] O0_N4_S0;		always @(posedge clk) O0_N4_S0 <=     O0_I0_R1_C1_SM1   +  O0_I0_R1_C2_SM1  ;
 logic signed [31:0] O0_N6_S0;		always @(posedge clk) O0_N6_S0 <=     O0_I0_R2_C0_SM1   +  O0_I0_R2_C1_SM1  ;
 logic signed [31:0] O0_N8_S0;		always @(posedge clk) O0_N8_S0 <=     O0_I0_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O0_N0_S1;		always @(posedge clk) O0_N0_S1 <=     O0_N0_S0  +  O0_N2_S0 ;
 logic signed [31:0] O0_N2_S1;		always @(posedge clk) O0_N2_S1 <=     O0_N4_S0  +  O0_N6_S0 ;
 logic signed [31:0] O0_N4_S1;		always @(posedge clk) O0_N4_S1 <=     O0_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O0_N0_S2;		always @(posedge clk) O0_N0_S2 <=     O0_N0_S1  +  O0_N2_S1 ;
 logic signed [31:0] O0_N2_S2;		always @(posedge clk) O0_N2_S2 <=     O0_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O0_N0_S3;		always @(posedge clk) O0_N0_S3 <=     O0_N0_S2  +  O0_N2_S2 ;
 assign conv_mac_0 = O0_N0_S3;

logic signed [31:0] conv_mac_1;
logic signed [31:0] O1_N0_S0;		always @(posedge clk) O1_N0_S0 <=     O1_I1_R0_C0_SM1   +  O1_I1_R0_C1_SM1  ;
 logic signed [31:0] O1_N2_S0;		always @(posedge clk) O1_N2_S0 <=     O1_I1_R0_C2_SM1   +  O1_I1_R1_C0_SM1  ;
 logic signed [31:0] O1_N4_S0;		always @(posedge clk) O1_N4_S0 <=     O1_I1_R1_C1_SM1   +  O1_I1_R1_C2_SM1  ;
 logic signed [31:0] O1_N6_S0;		always @(posedge clk) O1_N6_S0 <=     O1_I1_R2_C0_SM1   +  O1_I1_R2_C1_SM1  ;
 logic signed [31:0] O1_N8_S0;		always @(posedge clk) O1_N8_S0 <=     O1_I1_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O1_N0_S1;		always @(posedge clk) O1_N0_S1 <=     O1_N0_S0  +  O1_N2_S0 ;
 logic signed [31:0] O1_N2_S1;		always @(posedge clk) O1_N2_S1 <=     O1_N4_S0  +  O1_N6_S0 ;
 logic signed [31:0] O1_N4_S1;		always @(posedge clk) O1_N4_S1 <=     O1_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O1_N0_S2;		always @(posedge clk) O1_N0_S2 <=     O1_N0_S1  +  O1_N2_S1 ;
 logic signed [31:0] O1_N2_S2;		always @(posedge clk) O1_N2_S2 <=     O1_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O1_N0_S3;		always @(posedge clk) O1_N0_S3 <=     O1_N0_S2  +  O1_N2_S2 ;
 assign conv_mac_1 = O1_N0_S3;

logic signed [31:0] conv_mac_2;
logic signed [31:0] O2_N0_S0;		always @(posedge clk) O2_N0_S0 <=     O2_I2_R0_C0_SM1   +  O2_I2_R0_C1_SM1  ;
 logic signed [31:0] O2_N2_S0;		always @(posedge clk) O2_N2_S0 <=     O2_I2_R0_C2_SM1   +  O2_I2_R1_C0_SM1  ;
 logic signed [31:0] O2_N4_S0;		always @(posedge clk) O2_N4_S0 <=     O2_I2_R1_C1_SM1   +  O2_I2_R1_C2_SM1  ;
 logic signed [31:0] O2_N6_S0;		always @(posedge clk) O2_N6_S0 <=     O2_I2_R2_C0_SM1   +  O2_I2_R2_C1_SM1  ;
 logic signed [31:0] O2_N8_S0;		always @(posedge clk) O2_N8_S0 <=     O2_I2_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O2_N0_S1;		always @(posedge clk) O2_N0_S1 <=     O2_N0_S0  +  O2_N2_S0 ;
 logic signed [31:0] O2_N2_S1;		always @(posedge clk) O2_N2_S1 <=     O2_N4_S0  +  O2_N6_S0 ;
 logic signed [31:0] O2_N4_S1;		always @(posedge clk) O2_N4_S1 <=     O2_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O2_N0_S2;		always @(posedge clk) O2_N0_S2 <=     O2_N0_S1  +  O2_N2_S1 ;
 logic signed [31:0] O2_N2_S2;		always @(posedge clk) O2_N2_S2 <=     O2_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O2_N0_S3;		always @(posedge clk) O2_N0_S3 <=     O2_N0_S2  +  O2_N2_S2 ;
 assign conv_mac_2 = O2_N0_S3;

logic signed [31:0] conv_mac_3;
logic signed [31:0] O3_N0_S0;		always @(posedge clk) O3_N0_S0 <=     O3_I3_R0_C0_SM1   +  O3_I3_R0_C1_SM1  ;
 logic signed [31:0] O3_N2_S0;		always @(posedge clk) O3_N2_S0 <=     O3_I3_R0_C2_SM1   +  O3_I3_R1_C0_SM1  ;
 logic signed [31:0] O3_N4_S0;		always @(posedge clk) O3_N4_S0 <=     O3_I3_R1_C1_SM1   +  O3_I3_R1_C2_SM1  ;
 logic signed [31:0] O3_N6_S0;		always @(posedge clk) O3_N6_S0 <=     O3_I3_R2_C0_SM1   +  O3_I3_R2_C1_SM1  ;
 logic signed [31:0] O3_N8_S0;		always @(posedge clk) O3_N8_S0 <=     O3_I3_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O3_N0_S1;		always @(posedge clk) O3_N0_S1 <=     O3_N0_S0  +  O3_N2_S0 ;
 logic signed [31:0] O3_N2_S1;		always @(posedge clk) O3_N2_S1 <=     O3_N4_S0  +  O3_N6_S0 ;
 logic signed [31:0] O3_N4_S1;		always @(posedge clk) O3_N4_S1 <=     O3_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O3_N0_S2;		always @(posedge clk) O3_N0_S2 <=     O3_N0_S1  +  O3_N2_S1 ;
 logic signed [31:0] O3_N2_S2;		always @(posedge clk) O3_N2_S2 <=     O3_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O3_N0_S3;		always @(posedge clk) O3_N0_S3 <=     O3_N0_S2  +  O3_N2_S2 ;
 assign conv_mac_3 = O3_N0_S3;

logic signed [31:0] conv_mac_4;
logic signed [31:0] O4_N0_S0;		always @(posedge clk) O4_N0_S0 <=     O4_I4_R0_C0_SM1   +  O4_I4_R0_C1_SM1  ;
 logic signed [31:0] O4_N2_S0;		always @(posedge clk) O4_N2_S0 <=     O4_I4_R0_C2_SM1   +  O4_I4_R1_C0_SM1  ;
 logic signed [31:0] O4_N4_S0;		always @(posedge clk) O4_N4_S0 <=     O4_I4_R1_C1_SM1   +  O4_I4_R1_C2_SM1  ;
 logic signed [31:0] O4_N6_S0;		always @(posedge clk) O4_N6_S0 <=     O4_I4_R2_C0_SM1   +  O4_I4_R2_C1_SM1  ;
 logic signed [31:0] O4_N8_S0;		always @(posedge clk) O4_N8_S0 <=     O4_I4_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O4_N0_S1;		always @(posedge clk) O4_N0_S1 <=     O4_N0_S0  +  O4_N2_S0 ;
 logic signed [31:0] O4_N2_S1;		always @(posedge clk) O4_N2_S1 <=     O4_N4_S0  +  O4_N6_S0 ;
 logic signed [31:0] O4_N4_S1;		always @(posedge clk) O4_N4_S1 <=     O4_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O4_N0_S2;		always @(posedge clk) O4_N0_S2 <=     O4_N0_S1  +  O4_N2_S1 ;
 logic signed [31:0] O4_N2_S2;		always @(posedge clk) O4_N2_S2 <=     O4_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O4_N0_S3;		always @(posedge clk) O4_N0_S3 <=     O4_N0_S2  +  O4_N2_S2 ;
 assign conv_mac_4 = O4_N0_S3;

logic signed [31:0] conv_mac_5;
logic signed [31:0] O5_N0_S0;		always @(posedge clk) O5_N0_S0 <=     O5_I5_R0_C0_SM1   +  O5_I5_R0_C1_SM1  ;
 logic signed [31:0] O5_N2_S0;		always @(posedge clk) O5_N2_S0 <=     O5_I5_R0_C2_SM1   +  O5_I5_R1_C0_SM1  ;
 logic signed [31:0] O5_N4_S0;		always @(posedge clk) O5_N4_S0 <=     O5_I5_R1_C1_SM1   +  O5_I5_R1_C2_SM1  ;
 logic signed [31:0] O5_N6_S0;		always @(posedge clk) O5_N6_S0 <=     O5_I5_R2_C0_SM1   +  O5_I5_R2_C1_SM1  ;
 logic signed [31:0] O5_N8_S0;		always @(posedge clk) O5_N8_S0 <=     O5_I5_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O5_N0_S1;		always @(posedge clk) O5_N0_S1 <=     O5_N0_S0  +  O5_N2_S0 ;
 logic signed [31:0] O5_N2_S1;		always @(posedge clk) O5_N2_S1 <=     O5_N4_S0  +  O5_N6_S0 ;
 logic signed [31:0] O5_N4_S1;		always @(posedge clk) O5_N4_S1 <=     O5_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O5_N0_S2;		always @(posedge clk) O5_N0_S2 <=     O5_N0_S1  +  O5_N2_S1 ;
 logic signed [31:0] O5_N2_S2;		always @(posedge clk) O5_N2_S2 <=     O5_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O5_N0_S3;		always @(posedge clk) O5_N0_S3 <=     O5_N0_S2  +  O5_N2_S2 ;
 assign conv_mac_5 = O5_N0_S3;

logic signed [31:0] conv_mac_6;
logic signed [31:0] O6_N0_S0;		always @(posedge clk) O6_N0_S0 <=     O6_I6_R0_C0_SM1   +  O6_I6_R0_C1_SM1  ;
 logic signed [31:0] O6_N2_S0;		always @(posedge clk) O6_N2_S0 <=     O6_I6_R0_C2_SM1   +  O6_I6_R1_C0_SM1  ;
 logic signed [31:0] O6_N4_S0;		always @(posedge clk) O6_N4_S0 <=     O6_I6_R1_C1_SM1   +  O6_I6_R1_C2_SM1  ;
 logic signed [31:0] O6_N6_S0;		always @(posedge clk) O6_N6_S0 <=     O6_I6_R2_C0_SM1   +  O6_I6_R2_C1_SM1  ;
 logic signed [31:0] O6_N8_S0;		always @(posedge clk) O6_N8_S0 <=     O6_I6_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O6_N0_S1;		always @(posedge clk) O6_N0_S1 <=     O6_N0_S0  +  O6_N2_S0 ;
 logic signed [31:0] O6_N2_S1;		always @(posedge clk) O6_N2_S1 <=     O6_N4_S0  +  O6_N6_S0 ;
 logic signed [31:0] O6_N4_S1;		always @(posedge clk) O6_N4_S1 <=     O6_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O6_N0_S2;		always @(posedge clk) O6_N0_S2 <=     O6_N0_S1  +  O6_N2_S1 ;
 logic signed [31:0] O6_N2_S2;		always @(posedge clk) O6_N2_S2 <=     O6_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O6_N0_S3;		always @(posedge clk) O6_N0_S3 <=     O6_N0_S2  +  O6_N2_S2 ;
 assign conv_mac_6 = O6_N0_S3;

logic signed [31:0] conv_mac_7;
logic signed [31:0] O7_N0_S0;		always @(posedge clk) O7_N0_S0 <=     O7_I7_R0_C0_SM1   +  O7_I7_R0_C1_SM1  ;
 logic signed [31:0] O7_N2_S0;		always @(posedge clk) O7_N2_S0 <=     O7_I7_R0_C2_SM1   +  O7_I7_R1_C0_SM1  ;
 logic signed [31:0] O7_N4_S0;		always @(posedge clk) O7_N4_S0 <=     O7_I7_R1_C1_SM1   +  O7_I7_R1_C2_SM1  ;
 logic signed [31:0] O7_N6_S0;		always @(posedge clk) O7_N6_S0 <=     O7_I7_R2_C0_SM1   +  O7_I7_R2_C1_SM1  ;
 logic signed [31:0] O7_N8_S0;		always @(posedge clk) O7_N8_S0 <=     O7_I7_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O7_N0_S1;		always @(posedge clk) O7_N0_S1 <=     O7_N0_S0  +  O7_N2_S0 ;
 logic signed [31:0] O7_N2_S1;		always @(posedge clk) O7_N2_S1 <=     O7_N4_S0  +  O7_N6_S0 ;
 logic signed [31:0] O7_N4_S1;		always @(posedge clk) O7_N4_S1 <=     O7_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O7_N0_S2;		always @(posedge clk) O7_N0_S2 <=     O7_N0_S1  +  O7_N2_S1 ;
 logic signed [31:0] O7_N2_S2;		always @(posedge clk) O7_N2_S2 <=     O7_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O7_N0_S3;		always @(posedge clk) O7_N0_S3 <=     O7_N0_S2  +  O7_N2_S2 ;
 assign conv_mac_7 = O7_N0_S3;

logic signed [31:0] conv_mac_8;
logic signed [31:0] O8_N0_S0;		always @(posedge clk) O8_N0_S0 <=     O8_I8_R0_C0_SM1   +  O8_I8_R0_C1_SM1  ;
 logic signed [31:0] O8_N2_S0;		always @(posedge clk) O8_N2_S0 <=     O8_I8_R1_C0_SM1   +  O8_I8_R1_C1_SM1  ;
 logic signed [31:0] O8_N4_S0;		always @(posedge clk) O8_N4_S0 <=     O8_I8_R2_C0_SM1   +  O8_I8_R2_C1_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O8_N0_S1;		always @(posedge clk) O8_N0_S1 <=     O8_N0_S0  +  O8_N2_S0 ;
 logic signed [31:0] O8_N2_S1;		always @(posedge clk) O8_N2_S1 <=     O8_N4_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O8_N0_S2;		always @(posedge clk) O8_N0_S2 <=     O8_N0_S1  +  O8_N2_S1 ;
 assign conv_mac_8 = O8_N0_S2;

logic signed [31:0] conv_mac_9;
logic signed [31:0] O9_N0_S0;		always @(posedge clk) O9_N0_S0 <=     O9_I9_R0_C1_SM1   +  O9_I9_R0_C2_SM1  ;
 logic signed [31:0] O9_N2_S0;		always @(posedge clk) O9_N2_S0 <=     O9_I9_R1_C0_SM1   +  O9_I9_R1_C1_SM1  ;
 logic signed [31:0] O9_N4_S0;		always @(posedge clk) O9_N4_S0 <=     O9_I9_R1_C2_SM1   +  O9_I9_R2_C0_SM1  ;
 logic signed [31:0] O9_N6_S0;		always @(posedge clk) O9_N6_S0 <=     O9_I9_R2_C1_SM1   +  O9_I9_R2_C2_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O9_N0_S1;		always @(posedge clk) O9_N0_S1 <=     O9_N0_S0  +  O9_N2_S0 ;
 logic signed [31:0] O9_N2_S1;		always @(posedge clk) O9_N2_S1 <=     O9_N4_S0  +  O9_N6_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O9_N0_S2;		always @(posedge clk) O9_N0_S2 <=     O9_N0_S1  +  O9_N2_S1 ;
 assign conv_mac_9 = O9_N0_S2;

logic signed [31:0] conv_mac_10;
logic signed [31:0] O10_N0_S0;		always @(posedge clk) O10_N0_S0 <=     O10_I10_R0_C0_SM1   +  O10_I10_R0_C1_SM1  ;
 logic signed [31:0] O10_N2_S0;		always @(posedge clk) O10_N2_S0 <=     O10_I10_R0_C2_SM1   +  O10_I10_R1_C0_SM1  ;
 logic signed [31:0] O10_N4_S0;		always @(posedge clk) O10_N4_S0 <=     O10_I10_R1_C1_SM1   +  O10_I10_R1_C2_SM1  ;
 logic signed [31:0] O10_N6_S0;		always @(posedge clk) O10_N6_S0 <=     O10_I10_R2_C0_SM1   +  O10_I10_R2_C1_SM1  ;
 logic signed [31:0] O10_N8_S0;		always @(posedge clk) O10_N8_S0 <=     O10_I10_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O10_N0_S1;		always @(posedge clk) O10_N0_S1 <=     O10_N0_S0  +  O10_N2_S0 ;
 logic signed [31:0] O10_N2_S1;		always @(posedge clk) O10_N2_S1 <=     O10_N4_S0  +  O10_N6_S0 ;
 logic signed [31:0] O10_N4_S1;		always @(posedge clk) O10_N4_S1 <=     O10_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O10_N0_S2;		always @(posedge clk) O10_N0_S2 <=     O10_N0_S1  +  O10_N2_S1 ;
 logic signed [31:0] O10_N2_S2;		always @(posedge clk) O10_N2_S2 <=     O10_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O10_N0_S3;		always @(posedge clk) O10_N0_S3 <=     O10_N0_S2  +  O10_N2_S2 ;
 assign conv_mac_10 = O10_N0_S3;

logic signed [31:0] conv_mac_11;
logic signed [31:0] O11_N0_S0;		always @(posedge clk) O11_N0_S0 <=     O11_I11_R0_C0_SM1   +  O11_I11_R0_C1_SM1  ;
 logic signed [31:0] O11_N2_S0;		always @(posedge clk) O11_N2_S0 <=     O11_I11_R0_C2_SM1   +  O11_I11_R1_C0_SM1  ;
 logic signed [31:0] O11_N4_S0;		always @(posedge clk) O11_N4_S0 <=     O11_I11_R1_C1_SM1   +  O11_I11_R1_C2_SM1  ;
 logic signed [31:0] O11_N6_S0;		always @(posedge clk) O11_N6_S0 <=     O11_I11_R2_C0_SM1   +  O11_I11_R2_C1_SM1  ;
 logic signed [31:0] O11_N8_S0;		always @(posedge clk) O11_N8_S0 <=     O11_I11_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O11_N0_S1;		always @(posedge clk) O11_N0_S1 <=     O11_N0_S0  +  O11_N2_S0 ;
 logic signed [31:0] O11_N2_S1;		always @(posedge clk) O11_N2_S1 <=     O11_N4_S0  +  O11_N6_S0 ;
 logic signed [31:0] O11_N4_S1;		always @(posedge clk) O11_N4_S1 <=     O11_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O11_N0_S2;		always @(posedge clk) O11_N0_S2 <=     O11_N0_S1  +  O11_N2_S1 ;
 logic signed [31:0] O11_N2_S2;		always @(posedge clk) O11_N2_S2 <=     O11_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O11_N0_S3;		always @(posedge clk) O11_N0_S3 <=     O11_N0_S2  +  O11_N2_S2 ;
 assign conv_mac_11 = O11_N0_S3;

logic signed [31:0] conv_mac_12;
logic signed [31:0] O12_N0_S0;		always @(posedge clk) O12_N0_S0 <=     O12_I12_R0_C0_SM1   +  O12_I12_R0_C1_SM1  ;
 logic signed [31:0] O12_N2_S0;		always @(posedge clk) O12_N2_S0 <=     O12_I12_R0_C2_SM1   +  O12_I12_R1_C0_SM1  ;
 logic signed [31:0] O12_N4_S0;		always @(posedge clk) O12_N4_S0 <=     O12_I12_R1_C1_SM1   +  O12_I12_R1_C2_SM1  ;
 logic signed [31:0] O12_N6_S0;		always @(posedge clk) O12_N6_S0 <=     O12_I12_R2_C1_SM1   +  O12_I12_R2_C2_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O12_N0_S1;		always @(posedge clk) O12_N0_S1 <=     O12_N0_S0  +  O12_N2_S0 ;
 logic signed [31:0] O12_N2_S1;		always @(posedge clk) O12_N2_S1 <=     O12_N4_S0  +  O12_N6_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O12_N0_S2;		always @(posedge clk) O12_N0_S2 <=     O12_N0_S1  +  O12_N2_S1 ;
 assign conv_mac_12 = O12_N0_S2;

logic signed [31:0] conv_mac_13;
logic signed [31:0] O13_N0_S0;		always @(posedge clk) O13_N0_S0 <=     O13_I13_R0_C0_SM1   +  O13_I13_R0_C1_SM1  ;
 logic signed [31:0] O13_N2_S0;		always @(posedge clk) O13_N2_S0 <=     O13_I13_R0_C2_SM1   +  O13_I13_R1_C0_SM1  ;
 logic signed [31:0] O13_N4_S0;		always @(posedge clk) O13_N4_S0 <=     O13_I13_R1_C1_SM1   +  O13_I13_R1_C2_SM1  ;
 logic signed [31:0] O13_N6_S0;		always @(posedge clk) O13_N6_S0 <=     O13_I13_R2_C0_SM1   +  O13_I13_R2_C1_SM1  ;
 logic signed [31:0] O13_N8_S0;		always @(posedge clk) O13_N8_S0 <=     O13_I13_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O13_N0_S1;		always @(posedge clk) O13_N0_S1 <=     O13_N0_S0  +  O13_N2_S0 ;
 logic signed [31:0] O13_N2_S1;		always @(posedge clk) O13_N2_S1 <=     O13_N4_S0  +  O13_N6_S0 ;
 logic signed [31:0] O13_N4_S1;		always @(posedge clk) O13_N4_S1 <=     O13_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O13_N0_S2;		always @(posedge clk) O13_N0_S2 <=     O13_N0_S1  +  O13_N2_S1 ;
 logic signed [31:0] O13_N2_S2;		always @(posedge clk) O13_N2_S2 <=     O13_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O13_N0_S3;		always @(posedge clk) O13_N0_S3 <=     O13_N0_S2  +  O13_N2_S2 ;
 assign conv_mac_13 = O13_N0_S3;

logic signed [31:0] conv_mac_14;
logic signed [31:0] O14_N0_S0;		always @(posedge clk) O14_N0_S0 <=     O14_I14_R0_C0_SM1   +  O14_I14_R0_C1_SM1  ;
 logic signed [31:0] O14_N2_S0;		always @(posedge clk) O14_N2_S0 <=     O14_I14_R0_C2_SM1   +  O14_I14_R1_C0_SM1  ;
 logic signed [31:0] O14_N4_S0;		always @(posedge clk) O14_N4_S0 <=     O14_I14_R1_C1_SM1   +  O14_I14_R1_C2_SM1  ;
 logic signed [31:0] O14_N6_S0;		always @(posedge clk) O14_N6_S0 <=     O14_I14_R2_C0_SM1   +  O14_I14_R2_C1_SM1  ;
 logic signed [31:0] O14_N8_S0;		always @(posedge clk) O14_N8_S0 <=     O14_I14_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O14_N0_S1;		always @(posedge clk) O14_N0_S1 <=     O14_N0_S0  +  O14_N2_S0 ;
 logic signed [31:0] O14_N2_S1;		always @(posedge clk) O14_N2_S1 <=     O14_N4_S0  +  O14_N6_S0 ;
 logic signed [31:0] O14_N4_S1;		always @(posedge clk) O14_N4_S1 <=     O14_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O14_N0_S2;		always @(posedge clk) O14_N0_S2 <=     O14_N0_S1  +  O14_N2_S1 ;
 logic signed [31:0] O14_N2_S2;		always @(posedge clk) O14_N2_S2 <=     O14_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O14_N0_S3;		always @(posedge clk) O14_N0_S3 <=     O14_N0_S2  +  O14_N2_S2 ;
 assign conv_mac_14 = O14_N0_S3;

logic signed [31:0] conv_mac_15;
logic signed [31:0] O15_N0_S0;		always @(posedge clk) O15_N0_S0 <=     O15_I15_R0_C0_SM1   +  O15_I15_R0_C1_SM1  ;
 logic signed [31:0] O15_N2_S0;		always @(posedge clk) O15_N2_S0 <=     O15_I15_R0_C2_SM1   +  O15_I15_R1_C0_SM1  ;
 logic signed [31:0] O15_N4_S0;		always @(posedge clk) O15_N4_S0 <=     O15_I15_R1_C1_SM1   +  O15_I15_R1_C2_SM1  ;
 logic signed [31:0] O15_N6_S0;		always @(posedge clk) O15_N6_S0 <=     O15_I15_R2_C0_SM1   +  O15_I15_R2_C1_SM1  ;
 logic signed [31:0] O15_N8_S0;		always @(posedge clk) O15_N8_S0 <=     O15_I15_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O15_N0_S1;		always @(posedge clk) O15_N0_S1 <=     O15_N0_S0  +  O15_N2_S0 ;
 logic signed [31:0] O15_N2_S1;		always @(posedge clk) O15_N2_S1 <=     O15_N4_S0  +  O15_N6_S0 ;
 logic signed [31:0] O15_N4_S1;		always @(posedge clk) O15_N4_S1 <=     O15_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O15_N0_S2;		always @(posedge clk) O15_N0_S2 <=     O15_N0_S1  +  O15_N2_S1 ;
 logic signed [31:0] O15_N2_S2;		always @(posedge clk) O15_N2_S2 <=     O15_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O15_N0_S3;		always @(posedge clk) O15_N0_S3 <=     O15_N0_S2  +  O15_N2_S2 ;
 assign conv_mac_15 = O15_N0_S3;

logic valid_D1;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D1<= 0 ;
	else valid_D1<=valid;
end
logic valid_D2;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D2<= 0 ;
	else valid_D2<=valid_D1;
end
logic valid_D3;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D3<= 0 ;
	else valid_D3<=valid_D2;
end
logic valid_D4;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D4<= 0 ;
	else valid_D4<=valid_D3;
end
logic valid_D5;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D5<= 0 ;
	else valid_D5<=valid_D4;
end
always_ff @(posedge clk) begin
	if (rstn == 0) ready <= 0 ;
	else ready <=valid_D5;
end
logic [31:0] bias_add_0;
assign bias_add_0 = conv_mac_0 - 2'd1;
logic [31:0] bias_add_1;
assign bias_add_1 = conv_mac_1 + 8'd82;
logic [31:0] bias_add_2;
assign bias_add_2 = conv_mac_2 + 5'd12;
logic [31:0] bias_add_3;
assign bias_add_3 = conv_mac_3 + 4'd7;
logic [31:0] bias_add_4;
assign bias_add_4 = conv_mac_4 + 7'd57;
logic [31:0] bias_add_5;
assign bias_add_5 = conv_mac_5 + 5'd12;
logic [31:0] bias_add_6;
assign bias_add_6 = conv_mac_6 + 7'd45;
logic [31:0] bias_add_7;
assign bias_add_7 = conv_mac_7 + 5'd13;
logic [31:0] bias_add_8;
assign bias_add_8 = conv_mac_8 + 7'd47;
logic [31:0] bias_add_9;
assign bias_add_9 = conv_mac_9 + 4'd7;
logic [31:0] bias_add_10;
assign bias_add_10 = conv_mac_10 + 5'd9;
logic [31:0] bias_add_11;
assign bias_add_11 = conv_mac_11 + 6'd19;
logic [31:0] bias_add_12;
assign bias_add_12 = conv_mac_12 + 7'd36;
logic [31:0] bias_add_13;
assign bias_add_13 = conv_mac_13 - 4'd6;
logic [31:0] bias_add_14;
assign bias_add_14 = conv_mac_14 + 8'd77;
logic [31:0] bias_add_15;
assign bias_add_15 = conv_mac_15 + 7'd46;

logic [7:0] relu_0;
assign relu_0[7:0] = (bias_add_0[31]==0) ? ((bias_add_0<3'd6) ? {{bias_add_0[31],bias_add_0[10:4]}} :'d6) : '0;
logic [7:0] relu_1;
assign relu_1[7:0] = (bias_add_1[31]==0) ? ((bias_add_1<3'd6) ? {{bias_add_1[31],bias_add_1[10:4]}} :'d6) : '0;
logic [7:0] relu_2;
assign relu_2[7:0] = (bias_add_2[31]==0) ? ((bias_add_2<3'd6) ? {{bias_add_2[31],bias_add_2[10:4]}} :'d6) : '0;
logic [7:0] relu_3;
assign relu_3[7:0] = (bias_add_3[31]==0) ? ((bias_add_3<3'd6) ? {{bias_add_3[31],bias_add_3[10:4]}} :'d6) : '0;
logic [7:0] relu_4;
assign relu_4[7:0] = (bias_add_4[31]==0) ? ((bias_add_4<3'd6) ? {{bias_add_4[31],bias_add_4[10:4]}} :'d6) : '0;
logic [7:0] relu_5;
assign relu_5[7:0] = (bias_add_5[31]==0) ? ((bias_add_5<3'd6) ? {{bias_add_5[31],bias_add_5[10:4]}} :'d6) : '0;
logic [7:0] relu_6;
assign relu_6[7:0] = (bias_add_6[31]==0) ? ((bias_add_6<3'd6) ? {{bias_add_6[31],bias_add_6[10:4]}} :'d6) : '0;
logic [7:0] relu_7;
assign relu_7[7:0] = (bias_add_7[31]==0) ? ((bias_add_7<3'd6) ? {{bias_add_7[31],bias_add_7[10:4]}} :'d6) : '0;
logic [7:0] relu_8;
assign relu_8[7:0] = (bias_add_8[31]==0) ? ((bias_add_8<3'd6) ? {{bias_add_8[31],bias_add_8[10:4]}} :'d6) : '0;
logic [7:0] relu_9;
assign relu_9[7:0] = (bias_add_9[31]==0) ? ((bias_add_9<3'd6) ? {{bias_add_9[31],bias_add_9[10:4]}} :'d6) : '0;
logic [7:0] relu_10;
assign relu_10[7:0] = (bias_add_10[31]==0) ? ((bias_add_10<3'd6) ? {{bias_add_10[31],bias_add_10[10:4]}} :'d6) : '0;
logic [7:0] relu_11;
assign relu_11[7:0] = (bias_add_11[31]==0) ? ((bias_add_11<3'd6) ? {{bias_add_11[31],bias_add_11[10:4]}} :'d6) : '0;
logic [7:0] relu_12;
assign relu_12[7:0] = (bias_add_12[31]==0) ? ((bias_add_12<3'd6) ? {{bias_add_12[31],bias_add_12[10:4]}} :'d6) : '0;
logic [7:0] relu_13;
assign relu_13[7:0] = (bias_add_13[31]==0) ? ((bias_add_13<3'd6) ? {{bias_add_13[31],bias_add_13[10:4]}} :'d6) : '0;
logic [7:0] relu_14;
assign relu_14[7:0] = (bias_add_14[31]==0) ? ((bias_add_14<3'd6) ? {{bias_add_14[31],bias_add_14[10:4]}} :'d6) : '0;
logic [7:0] relu_15;
assign relu_15[7:0] = (bias_add_15[31]==0) ? ((bias_add_15<3'd6) ? {{bias_add_15[31],bias_add_15[10:4]}} :'d6) : '0;

assign output_act = {
	relu_15,
	relu_14,
	relu_13,
	relu_12,
	relu_11,
	relu_10,
	relu_9,
	relu_8,
	relu_7,
	relu_6,
	relu_5,
	relu_4,
	relu_3,
	relu_2,
	relu_1,
	relu_0
};

endmodule
module conv5_dw (
    input logic clk,
    input logic rstn,
    input logic valid,
    input logic [32*72-1:0] input_act,
    output logic [256-1:0] output_act,
    output logic ready
);
logic we;
logic [8:0] zero_number; 
assign zero_number = 9'd0; 
logic [32*72-1:0] input_act_ff;
genvar i;
generate
for (i=0;i<32;i++)
    begin: genblk_10
        always_ff @(posedge clk) begin
            if (rstn == 0) begin
                input_act_ff[(i+1)*72-1:i*72] <= '0;
            end
            else begin
                input_act_ff[(i+1)*72-1:i*72] <= input_act[(i+1)*72-1:i*72];
            end
        end
    end
endgenerate
logic [71:0] input_fmap_0;
assign input_fmap_0 = input_act_ff[71:0];
logic [71:0] input_fmap_1;
assign input_fmap_1 = input_act_ff[143:72];
logic [71:0] input_fmap_2;
assign input_fmap_2 = input_act_ff[215:144];
logic [71:0] input_fmap_3;
assign input_fmap_3 = input_act_ff[287:216];
logic [71:0] input_fmap_4;
assign input_fmap_4 = input_act_ff[359:288];
logic [71:0] input_fmap_5;
assign input_fmap_5 = input_act_ff[431:360];
logic [71:0] input_fmap_6;
assign input_fmap_6 = input_act_ff[503:432];
logic [71:0] input_fmap_7;
assign input_fmap_7 = input_act_ff[575:504];
logic [71:0] input_fmap_8;
assign input_fmap_8 = input_act_ff[647:576];
logic [71:0] input_fmap_9;
assign input_fmap_9 = input_act_ff[719:648];
logic [71:0] input_fmap_10;
assign input_fmap_10 = input_act_ff[791:720];
logic [71:0] input_fmap_11;
assign input_fmap_11 = input_act_ff[863:792];
logic [71:0] input_fmap_12;
assign input_fmap_12 = input_act_ff[935:864];
logic [71:0] input_fmap_13;
assign input_fmap_13 = input_act_ff[1007:936];
logic [71:0] input_fmap_14;
assign input_fmap_14 = input_act_ff[1079:1008];
logic [71:0] input_fmap_15;
assign input_fmap_15 = input_act_ff[1151:1080];
logic [71:0] input_fmap_16;
assign input_fmap_16 = input_act_ff[1223:1152];
logic [71:0] input_fmap_17;
assign input_fmap_17 = input_act_ff[1295:1224];
logic [71:0] input_fmap_18;
assign input_fmap_18 = input_act_ff[1367:1296];
logic [71:0] input_fmap_19;
assign input_fmap_19 = input_act_ff[1439:1368];
logic [71:0] input_fmap_20;
assign input_fmap_20 = input_act_ff[1511:1440];
logic [71:0] input_fmap_21;
assign input_fmap_21 = input_act_ff[1583:1512];
logic [71:0] input_fmap_22;
assign input_fmap_22 = input_act_ff[1655:1584];
logic [71:0] input_fmap_23;
assign input_fmap_23 = input_act_ff[1727:1656];
logic [71:0] input_fmap_24;
assign input_fmap_24 = input_act_ff[1799:1728];
logic [71:0] input_fmap_25;
assign input_fmap_25 = input_act_ff[1871:1800];
logic [71:0] input_fmap_26;
assign input_fmap_26 = input_act_ff[1943:1872];
logic [71:0] input_fmap_27;
assign input_fmap_27 = input_act_ff[2015:1944];
logic [71:0] input_fmap_28;
assign input_fmap_28 = input_act_ff[2087:2016];
logic [71:0] input_fmap_29;
assign input_fmap_29 = input_act_ff[2159:2088];
logic [71:0] input_fmap_30;
assign input_fmap_30 = input_act_ff[2231:2160];
logic [71:0] input_fmap_31;
assign input_fmap_31 = input_act_ff[2303:2232];

logic [11-1:0] O0_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O0_I0_R0_C03_rom_inst (.q(O0_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O0_I0_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O0_I0_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O0_I0_R0_C03_rom_inst (.q(O0_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [13-1:0] O0_I0_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O0_I0_R0_C18_rom_inst (.q(O0_I0_R0_C1_SM1 ),.address(input_fmap_0[15:8]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R0_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O0_I0_R0_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O0_I0_R0_C18_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O0_I0_R0_C18_rom_inst (.q(O0_I0_R0_C1_SM1 ),.address(input_fmap_0[15:8]),.clock  (clk));
logic [12-1:0] O0_I0_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O0_I0_R0_C26_rom_inst (.q(O0_I0_R0_C2_SM1 ),.address(input_fmap_0[23:16]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R0_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O0_I0_R0_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O0_I0_R0_C26_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O0_I0_R0_C26_rom_inst (.q(O0_I0_R0_C2_SM1 ),.address(input_fmap_0[23:16]),.clock  (clk));
logic [15-1:0] O0_I0_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(15),.INIT_FILE("deepfreeze_rom/deepfreeze_8_15.txt"))
    conv5_dw_O0_I0_R1_C053_rom_inst (.q(O0_I0_R1_C0_SM1 ),.address(input_fmap_0[31:24]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R1_C0_SM1  = 15'h1234;
//always@(posedge clk) begin 
//O0_I0_R1_C0_SM1  <= 15'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O0_I0_R1_C053_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(15))
//    conv5_dw_O0_I0_R1_C053_rom_inst (.q(O0_I0_R1_C0_SM1 ),.address(input_fmap_0[31:24]),.clock  (clk));
logic [15-1:0] O0_I0_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(15),.INIT_FILE("deepfreeze_rom/deepfreeze_8_15.txt"))
    conv5_dw_O0_I0_R1_C150_rom_inst (.q(O0_I0_R1_C1_SM1 ),.address(input_fmap_0[39:32]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R1_C1_SM1  = 15'h1234;
//always@(posedge clk) begin 
//O0_I0_R1_C1_SM1  <= 15'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O0_I0_R1_C150_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(15))
//    conv5_dw_O0_I0_R1_C150_rom_inst (.q(O0_I0_R1_C1_SM1 ),.address(input_fmap_0[39:32]),.clock  (clk));
logic [10-1:0] O0_I0_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_dw_O0_I0_R1_C21_rom_inst (.q(O0_I0_R1_C2_SM1 ),.address(input_fmap_0[47:40]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R1_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O0_I0_R1_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O0_I0_R1_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_dw_O0_I0_R1_C21_rom_inst (.q(O0_I0_R1_C2_SM1 ),.address(input_fmap_0[47:40]),.clock  (clk));
logic [14-1:0] O0_I0_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv5_dw_O0_I0_R2_C016_rom_inst (.q(O0_I0_R2_C0_SM1 ),.address(input_fmap_0[55:48]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R2_C0_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O0_I0_R2_C0_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O0_I0_R2_C016_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv5_dw_O0_I0_R2_C016_rom_inst (.q(O0_I0_R2_C0_SM1 ),.address(input_fmap_0[55:48]),.clock  (clk));
logic [14-1:0] O0_I0_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv5_dw_O0_I0_R2_C116_rom_inst (.q(O0_I0_R2_C1_SM1 ),.address(input_fmap_0[63:56]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R2_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O0_I0_R2_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O0_I0_R2_C116_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv5_dw_O0_I0_R2_C116_rom_inst (.q(O0_I0_R2_C1_SM1 ),.address(input_fmap_0[63:56]),.clock  (clk));
logic [12-1:0] O0_I0_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O0_I0_R2_C25_rom_inst (.q(O0_I0_R2_C2_SM1 ),.address(input_fmap_0[71:64]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R2_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O0_I0_R2_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O0_I0_R2_C25_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O0_I0_R2_C25_rom_inst (.q(O0_I0_R2_C2_SM1 ),.address(input_fmap_0[71:64]),.clock  (clk));
logic [12-1:0] O1_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O1_I1_R0_C05_rom_inst (.q(O1_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O1_I1_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O1_I1_R0_C05_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O1_I1_R0_C05_rom_inst (.q(O1_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [13-1:0] O1_I1_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O1_I1_R0_C114_rom_inst (.q(O1_I1_R0_C1_SM1 ),.address(input_fmap_1[15:8]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R0_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O1_I1_R0_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O1_I1_R0_C114_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O1_I1_R0_C114_rom_inst (.q(O1_I1_R0_C1_SM1 ),.address(input_fmap_1[15:8]),.clock  (clk));
logic [11-1:0] O1_I1_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O1_I1_R0_C23_rom_inst (.q(O1_I1_R0_C2_SM1 ),.address(input_fmap_1[23:16]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R0_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O1_I1_R0_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O1_I1_R0_C23_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O1_I1_R0_C23_rom_inst (.q(O1_I1_R0_C2_SM1 ),.address(input_fmap_1[23:16]),.clock  (clk));
logic [13-1:0] O1_I1_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O1_I1_R1_C08_rom_inst (.q(O1_I1_R1_C0_SM1 ),.address(input_fmap_1[31:24]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R1_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O1_I1_R1_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O1_I1_R1_C08_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O1_I1_R1_C08_rom_inst (.q(O1_I1_R1_C0_SM1 ),.address(input_fmap_1[31:24]),.clock  (clk));
logic [15-1:0] O1_I1_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(15),.INIT_FILE("deepfreeze_rom/deepfreeze_8_15.txt"))
    conv5_dw_O1_I1_R1_C135_rom_inst (.q(O1_I1_R1_C1_SM1 ),.address(input_fmap_1[39:32]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R1_C1_SM1  = 15'h1234;
//always@(posedge clk) begin 
//O1_I1_R1_C1_SM1  <= 15'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O1_I1_R1_C135_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(15))
//    conv5_dw_O1_I1_R1_C135_rom_inst (.q(O1_I1_R1_C1_SM1 ),.address(input_fmap_1[39:32]),.clock  (clk));
logic [13-1:0] O1_I1_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O1_I1_R1_C212_rom_inst (.q(O1_I1_R1_C2_SM1 ),.address(input_fmap_1[47:40]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R1_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O1_I1_R1_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O1_I1_R1_C212_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O1_I1_R1_C212_rom_inst (.q(O1_I1_R1_C2_SM1 ),.address(input_fmap_1[47:40]),.clock  (clk));
logic [13-1:0] O1_I1_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O1_I1_R2_C09_rom_inst (.q(O1_I1_R2_C0_SM1 ),.address(input_fmap_1[55:48]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R2_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O1_I1_R2_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O1_I1_R2_C09_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O1_I1_R2_C09_rom_inst (.q(O1_I1_R2_C0_SM1 ),.address(input_fmap_1[55:48]),.clock  (clk));
logic [11-1:0] O1_I1_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O1_I1_R2_C12_rom_inst (.q(O1_I1_R2_C1_SM1 ),.address(input_fmap_1[63:56]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R2_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O1_I1_R2_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O1_I1_R2_C12_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O1_I1_R2_C12_rom_inst (.q(O1_I1_R2_C1_SM1 ),.address(input_fmap_1[63:56]),.clock  (clk));
logic [12-1:0] O1_I1_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O1_I1_R2_C24_rom_inst (.q(O1_I1_R2_C2_SM1 ),.address(input_fmap_1[71:64]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R2_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O1_I1_R2_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O1_I1_R2_C24_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O1_I1_R2_C24_rom_inst (.q(O1_I1_R2_C2_SM1 ),.address(input_fmap_1[71:64]),.clock  (clk));
logic [13-1:0] O2_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O2_I2_R0_C014_rom_inst (.q(O2_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O2_I2_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O2_I2_R0_C014_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O2_I2_R0_C014_rom_inst (.q(O2_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [13-1:0] O2_I2_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O2_I2_R0_C113_rom_inst (.q(O2_I2_R0_C1_SM1 ),.address(input_fmap_2[15:8]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R0_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O2_I2_R0_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O2_I2_R0_C113_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O2_I2_R0_C113_rom_inst (.q(O2_I2_R0_C1_SM1 ),.address(input_fmap_2[15:8]),.clock  (clk));
logic [11-1:0] O2_I2_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O2_I2_R0_C22_rom_inst (.q(O2_I2_R0_C2_SM1 ),.address(input_fmap_2[23:16]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R0_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O2_I2_R0_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O2_I2_R0_C22_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O2_I2_R0_C22_rom_inst (.q(O2_I2_R0_C2_SM1 ),.address(input_fmap_2[23:16]),.clock  (clk));
logic [12-1:0] O2_I2_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O2_I2_R1_C04_rom_inst (.q(O2_I2_R1_C0_SM1 ),.address(input_fmap_2[31:24]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R1_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O2_I2_R1_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O2_I2_R1_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O2_I2_R1_C04_rom_inst (.q(O2_I2_R1_C0_SM1 ),.address(input_fmap_2[31:24]),.clock  (clk));
logic [12-1:0] O2_I2_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O2_I2_R1_C14_rom_inst (.q(O2_I2_R1_C1_SM1 ),.address(input_fmap_2[39:32]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R1_C1_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O2_I2_R1_C1_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O2_I2_R1_C14_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O2_I2_R1_C14_rom_inst (.q(O2_I2_R1_C1_SM1 ),.address(input_fmap_2[39:32]),.clock  (clk));
logic [12-1:0] O2_I2_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O2_I2_R1_C27_rom_inst (.q(O2_I2_R1_C2_SM1 ),.address(input_fmap_2[47:40]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R1_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O2_I2_R1_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O2_I2_R1_C27_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O2_I2_R1_C27_rom_inst (.q(O2_I2_R1_C2_SM1 ),.address(input_fmap_2[47:40]),.clock  (clk));
logic [11-1:0] O2_I2_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O2_I2_R2_C02_rom_inst (.q(O2_I2_R2_C0_SM1 ),.address(input_fmap_2[55:48]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R2_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O2_I2_R2_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O2_I2_R2_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O2_I2_R2_C02_rom_inst (.q(O2_I2_R2_C0_SM1 ),.address(input_fmap_2[55:48]),.clock  (clk));
logic [12-1:0] O2_I2_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O2_I2_R2_C17_rom_inst (.q(O2_I2_R2_C1_SM1 ),.address(input_fmap_2[63:56]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R2_C1_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O2_I2_R2_C1_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O2_I2_R2_C17_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O2_I2_R2_C17_rom_inst (.q(O2_I2_R2_C1_SM1 ),.address(input_fmap_2[63:56]),.clock  (clk));
logic [11-1:0] O2_I2_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O2_I2_R2_C22_rom_inst (.q(O2_I2_R2_C2_SM1 ),.address(input_fmap_2[71:64]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R2_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O2_I2_R2_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O2_I2_R2_C22_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O2_I2_R2_C22_rom_inst (.q(O2_I2_R2_C2_SM1 ),.address(input_fmap_2[71:64]),.clock  (clk));
logic [10-1:0] O3_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_dw_O3_I3_R0_C01_rom_inst (.q(O3_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O3_I3_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O3_I3_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_dw_O3_I3_R0_C01_rom_inst (.q(O3_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [13-1:0] O3_I3_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O3_I3_R0_C18_rom_inst (.q(O3_I3_R0_C1_SM1 ),.address(input_fmap_3[15:8]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R0_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O3_I3_R0_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O3_I3_R0_C18_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O3_I3_R0_C18_rom_inst (.q(O3_I3_R0_C1_SM1 ),.address(input_fmap_3[15:8]),.clock  (clk));
logic [11-1:0] O3_I3_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O3_I3_R0_C22_rom_inst (.q(O3_I3_R0_C2_SM1 ),.address(input_fmap_3[23:16]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R0_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O3_I3_R0_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O3_I3_R0_C22_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O3_I3_R0_C22_rom_inst (.q(O3_I3_R0_C2_SM1 ),.address(input_fmap_3[23:16]),.clock  (clk));
logic [13-1:0] O3_I3_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O3_I3_R1_C09_rom_inst (.q(O3_I3_R1_C0_SM1 ),.address(input_fmap_3[31:24]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R1_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O3_I3_R1_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O3_I3_R1_C09_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O3_I3_R1_C09_rom_inst (.q(O3_I3_R1_C0_SM1 ),.address(input_fmap_3[31:24]),.clock  (clk));
logic [13-1:0] O3_I3_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O3_I3_R1_C112_rom_inst (.q(O3_I3_R1_C1_SM1 ),.address(input_fmap_3[39:32]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R1_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O3_I3_R1_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O3_I3_R1_C112_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O3_I3_R1_C112_rom_inst (.q(O3_I3_R1_C1_SM1 ),.address(input_fmap_3[39:32]),.clock  (clk));
logic [10-1:0] O3_I3_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_dw_O3_I3_R2_C01_rom_inst (.q(O3_I3_R2_C0_SM1 ),.address(input_fmap_3[55:48]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R2_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O3_I3_R2_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O3_I3_R2_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_dw_O3_I3_R2_C01_rom_inst (.q(O3_I3_R2_C0_SM1 ),.address(input_fmap_3[55:48]),.clock  (clk));
logic [13-1:0] O3_I3_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O3_I3_R2_C112_rom_inst (.q(O3_I3_R2_C1_SM1 ),.address(input_fmap_3[63:56]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R2_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O3_I3_R2_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O3_I3_R2_C112_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O3_I3_R2_C112_rom_inst (.q(O3_I3_R2_C1_SM1 ),.address(input_fmap_3[63:56]),.clock  (clk));
logic [10-1:0] O3_I3_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_dw_O3_I3_R2_C21_rom_inst (.q(O3_I3_R2_C2_SM1 ),.address(input_fmap_3[71:64]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R2_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O3_I3_R2_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O3_I3_R2_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_dw_O3_I3_R2_C21_rom_inst (.q(O3_I3_R2_C2_SM1 ),.address(input_fmap_3[71:64]),.clock  (clk));
logic [14-1:0] O4_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv5_dw_O4_I4_R0_C018_rom_inst (.q(O4_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R0_C0_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O4_I4_R0_C0_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O4_I4_R0_C018_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv5_dw_O4_I4_R0_C018_rom_inst (.q(O4_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [14-1:0] O4_I4_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv5_dw_O4_I4_R0_C117_rom_inst (.q(O4_I4_R0_C1_SM1 ),.address(input_fmap_4[15:8]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R0_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O4_I4_R0_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O4_I4_R0_C117_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv5_dw_O4_I4_R0_C117_rom_inst (.q(O4_I4_R0_C1_SM1 ),.address(input_fmap_4[15:8]),.clock  (clk));
logic [11-1:0] O4_I4_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O4_I4_R0_C22_rom_inst (.q(O4_I4_R0_C2_SM1 ),.address(input_fmap_4[23:16]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R0_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O4_I4_R0_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O4_I4_R0_C22_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O4_I4_R0_C22_rom_inst (.q(O4_I4_R0_C2_SM1 ),.address(input_fmap_4[23:16]),.clock  (clk));
logic [14-1:0] O4_I4_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv5_dw_O4_I4_R1_C017_rom_inst (.q(O4_I4_R1_C0_SM1 ),.address(input_fmap_4[31:24]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R1_C0_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O4_I4_R1_C0_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O4_I4_R1_C017_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv5_dw_O4_I4_R1_C017_rom_inst (.q(O4_I4_R1_C0_SM1 ),.address(input_fmap_4[31:24]),.clock  (clk));
logic [14-1:0] O4_I4_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv5_dw_O4_I4_R1_C120_rom_inst (.q(O4_I4_R1_C1_SM1 ),.address(input_fmap_4[39:32]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R1_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O4_I4_R1_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O4_I4_R1_C120_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv5_dw_O4_I4_R1_C120_rom_inst (.q(O4_I4_R1_C1_SM1 ),.address(input_fmap_4[39:32]),.clock  (clk));
logic [12-1:0] O4_I4_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O4_I4_R1_C27_rom_inst (.q(O4_I4_R1_C2_SM1 ),.address(input_fmap_4[47:40]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R1_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O4_I4_R1_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O4_I4_R1_C27_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O4_I4_R1_C27_rom_inst (.q(O4_I4_R1_C2_SM1 ),.address(input_fmap_4[47:40]),.clock  (clk));
logic [11-1:0] O4_I4_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O4_I4_R2_C03_rom_inst (.q(O4_I4_R2_C0_SM1 ),.address(input_fmap_4[55:48]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R2_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O4_I4_R2_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O4_I4_R2_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O4_I4_R2_C03_rom_inst (.q(O4_I4_R2_C0_SM1 ),.address(input_fmap_4[55:48]),.clock  (clk));
logic [11-1:0] O4_I4_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O4_I4_R2_C12_rom_inst (.q(O4_I4_R2_C1_SM1 ),.address(input_fmap_4[63:56]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R2_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O4_I4_R2_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O4_I4_R2_C12_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O4_I4_R2_C12_rom_inst (.q(O4_I4_R2_C1_SM1 ),.address(input_fmap_4[63:56]),.clock  (clk));
logic [11-1:0] O4_I4_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O4_I4_R2_C22_rom_inst (.q(O4_I4_R2_C2_SM1 ),.address(input_fmap_4[71:64]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R2_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O4_I4_R2_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O4_I4_R2_C22_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O4_I4_R2_C22_rom_inst (.q(O4_I4_R2_C2_SM1 ),.address(input_fmap_4[71:64]),.clock  (clk));
logic [11-1:0] O5_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O5_I5_R0_C02_rom_inst (.q(O5_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O5_I5_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O5_I5_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O5_I5_R0_C02_rom_inst (.q(O5_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [12-1:0] O5_I5_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O5_I5_R0_C14_rom_inst (.q(O5_I5_R0_C1_SM1 ),.address(input_fmap_5[15:8]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R0_C1_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O5_I5_R0_C1_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O5_I5_R0_C14_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O5_I5_R0_C14_rom_inst (.q(O5_I5_R0_C1_SM1 ),.address(input_fmap_5[15:8]),.clock  (clk));
logic [12-1:0] O5_I5_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O5_I5_R0_C25_rom_inst (.q(O5_I5_R0_C2_SM1 ),.address(input_fmap_5[23:16]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R0_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O5_I5_R0_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O5_I5_R0_C25_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O5_I5_R0_C25_rom_inst (.q(O5_I5_R0_C2_SM1 ),.address(input_fmap_5[23:16]),.clock  (clk));
logic [13-1:0] O5_I5_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O5_I5_R1_C012_rom_inst (.q(O5_I5_R1_C0_SM1 ),.address(input_fmap_5[31:24]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R1_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O5_I5_R1_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O5_I5_R1_C012_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O5_I5_R1_C012_rom_inst (.q(O5_I5_R1_C0_SM1 ),.address(input_fmap_5[31:24]),.clock  (clk));
logic [14-1:0] O5_I5_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv5_dw_O5_I5_R1_C129_rom_inst (.q(O5_I5_R1_C1_SM1 ),.address(input_fmap_5[39:32]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R1_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O5_I5_R1_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O5_I5_R1_C129_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv5_dw_O5_I5_R1_C129_rom_inst (.q(O5_I5_R1_C1_SM1 ),.address(input_fmap_5[39:32]),.clock  (clk));
logic [11-1:0] O5_I5_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O5_I5_R1_C22_rom_inst (.q(O5_I5_R1_C2_SM1 ),.address(input_fmap_5[47:40]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R1_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O5_I5_R1_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O5_I5_R1_C22_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O5_I5_R1_C22_rom_inst (.q(O5_I5_R1_C2_SM1 ),.address(input_fmap_5[47:40]),.clock  (clk));
logic [13-1:0] O5_I5_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O5_I5_R2_C013_rom_inst (.q(O5_I5_R2_C0_SM1 ),.address(input_fmap_5[55:48]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R2_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O5_I5_R2_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O5_I5_R2_C013_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O5_I5_R2_C013_rom_inst (.q(O5_I5_R2_C0_SM1 ),.address(input_fmap_5[55:48]),.clock  (clk));
logic [14-1:0] O5_I5_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv5_dw_O5_I5_R2_C124_rom_inst (.q(O5_I5_R2_C1_SM1 ),.address(input_fmap_5[63:56]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R2_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O5_I5_R2_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O5_I5_R2_C124_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv5_dw_O5_I5_R2_C124_rom_inst (.q(O5_I5_R2_C1_SM1 ),.address(input_fmap_5[63:56]),.clock  (clk));
logic [10-1:0] O5_I5_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_dw_O5_I5_R2_C21_rom_inst (.q(O5_I5_R2_C2_SM1 ),.address(input_fmap_5[71:64]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R2_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I5_R2_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O5_I5_R2_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_dw_O5_I5_R2_C21_rom_inst (.q(O5_I5_R2_C2_SM1 ),.address(input_fmap_5[71:64]),.clock  (clk));
logic [13-1:0] O6_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O6_I6_R0_C013_rom_inst (.q(O6_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O6_I6_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O6_I6_R0_C013_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O6_I6_R0_C013_rom_inst (.q(O6_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [14-1:0] O6_I6_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv5_dw_O6_I6_R0_C119_rom_inst (.q(O6_I6_R0_C1_SM1 ),.address(input_fmap_6[15:8]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R0_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O6_I6_R0_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O6_I6_R0_C119_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv5_dw_O6_I6_R0_C119_rom_inst (.q(O6_I6_R0_C1_SM1 ),.address(input_fmap_6[15:8]),.clock  (clk));
logic [12-1:0] O6_I6_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O6_I6_R0_C27_rom_inst (.q(O6_I6_R0_C2_SM1 ),.address(input_fmap_6[23:16]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R0_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O6_I6_R0_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O6_I6_R0_C27_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O6_I6_R0_C27_rom_inst (.q(O6_I6_R0_C2_SM1 ),.address(input_fmap_6[23:16]),.clock  (clk));
logic [14-1:0] O6_I6_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv5_dw_O6_I6_R1_C022_rom_inst (.q(O6_I6_R1_C0_SM1 ),.address(input_fmap_6[31:24]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R1_C0_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O6_I6_R1_C0_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O6_I6_R1_C022_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv5_dw_O6_I6_R1_C022_rom_inst (.q(O6_I6_R1_C0_SM1 ),.address(input_fmap_6[31:24]),.clock  (clk));
logic [14-1:0] O6_I6_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv5_dw_O6_I6_R1_C129_rom_inst (.q(O6_I6_R1_C1_SM1 ),.address(input_fmap_6[39:32]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R1_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O6_I6_R1_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O6_I6_R1_C129_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv5_dw_O6_I6_R1_C129_rom_inst (.q(O6_I6_R1_C1_SM1 ),.address(input_fmap_6[39:32]),.clock  (clk));
logic [13-1:0] O6_I6_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O6_I6_R1_C28_rom_inst (.q(O6_I6_R1_C2_SM1 ),.address(input_fmap_6[47:40]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R1_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O6_I6_R1_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O6_I6_R1_C28_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O6_I6_R1_C28_rom_inst (.q(O6_I6_R1_C2_SM1 ),.address(input_fmap_6[47:40]),.clock  (clk));
logic [13-1:0] O6_I6_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O6_I6_R2_C012_rom_inst (.q(O6_I6_R2_C0_SM1 ),.address(input_fmap_6[55:48]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R2_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O6_I6_R2_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O6_I6_R2_C012_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O6_I6_R2_C012_rom_inst (.q(O6_I6_R2_C0_SM1 ),.address(input_fmap_6[55:48]),.clock  (clk));
logic [13-1:0] O6_I6_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O6_I6_R2_C110_rom_inst (.q(O6_I6_R2_C1_SM1 ),.address(input_fmap_6[63:56]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R2_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O6_I6_R2_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O6_I6_R2_C110_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O6_I6_R2_C110_rom_inst (.q(O6_I6_R2_C1_SM1 ),.address(input_fmap_6[63:56]),.clock  (clk));
logic [10-1:0] O6_I6_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_dw_O6_I6_R2_C21_rom_inst (.q(O6_I6_R2_C2_SM1 ),.address(input_fmap_6[71:64]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R2_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O6_I6_R2_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O6_I6_R2_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_dw_O6_I6_R2_C21_rom_inst (.q(O6_I6_R2_C2_SM1 ),.address(input_fmap_6[71:64]),.clock  (clk));
logic [10-1:0] O7_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_dw_O7_I7_R0_C01_rom_inst (.q(O7_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O7_I7_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O7_I7_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_dw_O7_I7_R0_C01_rom_inst (.q(O7_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [14-1:0] O7_I7_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv5_dw_O7_I7_R0_C119_rom_inst (.q(O7_I7_R0_C1_SM1 ),.address(input_fmap_7[15:8]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R0_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O7_I7_R0_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O7_I7_R0_C119_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv5_dw_O7_I7_R0_C119_rom_inst (.q(O7_I7_R0_C1_SM1 ),.address(input_fmap_7[15:8]),.clock  (clk));
logic [10-1:0] O7_I7_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_dw_O7_I7_R0_C21_rom_inst (.q(O7_I7_R0_C2_SM1 ),.address(input_fmap_7[23:16]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R0_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O7_I7_R0_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O7_I7_R0_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_dw_O7_I7_R0_C21_rom_inst (.q(O7_I7_R0_C2_SM1 ),.address(input_fmap_7[23:16]),.clock  (clk));
logic [13-1:0] O7_I7_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O7_I7_R1_C015_rom_inst (.q(O7_I7_R1_C0_SM1 ),.address(input_fmap_7[31:24]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R1_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O7_I7_R1_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O7_I7_R1_C015_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O7_I7_R1_C015_rom_inst (.q(O7_I7_R1_C0_SM1 ),.address(input_fmap_7[31:24]),.clock  (clk));
logic [13-1:0] O7_I7_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O7_I7_R1_C113_rom_inst (.q(O7_I7_R1_C1_SM1 ),.address(input_fmap_7[39:32]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R1_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O7_I7_R1_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O7_I7_R1_C113_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O7_I7_R1_C113_rom_inst (.q(O7_I7_R1_C1_SM1 ),.address(input_fmap_7[39:32]),.clock  (clk));
logic [11-1:0] O7_I7_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O7_I7_R1_C23_rom_inst (.q(O7_I7_R1_C2_SM1 ),.address(input_fmap_7[47:40]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R1_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O7_I7_R1_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O7_I7_R1_C23_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O7_I7_R1_C23_rom_inst (.q(O7_I7_R1_C2_SM1 ),.address(input_fmap_7[47:40]),.clock  (clk));
logic [10-1:0] O7_I7_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_dw_O7_I7_R2_C01_rom_inst (.q(O7_I7_R2_C0_SM1 ),.address(input_fmap_7[55:48]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R2_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O7_I7_R2_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O7_I7_R2_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_dw_O7_I7_R2_C01_rom_inst (.q(O7_I7_R2_C0_SM1 ),.address(input_fmap_7[55:48]),.clock  (clk));
logic [12-1:0] O7_I7_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O7_I7_R2_C15_rom_inst (.q(O7_I7_R2_C1_SM1 ),.address(input_fmap_7[63:56]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R2_C1_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O7_I7_R2_C1_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O7_I7_R2_C15_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O7_I7_R2_C15_rom_inst (.q(O7_I7_R2_C1_SM1 ),.address(input_fmap_7[63:56]),.clock  (clk));
logic [12-1:0] O7_I7_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O7_I7_R2_C26_rom_inst (.q(O7_I7_R2_C2_SM1 ),.address(input_fmap_7[71:64]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R2_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O7_I7_R2_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O7_I7_R2_C26_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O7_I7_R2_C26_rom_inst (.q(O7_I7_R2_C2_SM1 ),.address(input_fmap_7[71:64]),.clock  (clk));
logic [14-1:0] O8_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv5_dw_O8_I8_R0_C024_rom_inst (.q(O8_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O8_I8_R0_C0_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O8_I8_R0_C0_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O8_I8_R0_C024_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv5_dw_O8_I8_R0_C024_rom_inst (.q(O8_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [14-1:0] O8_I8_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv5_dw_O8_I8_R0_C121_rom_inst (.q(O8_I8_R0_C1_SM1 ),.address(input_fmap_8[15:8]),.clk(clk),.d(0),.we(0));
//assign O8_I8_R0_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O8_I8_R0_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O8_I8_R0_C121_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv5_dw_O8_I8_R0_C121_rom_inst (.q(O8_I8_R0_C1_SM1 ),.address(input_fmap_8[15:8]),.clock  (clk));
logic [12-1:0] O8_I8_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O8_I8_R0_C26_rom_inst (.q(O8_I8_R0_C2_SM1 ),.address(input_fmap_8[23:16]),.clk(clk),.d(0),.we(0));
//assign O8_I8_R0_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O8_I8_R0_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O8_I8_R0_C26_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O8_I8_R0_C26_rom_inst (.q(O8_I8_R0_C2_SM1 ),.address(input_fmap_8[23:16]),.clock  (clk));
logic [14-1:0] O8_I8_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv5_dw_O8_I8_R1_C023_rom_inst (.q(O8_I8_R1_C0_SM1 ),.address(input_fmap_8[31:24]),.clk(clk),.d(0),.we(0));
//assign O8_I8_R1_C0_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O8_I8_R1_C0_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O8_I8_R1_C023_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv5_dw_O8_I8_R1_C023_rom_inst (.q(O8_I8_R1_C0_SM1 ),.address(input_fmap_8[31:24]),.clock  (clk));
logic [14-1:0] O8_I8_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv5_dw_O8_I8_R1_C131_rom_inst (.q(O8_I8_R1_C1_SM1 ),.address(input_fmap_8[39:32]),.clk(clk),.d(0),.we(0));
//assign O8_I8_R1_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O8_I8_R1_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O8_I8_R1_C131_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv5_dw_O8_I8_R1_C131_rom_inst (.q(O8_I8_R1_C1_SM1 ),.address(input_fmap_8[39:32]),.clock  (clk));
logic [13-1:0] O8_I8_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O8_I8_R2_C012_rom_inst (.q(O8_I8_R2_C0_SM1 ),.address(input_fmap_8[55:48]),.clk(clk),.d(0),.we(0));
//assign O8_I8_R2_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O8_I8_R2_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O8_I8_R2_C012_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O8_I8_R2_C012_rom_inst (.q(O8_I8_R2_C0_SM1 ),.address(input_fmap_8[55:48]),.clock  (clk));
logic [10-1:0] O8_I8_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_dw_O8_I8_R2_C11_rom_inst (.q(O8_I8_R2_C1_SM1 ),.address(input_fmap_8[63:56]),.clk(clk),.d(0),.we(0));
//assign O8_I8_R2_C1_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O8_I8_R2_C1_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O8_I8_R2_C11_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_dw_O8_I8_R2_C11_rom_inst (.q(O8_I8_R2_C1_SM1 ),.address(input_fmap_8[63:56]),.clock  (clk));
logic [11-1:0] O8_I8_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O8_I8_R2_C23_rom_inst (.q(O8_I8_R2_C2_SM1 ),.address(input_fmap_8[71:64]),.clk(clk),.d(0),.we(0));
//assign O8_I8_R2_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O8_I8_R2_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O8_I8_R2_C23_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O8_I8_R2_C23_rom_inst (.q(O8_I8_R2_C2_SM1 ),.address(input_fmap_8[71:64]),.clock  (clk));
logic [12-1:0] O9_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O9_I9_R0_C06_rom_inst (.q(O9_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O9_I9_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O9_I9_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O9_I9_R0_C06_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O9_I9_R0_C06_rom_inst (.q(O9_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [11-1:0] O9_I9_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O9_I9_R0_C13_rom_inst (.q(O9_I9_R0_C1_SM1 ),.address(input_fmap_9[15:8]),.clk(clk),.d(0),.we(0));
//assign O9_I9_R0_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O9_I9_R0_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O9_I9_R0_C13_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O9_I9_R0_C13_rom_inst (.q(O9_I9_R0_C1_SM1 ),.address(input_fmap_9[15:8]),.clock  (clk));
logic [11-1:0] O9_I9_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O9_I9_R0_C23_rom_inst (.q(O9_I9_R0_C2_SM1 ),.address(input_fmap_9[23:16]),.clk(clk),.d(0),.we(0));
//assign O9_I9_R0_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O9_I9_R0_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O9_I9_R0_C23_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O9_I9_R0_C23_rom_inst (.q(O9_I9_R0_C2_SM1 ),.address(input_fmap_9[23:16]),.clock  (clk));
logic [14-1:0] O9_I9_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv5_dw_O9_I9_R1_C017_rom_inst (.q(O9_I9_R1_C0_SM1 ),.address(input_fmap_9[31:24]),.clk(clk),.d(0),.we(0));
//assign O9_I9_R1_C0_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O9_I9_R1_C0_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O9_I9_R1_C017_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv5_dw_O9_I9_R1_C017_rom_inst (.q(O9_I9_R1_C0_SM1 ),.address(input_fmap_9[31:24]),.clock  (clk));
logic [13-1:0] O9_I9_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O9_I9_R1_C113_rom_inst (.q(O9_I9_R1_C1_SM1 ),.address(input_fmap_9[39:32]),.clk(clk),.d(0),.we(0));
//assign O9_I9_R1_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O9_I9_R1_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O9_I9_R1_C113_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O9_I9_R1_C113_rom_inst (.q(O9_I9_R1_C1_SM1 ),.address(input_fmap_9[39:32]),.clock  (clk));
logic [10-1:0] O9_I9_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_dw_O9_I9_R1_C21_rom_inst (.q(O9_I9_R1_C2_SM1 ),.address(input_fmap_9[47:40]),.clk(clk),.d(0),.we(0));
//assign O9_I9_R1_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O9_I9_R1_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O9_I9_R1_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_dw_O9_I9_R1_C21_rom_inst (.q(O9_I9_R1_C2_SM1 ),.address(input_fmap_9[47:40]),.clock  (clk));
logic [12-1:0] O9_I9_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O9_I9_R2_C06_rom_inst (.q(O9_I9_R2_C0_SM1 ),.address(input_fmap_9[55:48]),.clk(clk),.d(0),.we(0));
//assign O9_I9_R2_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O9_I9_R2_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O9_I9_R2_C06_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O9_I9_R2_C06_rom_inst (.q(O9_I9_R2_C0_SM1 ),.address(input_fmap_9[55:48]),.clock  (clk));
logic [12-1:0] O9_I9_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O9_I9_R2_C17_rom_inst (.q(O9_I9_R2_C1_SM1 ),.address(input_fmap_9[63:56]),.clk(clk),.d(0),.we(0));
//assign O9_I9_R2_C1_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O9_I9_R2_C1_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O9_I9_R2_C17_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O9_I9_R2_C17_rom_inst (.q(O9_I9_R2_C1_SM1 ),.address(input_fmap_9[63:56]),.clock  (clk));
logic [11-1:0] O9_I9_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O9_I9_R2_C23_rom_inst (.q(O9_I9_R2_C2_SM1 ),.address(input_fmap_9[71:64]),.clk(clk),.d(0),.we(0));
//assign O9_I9_R2_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O9_I9_R2_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O9_I9_R2_C23_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O9_I9_R2_C23_rom_inst (.q(O9_I9_R2_C2_SM1 ),.address(input_fmap_9[71:64]),.clock  (clk));
logic [13-1:0] O10_I10_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O10_I10_R0_C012_rom_inst (.q(O10_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clk(clk),.d(0),.we(0));
//assign O10_I10_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O10_I10_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O10_I10_R0_C012_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O10_I10_R0_C012_rom_inst (.q(O10_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clock  (clk));
logic [12-1:0] O10_I10_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O10_I10_R0_C15_rom_inst (.q(O10_I10_R0_C1_SM1 ),.address(input_fmap_10[15:8]),.clk(clk),.d(0),.we(0));
//assign O10_I10_R0_C1_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O10_I10_R0_C1_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O10_I10_R0_C15_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O10_I10_R0_C15_rom_inst (.q(O10_I10_R0_C1_SM1 ),.address(input_fmap_10[15:8]),.clock  (clk));
logic [11-1:0] O10_I10_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O10_I10_R0_C23_rom_inst (.q(O10_I10_R0_C2_SM1 ),.address(input_fmap_10[23:16]),.clk(clk),.d(0),.we(0));
//assign O10_I10_R0_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O10_I10_R0_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O10_I10_R0_C23_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O10_I10_R0_C23_rom_inst (.q(O10_I10_R0_C2_SM1 ),.address(input_fmap_10[23:16]),.clock  (clk));
logic [14-1:0] O10_I10_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv5_dw_O10_I10_R1_C018_rom_inst (.q(O10_I10_R1_C0_SM1 ),.address(input_fmap_10[31:24]),.clk(clk),.d(0),.we(0));
//assign O10_I10_R1_C0_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O10_I10_R1_C0_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O10_I10_R1_C018_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv5_dw_O10_I10_R1_C018_rom_inst (.q(O10_I10_R1_C0_SM1 ),.address(input_fmap_10[31:24]),.clock  (clk));
logic [14-1:0] O10_I10_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv5_dw_O10_I10_R1_C127_rom_inst (.q(O10_I10_R1_C1_SM1 ),.address(input_fmap_10[39:32]),.clk(clk),.d(0),.we(0));
//assign O10_I10_R1_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O10_I10_R1_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O10_I10_R1_C127_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv5_dw_O10_I10_R1_C127_rom_inst (.q(O10_I10_R1_C1_SM1 ),.address(input_fmap_10[39:32]),.clock  (clk));
logic [13-1:0] O10_I10_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O10_I10_R1_C215_rom_inst (.q(O10_I10_R1_C2_SM1 ),.address(input_fmap_10[47:40]),.clk(clk),.d(0),.we(0));
//assign O10_I10_R1_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O10_I10_R1_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O10_I10_R1_C215_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O10_I10_R1_C215_rom_inst (.q(O10_I10_R1_C2_SM1 ),.address(input_fmap_10[47:40]),.clock  (clk));
logic [12-1:0] O10_I10_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O10_I10_R2_C05_rom_inst (.q(O10_I10_R2_C0_SM1 ),.address(input_fmap_10[55:48]),.clk(clk),.d(0),.we(0));
//assign O10_I10_R2_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O10_I10_R2_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O10_I10_R2_C05_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O10_I10_R2_C05_rom_inst (.q(O10_I10_R2_C0_SM1 ),.address(input_fmap_10[55:48]),.clock  (clk));
logic [13-1:0] O10_I10_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O10_I10_R2_C19_rom_inst (.q(O10_I10_R2_C1_SM1 ),.address(input_fmap_10[63:56]),.clk(clk),.d(0),.we(0));
//assign O10_I10_R2_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O10_I10_R2_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O10_I10_R2_C19_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O10_I10_R2_C19_rom_inst (.q(O10_I10_R2_C1_SM1 ),.address(input_fmap_10[63:56]),.clock  (clk));
logic [13-1:0] O10_I10_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O10_I10_R2_C210_rom_inst (.q(O10_I10_R2_C2_SM1 ),.address(input_fmap_10[71:64]),.clk(clk),.d(0),.we(0));
//assign O10_I10_R2_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O10_I10_R2_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O10_I10_R2_C210_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O10_I10_R2_C210_rom_inst (.q(O10_I10_R2_C2_SM1 ),.address(input_fmap_10[71:64]),.clock  (clk));
logic [13-1:0] O11_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O11_I11_R0_C010_rom_inst (.q(O11_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I11_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O11_I11_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O11_I11_R0_C010_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O11_I11_R0_C010_rom_inst (.q(O11_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [11-1:0] O11_I11_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O11_I11_R0_C23_rom_inst (.q(O11_I11_R0_C2_SM1 ),.address(input_fmap_11[23:16]),.clk(clk),.d(0),.we(0));
//assign O11_I11_R0_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O11_I11_R0_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O11_I11_R0_C23_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O11_I11_R0_C23_rom_inst (.q(O11_I11_R0_C2_SM1 ),.address(input_fmap_11[23:16]),.clock  (clk));
logic [14-1:0] O11_I11_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv5_dw_O11_I11_R1_C023_rom_inst (.q(O11_I11_R1_C0_SM1 ),.address(input_fmap_11[31:24]),.clk(clk),.d(0),.we(0));
//assign O11_I11_R1_C0_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O11_I11_R1_C0_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O11_I11_R1_C023_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv5_dw_O11_I11_R1_C023_rom_inst (.q(O11_I11_R1_C0_SM1 ),.address(input_fmap_11[31:24]),.clock  (clk));
logic [14-1:0] O11_I11_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv5_dw_O11_I11_R1_C130_rom_inst (.q(O11_I11_R1_C1_SM1 ),.address(input_fmap_11[39:32]),.clk(clk),.d(0),.we(0));
//assign O11_I11_R1_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O11_I11_R1_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O11_I11_R1_C130_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv5_dw_O11_I11_R1_C130_rom_inst (.q(O11_I11_R1_C1_SM1 ),.address(input_fmap_11[39:32]),.clock  (clk));
logic [13-1:0] O11_I11_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O11_I11_R1_C28_rom_inst (.q(O11_I11_R1_C2_SM1 ),.address(input_fmap_11[47:40]),.clk(clk),.d(0),.we(0));
//assign O11_I11_R1_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O11_I11_R1_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O11_I11_R1_C28_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O11_I11_R1_C28_rom_inst (.q(O11_I11_R1_C2_SM1 ),.address(input_fmap_11[47:40]),.clock  (clk));
logic [11-1:0] O11_I11_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O11_I11_R2_C03_rom_inst (.q(O11_I11_R2_C0_SM1 ),.address(input_fmap_11[55:48]),.clk(clk),.d(0),.we(0));
//assign O11_I11_R2_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O11_I11_R2_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O11_I11_R2_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O11_I11_R2_C03_rom_inst (.q(O11_I11_R2_C0_SM1 ),.address(input_fmap_11[55:48]),.clock  (clk));
logic [11-1:0] O11_I11_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O11_I11_R2_C13_rom_inst (.q(O11_I11_R2_C1_SM1 ),.address(input_fmap_11[63:56]),.clk(clk),.d(0),.we(0));
//assign O11_I11_R2_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O11_I11_R2_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O11_I11_R2_C13_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O11_I11_R2_C13_rom_inst (.q(O11_I11_R2_C1_SM1 ),.address(input_fmap_11[63:56]),.clock  (clk));
logic [12-1:0] O11_I11_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O11_I11_R2_C25_rom_inst (.q(O11_I11_R2_C2_SM1 ),.address(input_fmap_11[71:64]),.clk(clk),.d(0),.we(0));
//assign O11_I11_R2_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O11_I11_R2_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O11_I11_R2_C25_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O11_I11_R2_C25_rom_inst (.q(O11_I11_R2_C2_SM1 ),.address(input_fmap_11[71:64]),.clock  (clk));
logic [12-1:0] O12_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O12_I12_R0_C04_rom_inst (.q(O12_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I12_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O12_I12_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O12_I12_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O12_I12_R0_C04_rom_inst (.q(O12_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [13-1:0] O12_I12_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O12_I12_R0_C115_rom_inst (.q(O12_I12_R0_C1_SM1 ),.address(input_fmap_12[15:8]),.clk(clk),.d(0),.we(0));
//assign O12_I12_R0_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O12_I12_R0_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O12_I12_R0_C115_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O12_I12_R0_C115_rom_inst (.q(O12_I12_R0_C1_SM1 ),.address(input_fmap_12[15:8]),.clock  (clk));
logic [12-1:0] O12_I12_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O12_I12_R0_C24_rom_inst (.q(O12_I12_R0_C2_SM1 ),.address(input_fmap_12[23:16]),.clk(clk),.d(0),.we(0));
//assign O12_I12_R0_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O12_I12_R0_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O12_I12_R0_C24_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O12_I12_R0_C24_rom_inst (.q(O12_I12_R0_C2_SM1 ),.address(input_fmap_12[23:16]),.clock  (clk));
logic [13-1:0] O12_I12_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O12_I12_R1_C014_rom_inst (.q(O12_I12_R1_C0_SM1 ),.address(input_fmap_12[31:24]),.clk(clk),.d(0),.we(0));
//assign O12_I12_R1_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O12_I12_R1_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O12_I12_R1_C014_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O12_I12_R1_C014_rom_inst (.q(O12_I12_R1_C0_SM1 ),.address(input_fmap_12[31:24]),.clock  (clk));
logic [14-1:0] O12_I12_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv5_dw_O12_I12_R1_C129_rom_inst (.q(O12_I12_R1_C1_SM1 ),.address(input_fmap_12[39:32]),.clk(clk),.d(0),.we(0));
//assign O12_I12_R1_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O12_I12_R1_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O12_I12_R1_C129_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv5_dw_O12_I12_R1_C129_rom_inst (.q(O12_I12_R1_C1_SM1 ),.address(input_fmap_12[39:32]),.clock  (clk));
logic [10-1:0] O12_I12_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_dw_O12_I12_R1_C21_rom_inst (.q(O12_I12_R1_C2_SM1 ),.address(input_fmap_12[47:40]),.clk(clk),.d(0),.we(0));
//assign O12_I12_R1_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O12_I12_R1_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O12_I12_R1_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_dw_O12_I12_R1_C21_rom_inst (.q(O12_I12_R1_C2_SM1 ),.address(input_fmap_12[47:40]),.clock  (clk));
logic [13-1:0] O12_I12_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O12_I12_R2_C012_rom_inst (.q(O12_I12_R2_C0_SM1 ),.address(input_fmap_12[55:48]),.clk(clk),.d(0),.we(0));
//assign O12_I12_R2_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O12_I12_R2_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O12_I12_R2_C012_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O12_I12_R2_C012_rom_inst (.q(O12_I12_R2_C0_SM1 ),.address(input_fmap_12[55:48]),.clock  (clk));
logic [11-1:0] O12_I12_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O12_I12_R2_C13_rom_inst (.q(O12_I12_R2_C1_SM1 ),.address(input_fmap_12[63:56]),.clk(clk),.d(0),.we(0));
//assign O12_I12_R2_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O12_I12_R2_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O12_I12_R2_C13_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O12_I12_R2_C13_rom_inst (.q(O12_I12_R2_C1_SM1 ),.address(input_fmap_12[63:56]),.clock  (clk));
logic [12-1:0] O12_I12_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O12_I12_R2_C27_rom_inst (.q(O12_I12_R2_C2_SM1 ),.address(input_fmap_12[71:64]),.clk(clk),.d(0),.we(0));
//assign O12_I12_R2_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O12_I12_R2_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O12_I12_R2_C27_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O12_I12_R2_C27_rom_inst (.q(O12_I12_R2_C2_SM1 ),.address(input_fmap_12[71:64]),.clock  (clk));
logic [13-1:0] O13_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O13_I13_R0_C015_rom_inst (.q(O13_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O13_I13_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O13_I13_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O13_I13_R0_C015_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O13_I13_R0_C015_rom_inst (.q(O13_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [14-1:0] O13_I13_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv5_dw_O13_I13_R0_C117_rom_inst (.q(O13_I13_R0_C1_SM1 ),.address(input_fmap_13[15:8]),.clk(clk),.d(0),.we(0));
//assign O13_I13_R0_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O13_I13_R0_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O13_I13_R0_C117_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv5_dw_O13_I13_R0_C117_rom_inst (.q(O13_I13_R0_C1_SM1 ),.address(input_fmap_13[15:8]),.clock  (clk));
logic [11-1:0] O13_I13_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O13_I13_R0_C23_rom_inst (.q(O13_I13_R0_C2_SM1 ),.address(input_fmap_13[23:16]),.clk(clk),.d(0),.we(0));
//assign O13_I13_R0_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O13_I13_R0_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O13_I13_R0_C23_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O13_I13_R0_C23_rom_inst (.q(O13_I13_R0_C2_SM1 ),.address(input_fmap_13[23:16]),.clock  (clk));
logic [15-1:0] O13_I13_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(15),.INIT_FILE("deepfreeze_rom/deepfreeze_8_15.txt"))
    conv5_dw_O13_I13_R1_C040_rom_inst (.q(O13_I13_R1_C0_SM1 ),.address(input_fmap_13[31:24]),.clk(clk),.d(0),.we(0));
//assign O13_I13_R1_C0_SM1  = 15'h1234;
//always@(posedge clk) begin 
//O13_I13_R1_C0_SM1  <= 15'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O13_I13_R1_C040_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(15))
//    conv5_dw_O13_I13_R1_C040_rom_inst (.q(O13_I13_R1_C0_SM1 ),.address(input_fmap_13[31:24]),.clock  (clk));
logic [14-1:0] O13_I13_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv5_dw_O13_I13_R1_C129_rom_inst (.q(O13_I13_R1_C1_SM1 ),.address(input_fmap_13[39:32]),.clk(clk),.d(0),.we(0));
//assign O13_I13_R1_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O13_I13_R1_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O13_I13_R1_C129_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv5_dw_O13_I13_R1_C129_rom_inst (.q(O13_I13_R1_C1_SM1 ),.address(input_fmap_13[39:32]),.clock  (clk));
logic [13-1:0] O13_I13_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O13_I13_R1_C211_rom_inst (.q(O13_I13_R1_C2_SM1 ),.address(input_fmap_13[47:40]),.clk(clk),.d(0),.we(0));
//assign O13_I13_R1_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O13_I13_R1_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O13_I13_R1_C211_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O13_I13_R1_C211_rom_inst (.q(O13_I13_R1_C2_SM1 ),.address(input_fmap_13[47:40]),.clock  (clk));
logic [13-1:0] O13_I13_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O13_I13_R2_C013_rom_inst (.q(O13_I13_R2_C0_SM1 ),.address(input_fmap_13[55:48]),.clk(clk),.d(0),.we(0));
//assign O13_I13_R2_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O13_I13_R2_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O13_I13_R2_C013_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O13_I13_R2_C013_rom_inst (.q(O13_I13_R2_C0_SM1 ),.address(input_fmap_13[55:48]),.clock  (clk));
logic [13-1:0] O13_I13_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O13_I13_R2_C19_rom_inst (.q(O13_I13_R2_C1_SM1 ),.address(input_fmap_13[63:56]),.clk(clk),.d(0),.we(0));
//assign O13_I13_R2_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O13_I13_R2_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O13_I13_R2_C19_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O13_I13_R2_C19_rom_inst (.q(O13_I13_R2_C1_SM1 ),.address(input_fmap_13[63:56]),.clock  (clk));
logic [13-1:0] O13_I13_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O13_I13_R2_C28_rom_inst (.q(O13_I13_R2_C2_SM1 ),.address(input_fmap_13[71:64]),.clk(clk),.d(0),.we(0));
//assign O13_I13_R2_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O13_I13_R2_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O13_I13_R2_C28_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O13_I13_R2_C28_rom_inst (.q(O13_I13_R2_C2_SM1 ),.address(input_fmap_13[71:64]),.clock  (clk));
logic [14-1:0] O14_I14_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv5_dw_O14_I14_R0_C118_rom_inst (.q(O14_I14_R0_C1_SM1 ),.address(input_fmap_14[15:8]),.clk(clk),.d(0),.we(0));
//assign O14_I14_R0_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O14_I14_R0_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O14_I14_R0_C118_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv5_dw_O14_I14_R0_C118_rom_inst (.q(O14_I14_R0_C1_SM1 ),.address(input_fmap_14[15:8]),.clock  (clk));
logic [10-1:0] O14_I14_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_dw_O14_I14_R0_C21_rom_inst (.q(O14_I14_R0_C2_SM1 ),.address(input_fmap_14[23:16]),.clk(clk),.d(0),.we(0));
//assign O14_I14_R0_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O14_I14_R0_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O14_I14_R0_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_dw_O14_I14_R0_C21_rom_inst (.q(O14_I14_R0_C2_SM1 ),.address(input_fmap_14[23:16]),.clock  (clk));
logic [12-1:0] O14_I14_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O14_I14_R1_C06_rom_inst (.q(O14_I14_R1_C0_SM1 ),.address(input_fmap_14[31:24]),.clk(clk),.d(0),.we(0));
//assign O14_I14_R1_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O14_I14_R1_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O14_I14_R1_C06_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O14_I14_R1_C06_rom_inst (.q(O14_I14_R1_C0_SM1 ),.address(input_fmap_14[31:24]),.clock  (clk));
logic [15-1:0] O14_I14_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(15),.INIT_FILE("deepfreeze_rom/deepfreeze_8_15.txt"))
    conv5_dw_O14_I14_R1_C144_rom_inst (.q(O14_I14_R1_C1_SM1 ),.address(input_fmap_14[39:32]),.clk(clk),.d(0),.we(0));
//assign O14_I14_R1_C1_SM1  = 15'h1234;
//always@(posedge clk) begin 
//O14_I14_R1_C1_SM1  <= 15'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O14_I14_R1_C144_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(15))
//    conv5_dw_O14_I14_R1_C144_rom_inst (.q(O14_I14_R1_C1_SM1 ),.address(input_fmap_14[39:32]),.clock  (clk));
logic [13-1:0] O14_I14_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O14_I14_R1_C28_rom_inst (.q(O14_I14_R1_C2_SM1 ),.address(input_fmap_14[47:40]),.clk(clk),.d(0),.we(0));
//assign O14_I14_R1_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O14_I14_R1_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O14_I14_R1_C28_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O14_I14_R1_C28_rom_inst (.q(O14_I14_R1_C2_SM1 ),.address(input_fmap_14[47:40]),.clock  (clk));
logic [13-1:0] O14_I14_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O14_I14_R2_C08_rom_inst (.q(O14_I14_R2_C0_SM1 ),.address(input_fmap_14[55:48]),.clk(clk),.d(0),.we(0));
//assign O14_I14_R2_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O14_I14_R2_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O14_I14_R2_C08_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O14_I14_R2_C08_rom_inst (.q(O14_I14_R2_C0_SM1 ),.address(input_fmap_14[55:48]),.clock  (clk));
logic [13-1:0] O14_I14_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O14_I14_R2_C113_rom_inst (.q(O14_I14_R2_C1_SM1 ),.address(input_fmap_14[63:56]),.clk(clk),.d(0),.we(0));
//assign O14_I14_R2_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O14_I14_R2_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O14_I14_R2_C113_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O14_I14_R2_C113_rom_inst (.q(O14_I14_R2_C1_SM1 ),.address(input_fmap_14[63:56]),.clock  (clk));
logic [12-1:0] O15_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O15_I15_R0_C06_rom_inst (.q(O15_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I15_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O15_I15_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O15_I15_R0_C06_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O15_I15_R0_C06_rom_inst (.q(O15_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [10-1:0] O15_I15_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_dw_O15_I15_R0_C21_rom_inst (.q(O15_I15_R0_C2_SM1 ),.address(input_fmap_15[23:16]),.clk(clk),.d(0),.we(0));
//assign O15_I15_R0_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O15_I15_R0_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O15_I15_R0_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_dw_O15_I15_R0_C21_rom_inst (.q(O15_I15_R0_C2_SM1 ),.address(input_fmap_15[23:16]),.clock  (clk));
logic [12-1:0] O15_I15_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O15_I15_R1_C05_rom_inst (.q(O15_I15_R1_C0_SM1 ),.address(input_fmap_15[31:24]),.clk(clk),.d(0),.we(0));
//assign O15_I15_R1_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O15_I15_R1_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O15_I15_R1_C05_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O15_I15_R1_C05_rom_inst (.q(O15_I15_R1_C0_SM1 ),.address(input_fmap_15[31:24]),.clock  (clk));
logic [14-1:0] O15_I15_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv5_dw_O15_I15_R1_C126_rom_inst (.q(O15_I15_R1_C1_SM1 ),.address(input_fmap_15[39:32]),.clk(clk),.d(0),.we(0));
//assign O15_I15_R1_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O15_I15_R1_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O15_I15_R1_C126_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv5_dw_O15_I15_R1_C126_rom_inst (.q(O15_I15_R1_C1_SM1 ),.address(input_fmap_15[39:32]),.clock  (clk));
logic [11-1:0] O15_I15_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O15_I15_R1_C23_rom_inst (.q(O15_I15_R1_C2_SM1 ),.address(input_fmap_15[47:40]),.clk(clk),.d(0),.we(0));
//assign O15_I15_R1_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O15_I15_R1_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O15_I15_R1_C23_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O15_I15_R1_C23_rom_inst (.q(O15_I15_R1_C2_SM1 ),.address(input_fmap_15[47:40]),.clock  (clk));
logic [11-1:0] O15_I15_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O15_I15_R2_C03_rom_inst (.q(O15_I15_R2_C0_SM1 ),.address(input_fmap_15[55:48]),.clk(clk),.d(0),.we(0));
//assign O15_I15_R2_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O15_I15_R2_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O15_I15_R2_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O15_I15_R2_C03_rom_inst (.q(O15_I15_R2_C0_SM1 ),.address(input_fmap_15[55:48]),.clock  (clk));
logic [13-1:0] O15_I15_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O15_I15_R2_C110_rom_inst (.q(O15_I15_R2_C1_SM1 ),.address(input_fmap_15[63:56]),.clk(clk),.d(0),.we(0));
//assign O15_I15_R2_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O15_I15_R2_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O15_I15_R2_C110_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O15_I15_R2_C110_rom_inst (.q(O15_I15_R2_C1_SM1 ),.address(input_fmap_15[63:56]),.clock  (clk));
logic [13-1:0] O15_I15_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O15_I15_R2_C28_rom_inst (.q(O15_I15_R2_C2_SM1 ),.address(input_fmap_15[71:64]),.clk(clk),.d(0),.we(0));
//assign O15_I15_R2_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O15_I15_R2_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O15_I15_R2_C28_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O15_I15_R2_C28_rom_inst (.q(O15_I15_R2_C2_SM1 ),.address(input_fmap_15[71:64]),.clock  (clk));
logic [12-1:0] O16_I16_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O16_I16_R0_C06_rom_inst (.q(O16_I16_R0_C0_SM1 ),.address(input_fmap_16[7:0]),.clk(clk),.d(0),.we(0));
//assign O16_I16_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O16_I16_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O16_I16_R0_C06_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O16_I16_R0_C06_rom_inst (.q(O16_I16_R0_C0_SM1 ),.address(input_fmap_16[7:0]),.clock  (clk));
logic [14-1:0] O16_I16_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv5_dw_O16_I16_R0_C121_rom_inst (.q(O16_I16_R0_C1_SM1 ),.address(input_fmap_16[15:8]),.clk(clk),.d(0),.we(0));
//assign O16_I16_R0_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O16_I16_R0_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O16_I16_R0_C121_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv5_dw_O16_I16_R0_C121_rom_inst (.q(O16_I16_R0_C1_SM1 ),.address(input_fmap_16[15:8]),.clock  (clk));
logic [11-1:0] O16_I16_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O16_I16_R0_C22_rom_inst (.q(O16_I16_R0_C2_SM1 ),.address(input_fmap_16[23:16]),.clk(clk),.d(0),.we(0));
//assign O16_I16_R0_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O16_I16_R0_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O16_I16_R0_C22_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O16_I16_R0_C22_rom_inst (.q(O16_I16_R0_C2_SM1 ),.address(input_fmap_16[23:16]),.clock  (clk));
logic [15-1:0] O16_I16_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(15),.INIT_FILE("deepfreeze_rom/deepfreeze_8_15.txt"))
    conv5_dw_O16_I16_R1_C042_rom_inst (.q(O16_I16_R1_C0_SM1 ),.address(input_fmap_16[31:24]),.clk(clk),.d(0),.we(0));
//assign O16_I16_R1_C0_SM1  = 15'h1234;
//always@(posedge clk) begin 
//O16_I16_R1_C0_SM1  <= 15'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O16_I16_R1_C042_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(15))
//    conv5_dw_O16_I16_R1_C042_rom_inst (.q(O16_I16_R1_C0_SM1 ),.address(input_fmap_16[31:24]),.clock  (clk));
logic [12-1:0] O16_I16_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O16_I16_R1_C17_rom_inst (.q(O16_I16_R1_C1_SM1 ),.address(input_fmap_16[39:32]),.clk(clk),.d(0),.we(0));
//assign O16_I16_R1_C1_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O16_I16_R1_C1_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O16_I16_R1_C17_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O16_I16_R1_C17_rom_inst (.q(O16_I16_R1_C1_SM1 ),.address(input_fmap_16[39:32]),.clock  (clk));
logic [12-1:0] O16_I16_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O16_I16_R1_C26_rom_inst (.q(O16_I16_R1_C2_SM1 ),.address(input_fmap_16[47:40]),.clk(clk),.d(0),.we(0));
//assign O16_I16_R1_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O16_I16_R1_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O16_I16_R1_C26_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O16_I16_R1_C26_rom_inst (.q(O16_I16_R1_C2_SM1 ),.address(input_fmap_16[47:40]),.clock  (clk));
logic [14-1:0] O16_I16_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv5_dw_O16_I16_R2_C116_rom_inst (.q(O16_I16_R2_C1_SM1 ),.address(input_fmap_16[63:56]),.clk(clk),.d(0),.we(0));
//assign O16_I16_R2_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O16_I16_R2_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O16_I16_R2_C116_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv5_dw_O16_I16_R2_C116_rom_inst (.q(O16_I16_R2_C1_SM1 ),.address(input_fmap_16[63:56]),.clock  (clk));
logic [11-1:0] O16_I16_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O16_I16_R2_C22_rom_inst (.q(O16_I16_R2_C2_SM1 ),.address(input_fmap_16[71:64]),.clk(clk),.d(0),.we(0));
//assign O16_I16_R2_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O16_I16_R2_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O16_I16_R2_C22_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O16_I16_R2_C22_rom_inst (.q(O16_I16_R2_C2_SM1 ),.address(input_fmap_16[71:64]),.clock  (clk));
logic [12-1:0] O17_I17_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O17_I17_R0_C05_rom_inst (.q(O17_I17_R0_C0_SM1 ),.address(input_fmap_17[7:0]),.clk(clk),.d(0),.we(0));
//assign O17_I17_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O17_I17_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O17_I17_R0_C05_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O17_I17_R0_C05_rom_inst (.q(O17_I17_R0_C0_SM1 ),.address(input_fmap_17[7:0]),.clock  (clk));
logic [13-1:0] O17_I17_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O17_I17_R0_C110_rom_inst (.q(O17_I17_R0_C1_SM1 ),.address(input_fmap_17[15:8]),.clk(clk),.d(0),.we(0));
//assign O17_I17_R0_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O17_I17_R0_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O17_I17_R0_C110_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O17_I17_R0_C110_rom_inst (.q(O17_I17_R0_C1_SM1 ),.address(input_fmap_17[15:8]),.clock  (clk));
logic [11-1:0] O17_I17_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O17_I17_R0_C23_rom_inst (.q(O17_I17_R0_C2_SM1 ),.address(input_fmap_17[23:16]),.clk(clk),.d(0),.we(0));
//assign O17_I17_R0_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O17_I17_R0_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O17_I17_R0_C23_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O17_I17_R0_C23_rom_inst (.q(O17_I17_R0_C2_SM1 ),.address(input_fmap_17[23:16]),.clock  (clk));
logic [13-1:0] O17_I17_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O17_I17_R1_C011_rom_inst (.q(O17_I17_R1_C0_SM1 ),.address(input_fmap_17[31:24]),.clk(clk),.d(0),.we(0));
//assign O17_I17_R1_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O17_I17_R1_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O17_I17_R1_C011_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O17_I17_R1_C011_rom_inst (.q(O17_I17_R1_C0_SM1 ),.address(input_fmap_17[31:24]),.clock  (clk));
logic [15-1:0] O17_I17_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(15),.INIT_FILE("deepfreeze_rom/deepfreeze_8_15.txt"))
    conv5_dw_O17_I17_R1_C135_rom_inst (.q(O17_I17_R1_C1_SM1 ),.address(input_fmap_17[39:32]),.clk(clk),.d(0),.we(0));
//assign O17_I17_R1_C1_SM1  = 15'h1234;
//always@(posedge clk) begin 
//O17_I17_R1_C1_SM1  <= 15'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O17_I17_R1_C135_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(15))
//    conv5_dw_O17_I17_R1_C135_rom_inst (.q(O17_I17_R1_C1_SM1 ),.address(input_fmap_17[39:32]),.clock  (clk));
logic [11-1:0] O17_I17_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O17_I17_R1_C23_rom_inst (.q(O17_I17_R1_C2_SM1 ),.address(input_fmap_17[47:40]),.clk(clk),.d(0),.we(0));
//assign O17_I17_R1_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O17_I17_R1_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O17_I17_R1_C23_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O17_I17_R1_C23_rom_inst (.q(O17_I17_R1_C2_SM1 ),.address(input_fmap_17[47:40]),.clock  (clk));
logic [13-1:0] O17_I17_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O17_I17_R2_C08_rom_inst (.q(O17_I17_R2_C0_SM1 ),.address(input_fmap_17[55:48]),.clk(clk),.d(0),.we(0));
//assign O17_I17_R2_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O17_I17_R2_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O17_I17_R2_C08_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O17_I17_R2_C08_rom_inst (.q(O17_I17_R2_C0_SM1 ),.address(input_fmap_17[55:48]),.clock  (clk));
logic [13-1:0] O17_I17_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O17_I17_R2_C113_rom_inst (.q(O17_I17_R2_C1_SM1 ),.address(input_fmap_17[63:56]),.clk(clk),.d(0),.we(0));
//assign O17_I17_R2_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O17_I17_R2_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O17_I17_R2_C113_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O17_I17_R2_C113_rom_inst (.q(O17_I17_R2_C1_SM1 ),.address(input_fmap_17[63:56]),.clock  (clk));
logic [11-1:0] O17_I17_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O17_I17_R2_C22_rom_inst (.q(O17_I17_R2_C2_SM1 ),.address(input_fmap_17[71:64]),.clk(clk),.d(0),.we(0));
//assign O17_I17_R2_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O17_I17_R2_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O17_I17_R2_C22_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O17_I17_R2_C22_rom_inst (.q(O17_I17_R2_C2_SM1 ),.address(input_fmap_17[71:64]),.clock  (clk));
logic [13-1:0] O18_I18_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O18_I18_R0_C013_rom_inst (.q(O18_I18_R0_C0_SM1 ),.address(input_fmap_18[7:0]),.clk(clk),.d(0),.we(0));
//assign O18_I18_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O18_I18_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O18_I18_R0_C013_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O18_I18_R0_C013_rom_inst (.q(O18_I18_R0_C0_SM1 ),.address(input_fmap_18[7:0]),.clock  (clk));
logic [11-1:0] O18_I18_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O18_I18_R0_C12_rom_inst (.q(O18_I18_R0_C1_SM1 ),.address(input_fmap_18[15:8]),.clk(clk),.d(0),.we(0));
//assign O18_I18_R0_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O18_I18_R0_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O18_I18_R0_C12_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O18_I18_R0_C12_rom_inst (.q(O18_I18_R0_C1_SM1 ),.address(input_fmap_18[15:8]),.clock  (clk));
logic [11-1:0] O18_I18_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O18_I18_R0_C22_rom_inst (.q(O18_I18_R0_C2_SM1 ),.address(input_fmap_18[23:16]),.clk(clk),.d(0),.we(0));
//assign O18_I18_R0_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O18_I18_R0_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O18_I18_R0_C22_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O18_I18_R0_C22_rom_inst (.q(O18_I18_R0_C2_SM1 ),.address(input_fmap_18[23:16]),.clock  (clk));
logic [14-1:0] O18_I18_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv5_dw_O18_I18_R1_C017_rom_inst (.q(O18_I18_R1_C0_SM1 ),.address(input_fmap_18[31:24]),.clk(clk),.d(0),.we(0));
//assign O18_I18_R1_C0_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O18_I18_R1_C0_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O18_I18_R1_C017_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv5_dw_O18_I18_R1_C017_rom_inst (.q(O18_I18_R1_C0_SM1 ),.address(input_fmap_18[31:24]),.clock  (clk));
logic [15-1:0] O18_I18_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(15),.INIT_FILE("deepfreeze_rom/deepfreeze_8_15.txt"))
    conv5_dw_O18_I18_R1_C140_rom_inst (.q(O18_I18_R1_C1_SM1 ),.address(input_fmap_18[39:32]),.clk(clk),.d(0),.we(0));
//assign O18_I18_R1_C1_SM1  = 15'h1234;
//always@(posedge clk) begin 
//O18_I18_R1_C1_SM1  <= 15'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O18_I18_R1_C140_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(15))
//    conv5_dw_O18_I18_R1_C140_rom_inst (.q(O18_I18_R1_C1_SM1 ),.address(input_fmap_18[39:32]),.clock  (clk));
logic [13-1:0] O18_I18_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O18_I18_R1_C29_rom_inst (.q(O18_I18_R1_C2_SM1 ),.address(input_fmap_18[47:40]),.clk(clk),.d(0),.we(0));
//assign O18_I18_R1_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O18_I18_R1_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O18_I18_R1_C29_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O18_I18_R1_C29_rom_inst (.q(O18_I18_R1_C2_SM1 ),.address(input_fmap_18[47:40]),.clock  (clk));
logic [12-1:0] O18_I18_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O18_I18_R2_C05_rom_inst (.q(O18_I18_R2_C0_SM1 ),.address(input_fmap_18[55:48]),.clk(clk),.d(0),.we(0));
//assign O18_I18_R2_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O18_I18_R2_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O18_I18_R2_C05_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O18_I18_R2_C05_rom_inst (.q(O18_I18_R2_C0_SM1 ),.address(input_fmap_18[55:48]),.clock  (clk));
logic [13-1:0] O18_I18_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O18_I18_R2_C111_rom_inst (.q(O18_I18_R2_C1_SM1 ),.address(input_fmap_18[63:56]),.clk(clk),.d(0),.we(0));
//assign O18_I18_R2_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O18_I18_R2_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O18_I18_R2_C111_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O18_I18_R2_C111_rom_inst (.q(O18_I18_R2_C1_SM1 ),.address(input_fmap_18[63:56]),.clock  (clk));
logic [13-1:0] O18_I18_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O18_I18_R2_C210_rom_inst (.q(O18_I18_R2_C2_SM1 ),.address(input_fmap_18[71:64]),.clk(clk),.d(0),.we(0));
//assign O18_I18_R2_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O18_I18_R2_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O18_I18_R2_C210_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O18_I18_R2_C210_rom_inst (.q(O18_I18_R2_C2_SM1 ),.address(input_fmap_18[71:64]),.clock  (clk));
logic [13-1:0] O19_I19_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O19_I19_R0_C09_rom_inst (.q(O19_I19_R0_C0_SM1 ),.address(input_fmap_19[7:0]),.clk(clk),.d(0),.we(0));
//assign O19_I19_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O19_I19_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O19_I19_R0_C09_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O19_I19_R0_C09_rom_inst (.q(O19_I19_R0_C0_SM1 ),.address(input_fmap_19[7:0]),.clock  (clk));
logic [13-1:0] O19_I19_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O19_I19_R0_C113_rom_inst (.q(O19_I19_R0_C1_SM1 ),.address(input_fmap_19[15:8]),.clk(clk),.d(0),.we(0));
//assign O19_I19_R0_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O19_I19_R0_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O19_I19_R0_C113_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O19_I19_R0_C113_rom_inst (.q(O19_I19_R0_C1_SM1 ),.address(input_fmap_19[15:8]),.clock  (clk));
logic [11-1:0] O19_I19_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O19_I19_R0_C22_rom_inst (.q(O19_I19_R0_C2_SM1 ),.address(input_fmap_19[23:16]),.clk(clk),.d(0),.we(0));
//assign O19_I19_R0_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O19_I19_R0_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O19_I19_R0_C22_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O19_I19_R0_C22_rom_inst (.q(O19_I19_R0_C2_SM1 ),.address(input_fmap_19[23:16]),.clock  (clk));
logic [15-1:0] O19_I19_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(15),.INIT_FILE("deepfreeze_rom/deepfreeze_8_15.txt"))
    conv5_dw_O19_I19_R1_C044_rom_inst (.q(O19_I19_R1_C0_SM1 ),.address(input_fmap_19[31:24]),.clk(clk),.d(0),.we(0));
//assign O19_I19_R1_C0_SM1  = 15'h1234;
//always@(posedge clk) begin 
//O19_I19_R1_C0_SM1  <= 15'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O19_I19_R1_C044_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(15))
//    conv5_dw_O19_I19_R1_C044_rom_inst (.q(O19_I19_R1_C0_SM1 ),.address(input_fmap_19[31:24]),.clock  (clk));
logic [12-1:0] O19_I19_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O19_I19_R1_C16_rom_inst (.q(O19_I19_R1_C1_SM1 ),.address(input_fmap_19[39:32]),.clk(clk),.d(0),.we(0));
//assign O19_I19_R1_C1_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O19_I19_R1_C1_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O19_I19_R1_C16_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O19_I19_R1_C16_rom_inst (.q(O19_I19_R1_C1_SM1 ),.address(input_fmap_19[39:32]),.clock  (clk));
logic [12-1:0] O19_I19_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O19_I19_R1_C24_rom_inst (.q(O19_I19_R1_C2_SM1 ),.address(input_fmap_19[47:40]),.clk(clk),.d(0),.we(0));
//assign O19_I19_R1_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O19_I19_R1_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O19_I19_R1_C24_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O19_I19_R1_C24_rom_inst (.q(O19_I19_R1_C2_SM1 ),.address(input_fmap_19[47:40]),.clock  (clk));
logic [13-1:0] O19_I19_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O19_I19_R2_C09_rom_inst (.q(O19_I19_R2_C0_SM1 ),.address(input_fmap_19[55:48]),.clk(clk),.d(0),.we(0));
//assign O19_I19_R2_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O19_I19_R2_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O19_I19_R2_C09_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O19_I19_R2_C09_rom_inst (.q(O19_I19_R2_C0_SM1 ),.address(input_fmap_19[55:48]),.clock  (clk));
logic [13-1:0] O19_I19_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O19_I19_R2_C114_rom_inst (.q(O19_I19_R2_C1_SM1 ),.address(input_fmap_19[63:56]),.clk(clk),.d(0),.we(0));
//assign O19_I19_R2_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O19_I19_R2_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O19_I19_R2_C114_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O19_I19_R2_C114_rom_inst (.q(O19_I19_R2_C1_SM1 ),.address(input_fmap_19[63:56]),.clock  (clk));
logic [11-1:0] O19_I19_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O19_I19_R2_C23_rom_inst (.q(O19_I19_R2_C2_SM1 ),.address(input_fmap_19[71:64]),.clk(clk),.d(0),.we(0));
//assign O19_I19_R2_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O19_I19_R2_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O19_I19_R2_C23_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O19_I19_R2_C23_rom_inst (.q(O19_I19_R2_C2_SM1 ),.address(input_fmap_19[71:64]),.clock  (clk));
logic [11-1:0] O20_I20_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O20_I20_R0_C02_rom_inst (.q(O20_I20_R0_C0_SM1 ),.address(input_fmap_20[7:0]),.clk(clk),.d(0),.we(0));
//assign O20_I20_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O20_I20_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O20_I20_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O20_I20_R0_C02_rom_inst (.q(O20_I20_R0_C0_SM1 ),.address(input_fmap_20[7:0]),.clock  (clk));
logic [11-1:0] O20_I20_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O20_I20_R0_C12_rom_inst (.q(O20_I20_R0_C1_SM1 ),.address(input_fmap_20[15:8]),.clk(clk),.d(0),.we(0));
//assign O20_I20_R0_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O20_I20_R0_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O20_I20_R0_C12_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O20_I20_R0_C12_rom_inst (.q(O20_I20_R0_C1_SM1 ),.address(input_fmap_20[15:8]),.clock  (clk));
logic [12-1:0] O20_I20_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O20_I20_R0_C24_rom_inst (.q(O20_I20_R0_C2_SM1 ),.address(input_fmap_20[23:16]),.clk(clk),.d(0),.we(0));
//assign O20_I20_R0_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O20_I20_R0_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O20_I20_R0_C24_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O20_I20_R0_C24_rom_inst (.q(O20_I20_R0_C2_SM1 ),.address(input_fmap_20[23:16]),.clock  (clk));
logic [15-1:0] O20_I20_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(15),.INIT_FILE("deepfreeze_rom/deepfreeze_8_15.txt"))
    conv5_dw_O20_I20_R1_C034_rom_inst (.q(O20_I20_R1_C0_SM1 ),.address(input_fmap_20[31:24]),.clk(clk),.d(0),.we(0));
//assign O20_I20_R1_C0_SM1  = 15'h1234;
//always@(posedge clk) begin 
//O20_I20_R1_C0_SM1  <= 15'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O20_I20_R1_C034_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(15))
//    conv5_dw_O20_I20_R1_C034_rom_inst (.q(O20_I20_R1_C0_SM1 ),.address(input_fmap_20[31:24]),.clock  (clk));
logic [14-1:0] O20_I20_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv5_dw_O20_I20_R1_C126_rom_inst (.q(O20_I20_R1_C1_SM1 ),.address(input_fmap_20[39:32]),.clk(clk),.d(0),.we(0));
//assign O20_I20_R1_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O20_I20_R1_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O20_I20_R1_C126_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv5_dw_O20_I20_R1_C126_rom_inst (.q(O20_I20_R1_C1_SM1 ),.address(input_fmap_20[39:32]),.clock  (clk));
logic [11-1:0] O20_I20_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O20_I20_R1_C22_rom_inst (.q(O20_I20_R1_C2_SM1 ),.address(input_fmap_20[47:40]),.clk(clk),.d(0),.we(0));
//assign O20_I20_R1_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O20_I20_R1_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O20_I20_R1_C22_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O20_I20_R1_C22_rom_inst (.q(O20_I20_R1_C2_SM1 ),.address(input_fmap_20[47:40]),.clock  (clk));
logic [12-1:0] O20_I20_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O20_I20_R2_C06_rom_inst (.q(O20_I20_R2_C0_SM1 ),.address(input_fmap_20[55:48]),.clk(clk),.d(0),.we(0));
//assign O20_I20_R2_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O20_I20_R2_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O20_I20_R2_C06_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O20_I20_R2_C06_rom_inst (.q(O20_I20_R2_C0_SM1 ),.address(input_fmap_20[55:48]),.clock  (clk));
logic [10-1:0] O20_I20_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_dw_O20_I20_R2_C11_rom_inst (.q(O20_I20_R2_C1_SM1 ),.address(input_fmap_20[63:56]),.clk(clk),.d(0),.we(0));
//assign O20_I20_R2_C1_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O20_I20_R2_C1_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O20_I20_R2_C11_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_dw_O20_I20_R2_C11_rom_inst (.q(O20_I20_R2_C1_SM1 ),.address(input_fmap_20[63:56]),.clock  (clk));
logic [11-1:0] O20_I20_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O20_I20_R2_C23_rom_inst (.q(O20_I20_R2_C2_SM1 ),.address(input_fmap_20[71:64]),.clk(clk),.d(0),.we(0));
//assign O20_I20_R2_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O20_I20_R2_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O20_I20_R2_C23_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O20_I20_R2_C23_rom_inst (.q(O20_I20_R2_C2_SM1 ),.address(input_fmap_20[71:64]),.clock  (clk));
logic [11-1:0] O21_I21_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O21_I21_R0_C02_rom_inst (.q(O21_I21_R0_C0_SM1 ),.address(input_fmap_21[7:0]),.clk(clk),.d(0),.we(0));
//assign O21_I21_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O21_I21_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O21_I21_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O21_I21_R0_C02_rom_inst (.q(O21_I21_R0_C0_SM1 ),.address(input_fmap_21[7:0]),.clock  (clk));
logic [12-1:0] O21_I21_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O21_I21_R0_C15_rom_inst (.q(O21_I21_R0_C1_SM1 ),.address(input_fmap_21[15:8]),.clk(clk),.d(0),.we(0));
//assign O21_I21_R0_C1_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O21_I21_R0_C1_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O21_I21_R0_C15_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O21_I21_R0_C15_rom_inst (.q(O21_I21_R0_C1_SM1 ),.address(input_fmap_21[15:8]),.clock  (clk));
logic [13-1:0] O21_I21_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O21_I21_R0_C29_rom_inst (.q(O21_I21_R0_C2_SM1 ),.address(input_fmap_21[23:16]),.clk(clk),.d(0),.we(0));
//assign O21_I21_R0_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O21_I21_R0_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O21_I21_R0_C29_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O21_I21_R0_C29_rom_inst (.q(O21_I21_R0_C2_SM1 ),.address(input_fmap_21[23:16]),.clock  (clk));
logic [13-1:0] O21_I21_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O21_I21_R1_C014_rom_inst (.q(O21_I21_R1_C0_SM1 ),.address(input_fmap_21[31:24]),.clk(clk),.d(0),.we(0));
//assign O21_I21_R1_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O21_I21_R1_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O21_I21_R1_C014_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O21_I21_R1_C014_rom_inst (.q(O21_I21_R1_C0_SM1 ),.address(input_fmap_21[31:24]),.clock  (clk));
logic [14-1:0] O21_I21_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv5_dw_O21_I21_R1_C117_rom_inst (.q(O21_I21_R1_C1_SM1 ),.address(input_fmap_21[39:32]),.clk(clk),.d(0),.we(0));
//assign O21_I21_R1_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O21_I21_R1_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O21_I21_R1_C117_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv5_dw_O21_I21_R1_C117_rom_inst (.q(O21_I21_R1_C1_SM1 ),.address(input_fmap_21[39:32]),.clock  (clk));
logic [10-1:0] O21_I21_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_dw_O21_I21_R1_C21_rom_inst (.q(O21_I21_R1_C2_SM1 ),.address(input_fmap_21[47:40]),.clk(clk),.d(0),.we(0));
//assign O21_I21_R1_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O21_I21_R1_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O21_I21_R1_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_dw_O21_I21_R1_C21_rom_inst (.q(O21_I21_R1_C2_SM1 ),.address(input_fmap_21[47:40]),.clock  (clk));
logic [13-1:0] O21_I21_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O21_I21_R2_C010_rom_inst (.q(O21_I21_R2_C0_SM1 ),.address(input_fmap_21[55:48]),.clk(clk),.d(0),.we(0));
//assign O21_I21_R2_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O21_I21_R2_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O21_I21_R2_C010_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O21_I21_R2_C010_rom_inst (.q(O21_I21_R2_C0_SM1 ),.address(input_fmap_21[55:48]),.clock  (clk));
logic [12-1:0] O21_I21_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O21_I21_R2_C15_rom_inst (.q(O21_I21_R2_C1_SM1 ),.address(input_fmap_21[63:56]),.clk(clk),.d(0),.we(0));
//assign O21_I21_R2_C1_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O21_I21_R2_C1_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O21_I21_R2_C15_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O21_I21_R2_C15_rom_inst (.q(O21_I21_R2_C1_SM1 ),.address(input_fmap_21[63:56]),.clock  (clk));
logic [13-1:0] O21_I21_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O21_I21_R2_C28_rom_inst (.q(O21_I21_R2_C2_SM1 ),.address(input_fmap_21[71:64]),.clk(clk),.d(0),.we(0));
//assign O21_I21_R2_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O21_I21_R2_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O21_I21_R2_C28_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O21_I21_R2_C28_rom_inst (.q(O21_I21_R2_C2_SM1 ),.address(input_fmap_21[71:64]),.clock  (clk));
logic [12-1:0] O22_I22_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O22_I22_R0_C05_rom_inst (.q(O22_I22_R0_C0_SM1 ),.address(input_fmap_22[7:0]),.clk(clk),.d(0),.we(0));
//assign O22_I22_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O22_I22_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O22_I22_R0_C05_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O22_I22_R0_C05_rom_inst (.q(O22_I22_R0_C0_SM1 ),.address(input_fmap_22[7:0]),.clock  (clk));
logic [11-1:0] O22_I22_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O22_I22_R0_C13_rom_inst (.q(O22_I22_R0_C1_SM1 ),.address(input_fmap_22[15:8]),.clk(clk),.d(0),.we(0));
//assign O22_I22_R0_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O22_I22_R0_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O22_I22_R0_C13_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O22_I22_R0_C13_rom_inst (.q(O22_I22_R0_C1_SM1 ),.address(input_fmap_22[15:8]),.clock  (clk));
logic [11-1:0] O22_I22_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O22_I22_R0_C22_rom_inst (.q(O22_I22_R0_C2_SM1 ),.address(input_fmap_22[23:16]),.clk(clk),.d(0),.we(0));
//assign O22_I22_R0_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O22_I22_R0_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O22_I22_R0_C22_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O22_I22_R0_C22_rom_inst (.q(O22_I22_R0_C2_SM1 ),.address(input_fmap_22[23:16]),.clock  (clk));
logic [13-1:0] O22_I22_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O22_I22_R1_C09_rom_inst (.q(O22_I22_R1_C0_SM1 ),.address(input_fmap_22[31:24]),.clk(clk),.d(0),.we(0));
//assign O22_I22_R1_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O22_I22_R1_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O22_I22_R1_C09_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O22_I22_R1_C09_rom_inst (.q(O22_I22_R1_C0_SM1 ),.address(input_fmap_22[31:24]),.clock  (clk));
logic [14-1:0] O22_I22_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv5_dw_O22_I22_R1_C130_rom_inst (.q(O22_I22_R1_C1_SM1 ),.address(input_fmap_22[39:32]),.clk(clk),.d(0),.we(0));
//assign O22_I22_R1_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O22_I22_R1_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O22_I22_R1_C130_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv5_dw_O22_I22_R1_C130_rom_inst (.q(O22_I22_R1_C1_SM1 ),.address(input_fmap_22[39:32]),.clock  (clk));
logic [13-1:0] O22_I22_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O22_I22_R1_C29_rom_inst (.q(O22_I22_R1_C2_SM1 ),.address(input_fmap_22[47:40]),.clk(clk),.d(0),.we(0));
//assign O22_I22_R1_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O22_I22_R1_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O22_I22_R1_C29_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O22_I22_R1_C29_rom_inst (.q(O22_I22_R1_C2_SM1 ),.address(input_fmap_22[47:40]),.clock  (clk));
logic [10-1:0] O22_I22_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_dw_O22_I22_R2_C01_rom_inst (.q(O22_I22_R2_C0_SM1 ),.address(input_fmap_22[55:48]),.clk(clk),.d(0),.we(0));
//assign O22_I22_R2_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O22_I22_R2_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O22_I22_R2_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_dw_O22_I22_R2_C01_rom_inst (.q(O22_I22_R2_C0_SM1 ),.address(input_fmap_22[55:48]),.clock  (clk));
logic [12-1:0] O22_I22_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O22_I22_R2_C15_rom_inst (.q(O22_I22_R2_C1_SM1 ),.address(input_fmap_22[63:56]),.clk(clk),.d(0),.we(0));
//assign O22_I22_R2_C1_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O22_I22_R2_C1_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O22_I22_R2_C15_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O22_I22_R2_C15_rom_inst (.q(O22_I22_R2_C1_SM1 ),.address(input_fmap_22[63:56]),.clock  (clk));
logic [11-1:0] O22_I22_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O22_I22_R2_C22_rom_inst (.q(O22_I22_R2_C2_SM1 ),.address(input_fmap_22[71:64]),.clk(clk),.d(0),.we(0));
//assign O22_I22_R2_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O22_I22_R2_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O22_I22_R2_C22_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O22_I22_R2_C22_rom_inst (.q(O22_I22_R2_C2_SM1 ),.address(input_fmap_22[71:64]),.clock  (clk));
logic [13-1:0] O23_I23_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O23_I23_R0_C012_rom_inst (.q(O23_I23_R0_C0_SM1 ),.address(input_fmap_23[7:0]),.clk(clk),.d(0),.we(0));
//assign O23_I23_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O23_I23_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O23_I23_R0_C012_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O23_I23_R0_C012_rom_inst (.q(O23_I23_R0_C0_SM1 ),.address(input_fmap_23[7:0]),.clock  (clk));
logic [13-1:0] O23_I23_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O23_I23_R0_C115_rom_inst (.q(O23_I23_R0_C1_SM1 ),.address(input_fmap_23[15:8]),.clk(clk),.d(0),.we(0));
//assign O23_I23_R0_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O23_I23_R0_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O23_I23_R0_C115_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O23_I23_R0_C115_rom_inst (.q(O23_I23_R0_C1_SM1 ),.address(input_fmap_23[15:8]),.clock  (clk));
logic [11-1:0] O23_I23_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O23_I23_R0_C22_rom_inst (.q(O23_I23_R0_C2_SM1 ),.address(input_fmap_23[23:16]),.clk(clk),.d(0),.we(0));
//assign O23_I23_R0_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O23_I23_R0_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O23_I23_R0_C22_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O23_I23_R0_C22_rom_inst (.q(O23_I23_R0_C2_SM1 ),.address(input_fmap_23[23:16]),.clock  (clk));
logic [13-1:0] O23_I23_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O23_I23_R1_C014_rom_inst (.q(O23_I23_R1_C0_SM1 ),.address(input_fmap_23[31:24]),.clk(clk),.d(0),.we(0));
//assign O23_I23_R1_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O23_I23_R1_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O23_I23_R1_C014_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O23_I23_R1_C014_rom_inst (.q(O23_I23_R1_C0_SM1 ),.address(input_fmap_23[31:24]),.clock  (clk));
logic [12-1:0] O23_I23_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O23_I23_R1_C16_rom_inst (.q(O23_I23_R1_C1_SM1 ),.address(input_fmap_23[39:32]),.clk(clk),.d(0),.we(0));
//assign O23_I23_R1_C1_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O23_I23_R1_C1_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O23_I23_R1_C16_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O23_I23_R1_C16_rom_inst (.q(O23_I23_R1_C1_SM1 ),.address(input_fmap_23[39:32]),.clock  (clk));
logic [12-1:0] O23_I23_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O23_I23_R1_C24_rom_inst (.q(O23_I23_R1_C2_SM1 ),.address(input_fmap_23[47:40]),.clk(clk),.d(0),.we(0));
//assign O23_I23_R1_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O23_I23_R1_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O23_I23_R1_C24_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O23_I23_R1_C24_rom_inst (.q(O23_I23_R1_C2_SM1 ),.address(input_fmap_23[47:40]),.clock  (clk));
logic [11-1:0] O23_I23_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O23_I23_R2_C02_rom_inst (.q(O23_I23_R2_C0_SM1 ),.address(input_fmap_23[55:48]),.clk(clk),.d(0),.we(0));
//assign O23_I23_R2_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O23_I23_R2_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O23_I23_R2_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O23_I23_R2_C02_rom_inst (.q(O23_I23_R2_C0_SM1 ),.address(input_fmap_23[55:48]),.clock  (clk));
logic [11-1:0] O23_I23_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O23_I23_R2_C12_rom_inst (.q(O23_I23_R2_C1_SM1 ),.address(input_fmap_23[63:56]),.clk(clk),.d(0),.we(0));
//assign O23_I23_R2_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O23_I23_R2_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O23_I23_R2_C12_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O23_I23_R2_C12_rom_inst (.q(O23_I23_R2_C1_SM1 ),.address(input_fmap_23[63:56]),.clock  (clk));
logic [11-1:0] O23_I23_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O23_I23_R2_C23_rom_inst (.q(O23_I23_R2_C2_SM1 ),.address(input_fmap_23[71:64]),.clk(clk),.d(0),.we(0));
//assign O23_I23_R2_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O23_I23_R2_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O23_I23_R2_C23_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O23_I23_R2_C23_rom_inst (.q(O23_I23_R2_C2_SM1 ),.address(input_fmap_23[71:64]),.clock  (clk));
logic [13-1:0] O24_I24_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O24_I24_R0_C010_rom_inst (.q(O24_I24_R0_C0_SM1 ),.address(input_fmap_24[7:0]),.clk(clk),.d(0),.we(0));
//assign O24_I24_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O24_I24_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O24_I24_R0_C010_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O24_I24_R0_C010_rom_inst (.q(O24_I24_R0_C0_SM1 ),.address(input_fmap_24[7:0]),.clock  (clk));
logic [13-1:0] O24_I24_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O24_I24_R0_C19_rom_inst (.q(O24_I24_R0_C1_SM1 ),.address(input_fmap_24[15:8]),.clk(clk),.d(0),.we(0));
//assign O24_I24_R0_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O24_I24_R0_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O24_I24_R0_C19_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O24_I24_R0_C19_rom_inst (.q(O24_I24_R0_C1_SM1 ),.address(input_fmap_24[15:8]),.clock  (clk));
logic [11-1:0] O24_I24_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O24_I24_R0_C22_rom_inst (.q(O24_I24_R0_C2_SM1 ),.address(input_fmap_24[23:16]),.clk(clk),.d(0),.we(0));
//assign O24_I24_R0_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O24_I24_R0_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O24_I24_R0_C22_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O24_I24_R0_C22_rom_inst (.q(O24_I24_R0_C2_SM1 ),.address(input_fmap_24[23:16]),.clock  (clk));
logic [12-1:0] O24_I24_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O24_I24_R1_C07_rom_inst (.q(O24_I24_R1_C0_SM1 ),.address(input_fmap_24[31:24]),.clk(clk),.d(0),.we(0));
//assign O24_I24_R1_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O24_I24_R1_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O24_I24_R1_C07_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O24_I24_R1_C07_rom_inst (.q(O24_I24_R1_C0_SM1 ),.address(input_fmap_24[31:24]),.clock  (clk));
logic [13-1:0] O24_I24_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O24_I24_R1_C18_rom_inst (.q(O24_I24_R1_C1_SM1 ),.address(input_fmap_24[39:32]),.clk(clk),.d(0),.we(0));
//assign O24_I24_R1_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O24_I24_R1_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O24_I24_R1_C18_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O24_I24_R1_C18_rom_inst (.q(O24_I24_R1_C1_SM1 ),.address(input_fmap_24[39:32]),.clock  (clk));
logic [13-1:0] O24_I24_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O24_I24_R1_C211_rom_inst (.q(O24_I24_R1_C2_SM1 ),.address(input_fmap_24[47:40]),.clk(clk),.d(0),.we(0));
//assign O24_I24_R1_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O24_I24_R1_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O24_I24_R1_C211_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O24_I24_R1_C211_rom_inst (.q(O24_I24_R1_C2_SM1 ),.address(input_fmap_24[47:40]),.clock  (clk));
logic [11-1:0] O24_I24_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O24_I24_R2_C02_rom_inst (.q(O24_I24_R2_C0_SM1 ),.address(input_fmap_24[55:48]),.clk(clk),.d(0),.we(0));
//assign O24_I24_R2_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O24_I24_R2_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O24_I24_R2_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O24_I24_R2_C02_rom_inst (.q(O24_I24_R2_C0_SM1 ),.address(input_fmap_24[55:48]),.clock  (clk));
logic [11-1:0] O24_I24_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O24_I24_R2_C13_rom_inst (.q(O24_I24_R2_C1_SM1 ),.address(input_fmap_24[63:56]),.clk(clk),.d(0),.we(0));
//assign O24_I24_R2_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O24_I24_R2_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O24_I24_R2_C13_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O24_I24_R2_C13_rom_inst (.q(O24_I24_R2_C1_SM1 ),.address(input_fmap_24[63:56]),.clock  (clk));
logic [13-1:0] O25_I25_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O25_I25_R0_C08_rom_inst (.q(O25_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clk(clk),.d(0),.we(0));
//assign O25_I25_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O25_I25_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O25_I25_R0_C08_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O25_I25_R0_C08_rom_inst (.q(O25_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clock  (clk));
logic [13-1:0] O25_I25_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O25_I25_R0_C110_rom_inst (.q(O25_I25_R0_C1_SM1 ),.address(input_fmap_25[15:8]),.clk(clk),.d(0),.we(0));
//assign O25_I25_R0_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O25_I25_R0_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O25_I25_R0_C110_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O25_I25_R0_C110_rom_inst (.q(O25_I25_R0_C1_SM1 ),.address(input_fmap_25[15:8]),.clock  (clk));
logic [12-1:0] O25_I25_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O25_I25_R0_C27_rom_inst (.q(O25_I25_R0_C2_SM1 ),.address(input_fmap_25[23:16]),.clk(clk),.d(0),.we(0));
//assign O25_I25_R0_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O25_I25_R0_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O25_I25_R0_C27_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O25_I25_R0_C27_rom_inst (.q(O25_I25_R0_C2_SM1 ),.address(input_fmap_25[23:16]),.clock  (clk));
logic [14-1:0] O25_I25_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv5_dw_O25_I25_R1_C026_rom_inst (.q(O25_I25_R1_C0_SM1 ),.address(input_fmap_25[31:24]),.clk(clk),.d(0),.we(0));
//assign O25_I25_R1_C0_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O25_I25_R1_C0_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O25_I25_R1_C026_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv5_dw_O25_I25_R1_C026_rom_inst (.q(O25_I25_R1_C0_SM1 ),.address(input_fmap_25[31:24]),.clock  (clk));
logic [15-1:0] O25_I25_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(15),.INIT_FILE("deepfreeze_rom/deepfreeze_8_15.txt"))
    conv5_dw_O25_I25_R1_C142_rom_inst (.q(O25_I25_R1_C1_SM1 ),.address(input_fmap_25[39:32]),.clk(clk),.d(0),.we(0));
//assign O25_I25_R1_C1_SM1  = 15'h1234;
//always@(posedge clk) begin 
//O25_I25_R1_C1_SM1  <= 15'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O25_I25_R1_C142_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(15))
//    conv5_dw_O25_I25_R1_C142_rom_inst (.q(O25_I25_R1_C1_SM1 ),.address(input_fmap_25[39:32]),.clock  (clk));
logic [13-1:0] O25_I25_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O25_I25_R1_C214_rom_inst (.q(O25_I25_R1_C2_SM1 ),.address(input_fmap_25[47:40]),.clk(clk),.d(0),.we(0));
//assign O25_I25_R1_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O25_I25_R1_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O25_I25_R1_C214_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O25_I25_R1_C214_rom_inst (.q(O25_I25_R1_C2_SM1 ),.address(input_fmap_25[47:40]),.clock  (clk));
logic [14-1:0] O25_I25_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv5_dw_O25_I25_R2_C019_rom_inst (.q(O25_I25_R2_C0_SM1 ),.address(input_fmap_25[55:48]),.clk(clk),.d(0),.we(0));
//assign O25_I25_R2_C0_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O25_I25_R2_C0_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O25_I25_R2_C019_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv5_dw_O25_I25_R2_C019_rom_inst (.q(O25_I25_R2_C0_SM1 ),.address(input_fmap_25[55:48]),.clock  (clk));
logic [11-1:0] O25_I25_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O25_I25_R2_C12_rom_inst (.q(O25_I25_R2_C1_SM1 ),.address(input_fmap_25[63:56]),.clk(clk),.d(0),.we(0));
//assign O25_I25_R2_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O25_I25_R2_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O25_I25_R2_C12_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O25_I25_R2_C12_rom_inst (.q(O25_I25_R2_C1_SM1 ),.address(input_fmap_25[63:56]),.clock  (clk));
logic [12-1:0] O25_I25_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O25_I25_R2_C24_rom_inst (.q(O25_I25_R2_C2_SM1 ),.address(input_fmap_25[71:64]),.clk(clk),.d(0),.we(0));
//assign O25_I25_R2_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O25_I25_R2_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O25_I25_R2_C24_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O25_I25_R2_C24_rom_inst (.q(O25_I25_R2_C2_SM1 ),.address(input_fmap_25[71:64]),.clock  (clk));
logic [10-1:0] O26_I26_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_dw_O26_I26_R0_C01_rom_inst (.q(O26_I26_R0_C0_SM1 ),.address(input_fmap_26[7:0]),.clk(clk),.d(0),.we(0));
//assign O26_I26_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O26_I26_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O26_I26_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_dw_O26_I26_R0_C01_rom_inst (.q(O26_I26_R0_C0_SM1 ),.address(input_fmap_26[7:0]),.clock  (clk));
logic [13-1:0] O26_I26_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O26_I26_R0_C18_rom_inst (.q(O26_I26_R0_C1_SM1 ),.address(input_fmap_26[15:8]),.clk(clk),.d(0),.we(0));
//assign O26_I26_R0_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O26_I26_R0_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O26_I26_R0_C18_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O26_I26_R0_C18_rom_inst (.q(O26_I26_R0_C1_SM1 ),.address(input_fmap_26[15:8]),.clock  (clk));
logic [11-1:0] O26_I26_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O26_I26_R0_C22_rom_inst (.q(O26_I26_R0_C2_SM1 ),.address(input_fmap_26[23:16]),.clk(clk),.d(0),.we(0));
//assign O26_I26_R0_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O26_I26_R0_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O26_I26_R0_C22_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O26_I26_R0_C22_rom_inst (.q(O26_I26_R0_C2_SM1 ),.address(input_fmap_26[23:16]),.clock  (clk));
logic [13-1:0] O26_I26_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O26_I26_R1_C013_rom_inst (.q(O26_I26_R1_C0_SM1 ),.address(input_fmap_26[31:24]),.clk(clk),.d(0),.we(0));
//assign O26_I26_R1_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O26_I26_R1_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O26_I26_R1_C013_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O26_I26_R1_C013_rom_inst (.q(O26_I26_R1_C0_SM1 ),.address(input_fmap_26[31:24]),.clock  (clk));
logic [14-1:0] O26_I26_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv5_dw_O26_I26_R1_C123_rom_inst (.q(O26_I26_R1_C1_SM1 ),.address(input_fmap_26[39:32]),.clk(clk),.d(0),.we(0));
//assign O26_I26_R1_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O26_I26_R1_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O26_I26_R1_C123_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv5_dw_O26_I26_R1_C123_rom_inst (.q(O26_I26_R1_C1_SM1 ),.address(input_fmap_26[39:32]),.clock  (clk));
logic [13-1:0] O26_I26_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O26_I26_R1_C210_rom_inst (.q(O26_I26_R1_C2_SM1 ),.address(input_fmap_26[47:40]),.clk(clk),.d(0),.we(0));
//assign O26_I26_R1_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O26_I26_R1_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O26_I26_R1_C210_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O26_I26_R1_C210_rom_inst (.q(O26_I26_R1_C2_SM1 ),.address(input_fmap_26[47:40]),.clock  (clk));
logic [12-1:0] O26_I26_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O26_I26_R2_C04_rom_inst (.q(O26_I26_R2_C0_SM1 ),.address(input_fmap_26[55:48]),.clk(clk),.d(0),.we(0));
//assign O26_I26_R2_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O26_I26_R2_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O26_I26_R2_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O26_I26_R2_C04_rom_inst (.q(O26_I26_R2_C0_SM1 ),.address(input_fmap_26[55:48]),.clock  (clk));
logic [12-1:0] O26_I26_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O26_I26_R2_C17_rom_inst (.q(O26_I26_R2_C1_SM1 ),.address(input_fmap_26[63:56]),.clk(clk),.d(0),.we(0));
//assign O26_I26_R2_C1_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O26_I26_R2_C1_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O26_I26_R2_C17_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O26_I26_R2_C17_rom_inst (.q(O26_I26_R2_C1_SM1 ),.address(input_fmap_26[63:56]),.clock  (clk));
logic [10-1:0] O26_I26_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_dw_O26_I26_R2_C21_rom_inst (.q(O26_I26_R2_C2_SM1 ),.address(input_fmap_26[71:64]),.clk(clk),.d(0),.we(0));
//assign O26_I26_R2_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O26_I26_R2_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O26_I26_R2_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_dw_O26_I26_R2_C21_rom_inst (.q(O26_I26_R2_C2_SM1 ),.address(input_fmap_26[71:64]),.clock  (clk));
logic [10-1:0] O27_I27_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_dw_O27_I27_R0_C01_rom_inst (.q(O27_I27_R0_C0_SM1 ),.address(input_fmap_27[7:0]),.clk(clk),.d(0),.we(0));
//assign O27_I27_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O27_I27_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O27_I27_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_dw_O27_I27_R0_C01_rom_inst (.q(O27_I27_R0_C0_SM1 ),.address(input_fmap_27[7:0]),.clock  (clk));
logic [12-1:0] O27_I27_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O27_I27_R0_C17_rom_inst (.q(O27_I27_R0_C1_SM1 ),.address(input_fmap_27[15:8]),.clk(clk),.d(0),.we(0));
//assign O27_I27_R0_C1_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O27_I27_R0_C1_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O27_I27_R0_C17_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O27_I27_R0_C17_rom_inst (.q(O27_I27_R0_C1_SM1 ),.address(input_fmap_27[15:8]),.clock  (clk));
logic [11-1:0] O27_I27_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O27_I27_R0_C23_rom_inst (.q(O27_I27_R0_C2_SM1 ),.address(input_fmap_27[23:16]),.clk(clk),.d(0),.we(0));
//assign O27_I27_R0_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O27_I27_R0_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O27_I27_R0_C23_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O27_I27_R0_C23_rom_inst (.q(O27_I27_R0_C2_SM1 ),.address(input_fmap_27[23:16]),.clock  (clk));
logic [14-1:0] O27_I27_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv5_dw_O27_I27_R1_C017_rom_inst (.q(O27_I27_R1_C0_SM1 ),.address(input_fmap_27[31:24]),.clk(clk),.d(0),.we(0));
//assign O27_I27_R1_C0_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O27_I27_R1_C0_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O27_I27_R1_C017_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv5_dw_O27_I27_R1_C017_rom_inst (.q(O27_I27_R1_C0_SM1 ),.address(input_fmap_27[31:24]),.clock  (clk));
logic [14-1:0] O27_I27_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv5_dw_O27_I27_R1_C131_rom_inst (.q(O27_I27_R1_C1_SM1 ),.address(input_fmap_27[39:32]),.clk(clk),.d(0),.we(0));
//assign O27_I27_R1_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O27_I27_R1_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O27_I27_R1_C131_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv5_dw_O27_I27_R1_C131_rom_inst (.q(O27_I27_R1_C1_SM1 ),.address(input_fmap_27[39:32]),.clock  (clk));
logic [13-1:0] O27_I27_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O27_I27_R1_C214_rom_inst (.q(O27_I27_R1_C2_SM1 ),.address(input_fmap_27[47:40]),.clk(clk),.d(0),.we(0));
//assign O27_I27_R1_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O27_I27_R1_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O27_I27_R1_C214_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O27_I27_R1_C214_rom_inst (.q(O27_I27_R1_C2_SM1 ),.address(input_fmap_27[47:40]),.clock  (clk));
logic [13-1:0] O27_I27_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O27_I27_R2_C012_rom_inst (.q(O27_I27_R2_C0_SM1 ),.address(input_fmap_27[55:48]),.clk(clk),.d(0),.we(0));
//assign O27_I27_R2_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O27_I27_R2_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O27_I27_R2_C012_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O27_I27_R2_C012_rom_inst (.q(O27_I27_R2_C0_SM1 ),.address(input_fmap_27[55:48]),.clock  (clk));
logic [13-1:0] O27_I27_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O27_I27_R2_C113_rom_inst (.q(O27_I27_R2_C1_SM1 ),.address(input_fmap_27[63:56]),.clk(clk),.d(0),.we(0));
//assign O27_I27_R2_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O27_I27_R2_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O27_I27_R2_C113_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O27_I27_R2_C113_rom_inst (.q(O27_I27_R2_C1_SM1 ),.address(input_fmap_27[63:56]),.clock  (clk));
logic [12-1:0] O27_I27_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O27_I27_R2_C25_rom_inst (.q(O27_I27_R2_C2_SM1 ),.address(input_fmap_27[71:64]),.clk(clk),.d(0),.we(0));
//assign O27_I27_R2_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O27_I27_R2_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O27_I27_R2_C25_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O27_I27_R2_C25_rom_inst (.q(O27_I27_R2_C2_SM1 ),.address(input_fmap_27[71:64]),.clock  (clk));
logic [10-1:0] O28_I28_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_dw_O28_I28_R0_C01_rom_inst (.q(O28_I28_R0_C0_SM1 ),.address(input_fmap_28[7:0]),.clk(clk),.d(0),.we(0));
//assign O28_I28_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O28_I28_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O28_I28_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_dw_O28_I28_R0_C01_rom_inst (.q(O28_I28_R0_C0_SM1 ),.address(input_fmap_28[7:0]),.clock  (clk));
logic [13-1:0] O28_I28_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O28_I28_R0_C112_rom_inst (.q(O28_I28_R0_C1_SM1 ),.address(input_fmap_28[15:8]),.clk(clk),.d(0),.we(0));
//assign O28_I28_R0_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O28_I28_R0_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O28_I28_R0_C112_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O28_I28_R0_C112_rom_inst (.q(O28_I28_R0_C1_SM1 ),.address(input_fmap_28[15:8]),.clock  (clk));
logic [13-1:0] O28_I28_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O28_I28_R1_C09_rom_inst (.q(O28_I28_R1_C0_SM1 ),.address(input_fmap_28[31:24]),.clk(clk),.d(0),.we(0));
//assign O28_I28_R1_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O28_I28_R1_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O28_I28_R1_C09_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O28_I28_R1_C09_rom_inst (.q(O28_I28_R1_C0_SM1 ),.address(input_fmap_28[31:24]),.clock  (clk));
logic [13-1:0] O28_I28_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O28_I28_R1_C110_rom_inst (.q(O28_I28_R1_C1_SM1 ),.address(input_fmap_28[39:32]),.clk(clk),.d(0),.we(0));
//assign O28_I28_R1_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O28_I28_R1_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O28_I28_R1_C110_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O28_I28_R1_C110_rom_inst (.q(O28_I28_R1_C1_SM1 ),.address(input_fmap_28[39:32]),.clock  (clk));
logic [11-1:0] O28_I28_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O28_I28_R1_C23_rom_inst (.q(O28_I28_R1_C2_SM1 ),.address(input_fmap_28[47:40]),.clk(clk),.d(0),.we(0));
//assign O28_I28_R1_C2_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O28_I28_R1_C2_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O28_I28_R1_C23_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O28_I28_R1_C23_rom_inst (.q(O28_I28_R1_C2_SM1 ),.address(input_fmap_28[47:40]),.clock  (clk));
logic [10-1:0] O28_I28_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_dw_O28_I28_R2_C01_rom_inst (.q(O28_I28_R2_C0_SM1 ),.address(input_fmap_28[55:48]),.clk(clk),.d(0),.we(0));
//assign O28_I28_R2_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O28_I28_R2_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O28_I28_R2_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_dw_O28_I28_R2_C01_rom_inst (.q(O28_I28_R2_C0_SM1 ),.address(input_fmap_28[55:48]),.clock  (clk));
logic [13-1:0] O28_I28_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O28_I28_R2_C112_rom_inst (.q(O28_I28_R2_C1_SM1 ),.address(input_fmap_28[63:56]),.clk(clk),.d(0),.we(0));
//assign O28_I28_R2_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O28_I28_R2_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O28_I28_R2_C112_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O28_I28_R2_C112_rom_inst (.q(O28_I28_R2_C1_SM1 ),.address(input_fmap_28[63:56]),.clock  (clk));
logic [12-1:0] O28_I28_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O28_I28_R2_C24_rom_inst (.q(O28_I28_R2_C2_SM1 ),.address(input_fmap_28[71:64]),.clk(clk),.d(0),.we(0));
//assign O28_I28_R2_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O28_I28_R2_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O28_I28_R2_C24_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O28_I28_R2_C24_rom_inst (.q(O28_I28_R2_C2_SM1 ),.address(input_fmap_28[71:64]),.clock  (clk));
logic [13-1:0] O29_I29_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O29_I29_R0_C010_rom_inst (.q(O29_I29_R0_C0_SM1 ),.address(input_fmap_29[7:0]),.clk(clk),.d(0),.we(0));
//assign O29_I29_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O29_I29_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O29_I29_R0_C010_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O29_I29_R0_C010_rom_inst (.q(O29_I29_R0_C0_SM1 ),.address(input_fmap_29[7:0]),.clock  (clk));
logic [13-1:0] O29_I29_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O29_I29_R0_C110_rom_inst (.q(O29_I29_R0_C1_SM1 ),.address(input_fmap_29[15:8]),.clk(clk),.d(0),.we(0));
//assign O29_I29_R0_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O29_I29_R0_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O29_I29_R0_C110_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O29_I29_R0_C110_rom_inst (.q(O29_I29_R0_C1_SM1 ),.address(input_fmap_29[15:8]),.clock  (clk));
logic [10-1:0] O29_I29_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_dw_O29_I29_R0_C21_rom_inst (.q(O29_I29_R0_C2_SM1 ),.address(input_fmap_29[23:16]),.clk(clk),.d(0),.we(0));
//assign O29_I29_R0_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O29_I29_R0_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O29_I29_R0_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_dw_O29_I29_R0_C21_rom_inst (.q(O29_I29_R0_C2_SM1 ),.address(input_fmap_29[23:16]),.clock  (clk));
logic [13-1:0] O29_I29_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O29_I29_R1_C010_rom_inst (.q(O29_I29_R1_C0_SM1 ),.address(input_fmap_29[31:24]),.clk(clk),.d(0),.we(0));
//assign O29_I29_R1_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O29_I29_R1_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O29_I29_R1_C010_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O29_I29_R1_C010_rom_inst (.q(O29_I29_R1_C0_SM1 ),.address(input_fmap_29[31:24]),.clock  (clk));
logic [15-1:0] O29_I29_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(15),.INIT_FILE("deepfreeze_rom/deepfreeze_8_15.txt"))
    conv5_dw_O29_I29_R1_C136_rom_inst (.q(O29_I29_R1_C1_SM1 ),.address(input_fmap_29[39:32]),.clk(clk),.d(0),.we(0));
//assign O29_I29_R1_C1_SM1  = 15'h1234;
//always@(posedge clk) begin 
//O29_I29_R1_C1_SM1  <= 15'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O29_I29_R1_C136_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(15))
//    conv5_dw_O29_I29_R1_C136_rom_inst (.q(O29_I29_R1_C1_SM1 ),.address(input_fmap_29[39:32]),.clock  (clk));
logic [13-1:0] O29_I29_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O29_I29_R1_C210_rom_inst (.q(O29_I29_R1_C2_SM1 ),.address(input_fmap_29[47:40]),.clk(clk),.d(0),.we(0));
//assign O29_I29_R1_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O29_I29_R1_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O29_I29_R1_C210_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O29_I29_R1_C210_rom_inst (.q(O29_I29_R1_C2_SM1 ),.address(input_fmap_29[47:40]),.clock  (clk));
logic [11-1:0] O29_I29_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O29_I29_R2_C03_rom_inst (.q(O29_I29_R2_C0_SM1 ),.address(input_fmap_29[55:48]),.clk(clk),.d(0),.we(0));
//assign O29_I29_R2_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O29_I29_R2_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O29_I29_R2_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O29_I29_R2_C03_rom_inst (.q(O29_I29_R2_C0_SM1 ),.address(input_fmap_29[55:48]),.clock  (clk));
logic [13-1:0] O29_I29_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O29_I29_R2_C110_rom_inst (.q(O29_I29_R2_C1_SM1 ),.address(input_fmap_29[63:56]),.clk(clk),.d(0),.we(0));
//assign O29_I29_R2_C1_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O29_I29_R2_C1_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O29_I29_R2_C110_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O29_I29_R2_C110_rom_inst (.q(O29_I29_R2_C1_SM1 ),.address(input_fmap_29[63:56]),.clock  (clk));
logic [13-1:0] O29_I29_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O29_I29_R2_C211_rom_inst (.q(O29_I29_R2_C2_SM1 ),.address(input_fmap_29[71:64]),.clk(clk),.d(0),.we(0));
//assign O29_I29_R2_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O29_I29_R2_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O29_I29_R2_C211_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O29_I29_R2_C211_rom_inst (.q(O29_I29_R2_C2_SM1 ),.address(input_fmap_29[71:64]),.clock  (clk));
logic [13-1:0] O30_I30_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O30_I30_R0_C013_rom_inst (.q(O30_I30_R0_C0_SM1 ),.address(input_fmap_30[7:0]),.clk(clk),.d(0),.we(0));
//assign O30_I30_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O30_I30_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O30_I30_R0_C013_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O30_I30_R0_C013_rom_inst (.q(O30_I30_R0_C0_SM1 ),.address(input_fmap_30[7:0]),.clock  (clk));
logic [12-1:0] O30_I30_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O30_I30_R0_C17_rom_inst (.q(O30_I30_R0_C1_SM1 ),.address(input_fmap_30[15:8]),.clk(clk),.d(0),.we(0));
//assign O30_I30_R0_C1_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O30_I30_R0_C1_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O30_I30_R0_C17_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O30_I30_R0_C17_rom_inst (.q(O30_I30_R0_C1_SM1 ),.address(input_fmap_30[15:8]),.clock  (clk));
logic [13-1:0] O30_I30_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O30_I30_R0_C28_rom_inst (.q(O30_I30_R0_C2_SM1 ),.address(input_fmap_30[23:16]),.clk(clk),.d(0),.we(0));
//assign O30_I30_R0_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O30_I30_R0_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O30_I30_R0_C28_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O30_I30_R0_C28_rom_inst (.q(O30_I30_R0_C2_SM1 ),.address(input_fmap_30[23:16]),.clock  (clk));
logic [14-1:0] O30_I30_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv5_dw_O30_I30_R1_C028_rom_inst (.q(O30_I30_R1_C0_SM1 ),.address(input_fmap_30[31:24]),.clk(clk),.d(0),.we(0));
//assign O30_I30_R1_C0_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O30_I30_R1_C0_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O30_I30_R1_C028_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv5_dw_O30_I30_R1_C028_rom_inst (.q(O30_I30_R1_C0_SM1 ),.address(input_fmap_30[31:24]),.clock  (clk));
logic [12-1:0] O30_I30_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O30_I30_R1_C17_rom_inst (.q(O30_I30_R1_C1_SM1 ),.address(input_fmap_30[39:32]),.clk(clk),.d(0),.we(0));
//assign O30_I30_R1_C1_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O30_I30_R1_C1_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O30_I30_R1_C17_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O30_I30_R1_C17_rom_inst (.q(O30_I30_R1_C1_SM1 ),.address(input_fmap_30[39:32]),.clock  (clk));
logic [13-1:0] O30_I30_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O30_I30_R1_C29_rom_inst (.q(O30_I30_R1_C2_SM1 ),.address(input_fmap_30[47:40]),.clk(clk),.d(0),.we(0));
//assign O30_I30_R1_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O30_I30_R1_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O30_I30_R1_C29_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O30_I30_R1_C29_rom_inst (.q(O30_I30_R1_C2_SM1 ),.address(input_fmap_30[47:40]),.clock  (clk));
logic [12-1:0] O30_I30_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O30_I30_R2_C05_rom_inst (.q(O30_I30_R2_C0_SM1 ),.address(input_fmap_30[55:48]),.clk(clk),.d(0),.we(0));
//assign O30_I30_R2_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O30_I30_R2_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O30_I30_R2_C05_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O30_I30_R2_C05_rom_inst (.q(O30_I30_R2_C0_SM1 ),.address(input_fmap_30[55:48]),.clock  (clk));
logic [10-1:0] O30_I30_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_dw_O30_I30_R2_C11_rom_inst (.q(O30_I30_R2_C1_SM1 ),.address(input_fmap_30[63:56]),.clk(clk),.d(0),.we(0));
//assign O30_I30_R2_C1_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O30_I30_R2_C1_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O30_I30_R2_C11_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_dw_O30_I30_R2_C11_rom_inst (.q(O30_I30_R2_C1_SM1 ),.address(input_fmap_30[63:56]),.clock  (clk));
logic [13-1:0] O30_I30_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_dw_O30_I30_R2_C28_rom_inst (.q(O30_I30_R2_C2_SM1 ),.address(input_fmap_30[71:64]),.clk(clk),.d(0),.we(0));
//assign O30_I30_R2_C2_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O30_I30_R2_C2_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O30_I30_R2_C28_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_dw_O30_I30_R2_C28_rom_inst (.q(O30_I30_R2_C2_SM1 ),.address(input_fmap_30[71:64]),.clock  (clk));
logic [10-1:0] O31_I31_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_dw_O31_I31_R0_C01_rom_inst (.q(O31_I31_R0_C0_SM1 ),.address(input_fmap_31[7:0]),.clk(clk),.d(0),.we(0));
//assign O31_I31_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O31_I31_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O31_I31_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_dw_O31_I31_R0_C01_rom_inst (.q(O31_I31_R0_C0_SM1 ),.address(input_fmap_31[7:0]),.clock  (clk));
logic [11-1:0] O31_I31_R0_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O31_I31_R0_C13_rom_inst (.q(O31_I31_R0_C1_SM1 ),.address(input_fmap_31[15:8]),.clk(clk),.d(0),.we(0));
//assign O31_I31_R0_C1_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O31_I31_R0_C1_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O31_I31_R0_C13_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O31_I31_R0_C13_rom_inst (.q(O31_I31_R0_C1_SM1 ),.address(input_fmap_31[15:8]),.clock  (clk));
logic [10-1:0] O31_I31_R0_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_dw_O31_I31_R0_C21_rom_inst (.q(O31_I31_R0_C2_SM1 ),.address(input_fmap_31[23:16]),.clk(clk),.d(0),.we(0));
//assign O31_I31_R0_C2_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O31_I31_R0_C2_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O31_I31_R0_C21_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_dw_O31_I31_R0_C21_rom_inst (.q(O31_I31_R0_C2_SM1 ),.address(input_fmap_31[23:16]),.clock  (clk));
logic [14-1:0] O31_I31_R1_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv5_dw_O31_I31_R1_C021_rom_inst (.q(O31_I31_R1_C0_SM1 ),.address(input_fmap_31[31:24]),.clk(clk),.d(0),.we(0));
//assign O31_I31_R1_C0_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O31_I31_R1_C0_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O31_I31_R1_C021_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv5_dw_O31_I31_R1_C021_rom_inst (.q(O31_I31_R1_C0_SM1 ),.address(input_fmap_31[31:24]),.clock  (clk));
logic [14-1:0] O31_I31_R1_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(14),.INIT_FILE("deepfreeze_rom/deepfreeze_8_14.txt"))
    conv5_dw_O31_I31_R1_C117_rom_inst (.q(O31_I31_R1_C1_SM1 ),.address(input_fmap_31[39:32]),.clk(clk),.d(0),.we(0));
//assign O31_I31_R1_C1_SM1  = 14'h1234;
//always@(posedge clk) begin 
//O31_I31_R1_C1_SM1  <= 14'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O31_I31_R1_C117_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(14))
//    conv5_dw_O31_I31_R1_C117_rom_inst (.q(O31_I31_R1_C1_SM1 ),.address(input_fmap_31[39:32]),.clock  (clk));
logic [12-1:0] O31_I31_R1_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O31_I31_R1_C24_rom_inst (.q(O31_I31_R1_C2_SM1 ),.address(input_fmap_31[47:40]),.clk(clk),.d(0),.we(0));
//assign O31_I31_R1_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O31_I31_R1_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O31_I31_R1_C24_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O31_I31_R1_C24_rom_inst (.q(O31_I31_R1_C2_SM1 ),.address(input_fmap_31[47:40]),.clock  (clk));
logic [11-1:0] O31_I31_R2_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_dw_O31_I31_R2_C02_rom_inst (.q(O31_I31_R2_C0_SM1 ),.address(input_fmap_31[55:48]),.clk(clk),.d(0),.we(0));
//assign O31_I31_R2_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O31_I31_R2_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O31_I31_R2_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_dw_O31_I31_R2_C02_rom_inst (.q(O31_I31_R2_C0_SM1 ),.address(input_fmap_31[55:48]),.clock  (clk));
logic [12-1:0] O31_I31_R2_C1_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O31_I31_R2_C17_rom_inst (.q(O31_I31_R2_C1_SM1 ),.address(input_fmap_31[63:56]),.clk(clk),.d(0),.we(0));
//assign O31_I31_R2_C1_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O31_I31_R2_C1_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O31_I31_R2_C17_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O31_I31_R2_C17_rom_inst (.q(O31_I31_R2_C1_SM1 ),.address(input_fmap_31[63:56]),.clock  (clk));
logic [12-1:0] O31_I31_R2_C2_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_dw_O31_I31_R2_C25_rom_inst (.q(O31_I31_R2_C2_SM1 ),.address(input_fmap_31[71:64]),.clk(clk),.d(0),.we(0));
//assign O31_I31_R2_C2_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O31_I31_R2_C2_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_dw_O31_I31_R2_C25_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_dw_O31_I31_R2_C25_rom_inst (.q(O31_I31_R2_C2_SM1 ),.address(input_fmap_31[71:64]),.clock  (clk));
logic signed [31:0] conv_mac_0;
logic signed [31:0] O0_N0_S0;		always @(posedge clk) O0_N0_S0 <=     O0_I0_R0_C0_SM1   +  O0_I0_R0_C1_SM1  ;
 logic signed [31:0] O0_N2_S0;		always @(posedge clk) O0_N2_S0 <=     O0_I0_R0_C2_SM1   +  O0_I0_R1_C0_SM1  ;
 logic signed [31:0] O0_N4_S0;		always @(posedge clk) O0_N4_S0 <=     O0_I0_R1_C1_SM1   +  O0_I0_R1_C2_SM1  ;
 logic signed [31:0] O0_N6_S0;		always @(posedge clk) O0_N6_S0 <=     O0_I0_R2_C0_SM1   +  O0_I0_R2_C1_SM1  ;
 logic signed [31:0] O0_N8_S0;		always @(posedge clk) O0_N8_S0 <=     O0_I0_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O0_N0_S1;		always @(posedge clk) O0_N0_S1 <=     O0_N0_S0  +  O0_N2_S0 ;
 logic signed [31:0] O0_N2_S1;		always @(posedge clk) O0_N2_S1 <=     O0_N4_S0  +  O0_N6_S0 ;
 logic signed [31:0] O0_N4_S1;		always @(posedge clk) O0_N4_S1 <=     O0_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O0_N0_S2;		always @(posedge clk) O0_N0_S2 <=     O0_N0_S1  +  O0_N2_S1 ;
 logic signed [31:0] O0_N2_S2;		always @(posedge clk) O0_N2_S2 <=     O0_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O0_N0_S3;		always @(posedge clk) O0_N0_S3 <=     O0_N0_S2  +  O0_N2_S2 ;
 assign conv_mac_0 = O0_N0_S3;

logic signed [31:0] conv_mac_1;
logic signed [31:0] O1_N0_S0;		always @(posedge clk) O1_N0_S0 <=     O1_I1_R0_C0_SM1   +  O1_I1_R0_C1_SM1  ;
 logic signed [31:0] O1_N2_S0;		always @(posedge clk) O1_N2_S0 <=     O1_I1_R0_C2_SM1   +  O1_I1_R1_C0_SM1  ;
 logic signed [31:0] O1_N4_S0;		always @(posedge clk) O1_N4_S0 <=     O1_I1_R1_C1_SM1   +  O1_I1_R1_C2_SM1  ;
 logic signed [31:0] O1_N6_S0;		always @(posedge clk) O1_N6_S0 <=     O1_I1_R2_C0_SM1   +  O1_I1_R2_C1_SM1  ;
 logic signed [31:0] O1_N8_S0;		always @(posedge clk) O1_N8_S0 <=     O1_I1_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O1_N0_S1;		always @(posedge clk) O1_N0_S1 <=     O1_N0_S0  +  O1_N2_S0 ;
 logic signed [31:0] O1_N2_S1;		always @(posedge clk) O1_N2_S1 <=     O1_N4_S0  +  O1_N6_S0 ;
 logic signed [31:0] O1_N4_S1;		always @(posedge clk) O1_N4_S1 <=     O1_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O1_N0_S2;		always @(posedge clk) O1_N0_S2 <=     O1_N0_S1  +  O1_N2_S1 ;
 logic signed [31:0] O1_N2_S2;		always @(posedge clk) O1_N2_S2 <=     O1_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O1_N0_S3;		always @(posedge clk) O1_N0_S3 <=     O1_N0_S2  +  O1_N2_S2 ;
 assign conv_mac_1 = O1_N0_S3;

logic signed [31:0] conv_mac_2;
logic signed [31:0] O2_N0_S0;		always @(posedge clk) O2_N0_S0 <=     O2_I2_R0_C0_SM1   +  O2_I2_R0_C1_SM1  ;
 logic signed [31:0] O2_N2_S0;		always @(posedge clk) O2_N2_S0 <=     O2_I2_R0_C2_SM1   +  O2_I2_R1_C0_SM1  ;
 logic signed [31:0] O2_N4_S0;		always @(posedge clk) O2_N4_S0 <=     O2_I2_R1_C1_SM1   +  O2_I2_R1_C2_SM1  ;
 logic signed [31:0] O2_N6_S0;		always @(posedge clk) O2_N6_S0 <=     O2_I2_R2_C0_SM1   +  O2_I2_R2_C1_SM1  ;
 logic signed [31:0] O2_N8_S0;		always @(posedge clk) O2_N8_S0 <=     O2_I2_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O2_N0_S1;		always @(posedge clk) O2_N0_S1 <=     O2_N0_S0  +  O2_N2_S0 ;
 logic signed [31:0] O2_N2_S1;		always @(posedge clk) O2_N2_S1 <=     O2_N4_S0  +  O2_N6_S0 ;
 logic signed [31:0] O2_N4_S1;		always @(posedge clk) O2_N4_S1 <=     O2_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O2_N0_S2;		always @(posedge clk) O2_N0_S2 <=     O2_N0_S1  +  O2_N2_S1 ;
 logic signed [31:0] O2_N2_S2;		always @(posedge clk) O2_N2_S2 <=     O2_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O2_N0_S3;		always @(posedge clk) O2_N0_S3 <=     O2_N0_S2  +  O2_N2_S2 ;
 assign conv_mac_2 = O2_N0_S3;

logic signed [31:0] conv_mac_3;
logic signed [31:0] O3_N0_S0;		always @(posedge clk) O3_N0_S0 <=     O3_I3_R0_C0_SM1   +  O3_I3_R0_C1_SM1  ;
 logic signed [31:0] O3_N2_S0;		always @(posedge clk) O3_N2_S0 <=     O3_I3_R0_C2_SM1   +  O3_I3_R1_C0_SM1  ;
 logic signed [31:0] O3_N4_S0;		always @(posedge clk) O3_N4_S0 <=     O3_I3_R1_C1_SM1   +  O3_I3_R2_C0_SM1  ;
 logic signed [31:0] O3_N6_S0;		always @(posedge clk) O3_N6_S0 <=     O3_I3_R2_C1_SM1   +  O3_I3_R2_C2_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O3_N0_S1;		always @(posedge clk) O3_N0_S1 <=     O3_N0_S0  +  O3_N2_S0 ;
 logic signed [31:0] O3_N2_S1;		always @(posedge clk) O3_N2_S1 <=     O3_N4_S0  +  O3_N6_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O3_N0_S2;		always @(posedge clk) O3_N0_S2 <=     O3_N0_S1  +  O3_N2_S1 ;
 assign conv_mac_3 = O3_N0_S2;

logic signed [31:0] conv_mac_4;
logic signed [31:0] O4_N0_S0;		always @(posedge clk) O4_N0_S0 <=     O4_I4_R0_C0_SM1   +  O4_I4_R0_C1_SM1  ;
 logic signed [31:0] O4_N2_S0;		always @(posedge clk) O4_N2_S0 <=     O4_I4_R0_C2_SM1   +  O4_I4_R1_C0_SM1  ;
 logic signed [31:0] O4_N4_S0;		always @(posedge clk) O4_N4_S0 <=     O4_I4_R1_C1_SM1   +  O4_I4_R1_C2_SM1  ;
 logic signed [31:0] O4_N6_S0;		always @(posedge clk) O4_N6_S0 <=     O4_I4_R2_C0_SM1   +  O4_I4_R2_C1_SM1  ;
 logic signed [31:0] O4_N8_S0;		always @(posedge clk) O4_N8_S0 <=     O4_I4_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O4_N0_S1;		always @(posedge clk) O4_N0_S1 <=     O4_N0_S0  +  O4_N2_S0 ;
 logic signed [31:0] O4_N2_S1;		always @(posedge clk) O4_N2_S1 <=     O4_N4_S0  +  O4_N6_S0 ;
 logic signed [31:0] O4_N4_S1;		always @(posedge clk) O4_N4_S1 <=     O4_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O4_N0_S2;		always @(posedge clk) O4_N0_S2 <=     O4_N0_S1  +  O4_N2_S1 ;
 logic signed [31:0] O4_N2_S2;		always @(posedge clk) O4_N2_S2 <=     O4_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O4_N0_S3;		always @(posedge clk) O4_N0_S3 <=     O4_N0_S2  +  O4_N2_S2 ;
 assign conv_mac_4 = O4_N0_S3;

logic signed [31:0] conv_mac_5;
logic signed [31:0] O5_N0_S0;		always @(posedge clk) O5_N0_S0 <=     O5_I5_R0_C0_SM1   +  O5_I5_R0_C1_SM1  ;
 logic signed [31:0] O5_N2_S0;		always @(posedge clk) O5_N2_S0 <=     O5_I5_R0_C2_SM1   +  O5_I5_R1_C0_SM1  ;
 logic signed [31:0] O5_N4_S0;		always @(posedge clk) O5_N4_S0 <=     O5_I5_R1_C1_SM1   +  O5_I5_R1_C2_SM1  ;
 logic signed [31:0] O5_N6_S0;		always @(posedge clk) O5_N6_S0 <=     O5_I5_R2_C0_SM1   +  O5_I5_R2_C1_SM1  ;
 logic signed [31:0] O5_N8_S0;		always @(posedge clk) O5_N8_S0 <=     O5_I5_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O5_N0_S1;		always @(posedge clk) O5_N0_S1 <=     O5_N0_S0  +  O5_N2_S0 ;
 logic signed [31:0] O5_N2_S1;		always @(posedge clk) O5_N2_S1 <=     O5_N4_S0  +  O5_N6_S0 ;
 logic signed [31:0] O5_N4_S1;		always @(posedge clk) O5_N4_S1 <=     O5_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O5_N0_S2;		always @(posedge clk) O5_N0_S2 <=     O5_N0_S1  +  O5_N2_S1 ;
 logic signed [31:0] O5_N2_S2;		always @(posedge clk) O5_N2_S2 <=     O5_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O5_N0_S3;		always @(posedge clk) O5_N0_S3 <=     O5_N0_S2  +  O5_N2_S2 ;
 assign conv_mac_5 = O5_N0_S3;

logic signed [31:0] conv_mac_6;
logic signed [31:0] O6_N0_S0;		always @(posedge clk) O6_N0_S0 <=     O6_I6_R0_C0_SM1   +  O6_I6_R0_C1_SM1  ;
 logic signed [31:0] O6_N2_S0;		always @(posedge clk) O6_N2_S0 <=     O6_I6_R0_C2_SM1   +  O6_I6_R1_C0_SM1  ;
 logic signed [31:0] O6_N4_S0;		always @(posedge clk) O6_N4_S0 <=     O6_I6_R1_C1_SM1   +  O6_I6_R1_C2_SM1  ;
 logic signed [31:0] O6_N6_S0;		always @(posedge clk) O6_N6_S0 <=     O6_I6_R2_C0_SM1   +  O6_I6_R2_C1_SM1  ;
 logic signed [31:0] O6_N8_S0;		always @(posedge clk) O6_N8_S0 <=     O6_I6_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O6_N0_S1;		always @(posedge clk) O6_N0_S1 <=     O6_N0_S0  +  O6_N2_S0 ;
 logic signed [31:0] O6_N2_S1;		always @(posedge clk) O6_N2_S1 <=     O6_N4_S0  +  O6_N6_S0 ;
 logic signed [31:0] O6_N4_S1;		always @(posedge clk) O6_N4_S1 <=     O6_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O6_N0_S2;		always @(posedge clk) O6_N0_S2 <=     O6_N0_S1  +  O6_N2_S1 ;
 logic signed [31:0] O6_N2_S2;		always @(posedge clk) O6_N2_S2 <=     O6_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O6_N0_S3;		always @(posedge clk) O6_N0_S3 <=     O6_N0_S2  +  O6_N2_S2 ;
 assign conv_mac_6 = O6_N0_S3;

logic signed [31:0] conv_mac_7;
logic signed [31:0] O7_N0_S0;		always @(posedge clk) O7_N0_S0 <=     O7_I7_R0_C0_SM1   +  O7_I7_R0_C1_SM1  ;
 logic signed [31:0] O7_N2_S0;		always @(posedge clk) O7_N2_S0 <=     O7_I7_R0_C2_SM1   +  O7_I7_R1_C0_SM1  ;
 logic signed [31:0] O7_N4_S0;		always @(posedge clk) O7_N4_S0 <=     O7_I7_R1_C1_SM1   +  O7_I7_R1_C2_SM1  ;
 logic signed [31:0] O7_N6_S0;		always @(posedge clk) O7_N6_S0 <=     O7_I7_R2_C0_SM1   +  O7_I7_R2_C1_SM1  ;
 logic signed [31:0] O7_N8_S0;		always @(posedge clk) O7_N8_S0 <=     O7_I7_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O7_N0_S1;		always @(posedge clk) O7_N0_S1 <=     O7_N0_S0  +  O7_N2_S0 ;
 logic signed [31:0] O7_N2_S1;		always @(posedge clk) O7_N2_S1 <=     O7_N4_S0  +  O7_N6_S0 ;
 logic signed [31:0] O7_N4_S1;		always @(posedge clk) O7_N4_S1 <=     O7_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O7_N0_S2;		always @(posedge clk) O7_N0_S2 <=     O7_N0_S1  +  O7_N2_S1 ;
 logic signed [31:0] O7_N2_S2;		always @(posedge clk) O7_N2_S2 <=     O7_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O7_N0_S3;		always @(posedge clk) O7_N0_S3 <=     O7_N0_S2  +  O7_N2_S2 ;
 assign conv_mac_7 = O7_N0_S3;

logic signed [31:0] conv_mac_8;
logic signed [31:0] O8_N0_S0;		always @(posedge clk) O8_N0_S0 <=     O8_I8_R0_C0_SM1   +  O8_I8_R0_C1_SM1  ;
 logic signed [31:0] O8_N2_S0;		always @(posedge clk) O8_N2_S0 <=     O8_I8_R0_C2_SM1   +  O8_I8_R1_C0_SM1  ;
 logic signed [31:0] O8_N4_S0;		always @(posedge clk) O8_N4_S0 <=     O8_I8_R1_C1_SM1   +  O8_I8_R2_C0_SM1  ;
 logic signed [31:0] O8_N6_S0;		always @(posedge clk) O8_N6_S0 <=     O8_I8_R2_C1_SM1   +  O8_I8_R2_C2_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O8_N0_S1;		always @(posedge clk) O8_N0_S1 <=     O8_N0_S0  +  O8_N2_S0 ;
 logic signed [31:0] O8_N2_S1;		always @(posedge clk) O8_N2_S1 <=     O8_N4_S0  +  O8_N6_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O8_N0_S2;		always @(posedge clk) O8_N0_S2 <=     O8_N0_S1  +  O8_N2_S1 ;
 assign conv_mac_8 = O8_N0_S2;

logic signed [31:0] conv_mac_9;
logic signed [31:0] O9_N0_S0;		always @(posedge clk) O9_N0_S0 <=     O9_I9_R0_C0_SM1   +  O9_I9_R0_C1_SM1  ;
 logic signed [31:0] O9_N2_S0;		always @(posedge clk) O9_N2_S0 <=     O9_I9_R0_C2_SM1   +  O9_I9_R1_C0_SM1  ;
 logic signed [31:0] O9_N4_S0;		always @(posedge clk) O9_N4_S0 <=     O9_I9_R1_C1_SM1   +  O9_I9_R1_C2_SM1  ;
 logic signed [31:0] O9_N6_S0;		always @(posedge clk) O9_N6_S0 <=     O9_I9_R2_C0_SM1   +  O9_I9_R2_C1_SM1  ;
 logic signed [31:0] O9_N8_S0;		always @(posedge clk) O9_N8_S0 <=     O9_I9_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O9_N0_S1;		always @(posedge clk) O9_N0_S1 <=     O9_N0_S0  +  O9_N2_S0 ;
 logic signed [31:0] O9_N2_S1;		always @(posedge clk) O9_N2_S1 <=     O9_N4_S0  +  O9_N6_S0 ;
 logic signed [31:0] O9_N4_S1;		always @(posedge clk) O9_N4_S1 <=     O9_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O9_N0_S2;		always @(posedge clk) O9_N0_S2 <=     O9_N0_S1  +  O9_N2_S1 ;
 logic signed [31:0] O9_N2_S2;		always @(posedge clk) O9_N2_S2 <=     O9_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O9_N0_S3;		always @(posedge clk) O9_N0_S3 <=     O9_N0_S2  +  O9_N2_S2 ;
 assign conv_mac_9 = O9_N0_S3;

logic signed [31:0] conv_mac_10;
logic signed [31:0] O10_N0_S0;		always @(posedge clk) O10_N0_S0 <=     O10_I10_R0_C0_SM1   +  O10_I10_R0_C1_SM1  ;
 logic signed [31:0] O10_N2_S0;		always @(posedge clk) O10_N2_S0 <=     O10_I10_R0_C2_SM1   +  O10_I10_R1_C0_SM1  ;
 logic signed [31:0] O10_N4_S0;		always @(posedge clk) O10_N4_S0 <=     O10_I10_R1_C1_SM1   +  O10_I10_R1_C2_SM1  ;
 logic signed [31:0] O10_N6_S0;		always @(posedge clk) O10_N6_S0 <=     O10_I10_R2_C0_SM1   +  O10_I10_R2_C1_SM1  ;
 logic signed [31:0] O10_N8_S0;		always @(posedge clk) O10_N8_S0 <=     O10_I10_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O10_N0_S1;		always @(posedge clk) O10_N0_S1 <=     O10_N0_S0  +  O10_N2_S0 ;
 logic signed [31:0] O10_N2_S1;		always @(posedge clk) O10_N2_S1 <=     O10_N4_S0  +  O10_N6_S0 ;
 logic signed [31:0] O10_N4_S1;		always @(posedge clk) O10_N4_S1 <=     O10_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O10_N0_S2;		always @(posedge clk) O10_N0_S2 <=     O10_N0_S1  +  O10_N2_S1 ;
 logic signed [31:0] O10_N2_S2;		always @(posedge clk) O10_N2_S2 <=     O10_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O10_N0_S3;		always @(posedge clk) O10_N0_S3 <=     O10_N0_S2  +  O10_N2_S2 ;
 assign conv_mac_10 = O10_N0_S3;

logic signed [31:0] conv_mac_11;
logic signed [31:0] O11_N0_S0;		always @(posedge clk) O11_N0_S0 <=     O11_I11_R0_C0_SM1   +  O11_I11_R0_C2_SM1  ;
 logic signed [31:0] O11_N2_S0;		always @(posedge clk) O11_N2_S0 <=     O11_I11_R1_C0_SM1   +  O11_I11_R1_C1_SM1  ;
 logic signed [31:0] O11_N4_S0;		always @(posedge clk) O11_N4_S0 <=     O11_I11_R1_C2_SM1   +  O11_I11_R2_C0_SM1  ;
 logic signed [31:0] O11_N6_S0;		always @(posedge clk) O11_N6_S0 <=     O11_I11_R2_C1_SM1   +  O11_I11_R2_C2_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O11_N0_S1;		always @(posedge clk) O11_N0_S1 <=     O11_N0_S0  +  O11_N2_S0 ;
 logic signed [31:0] O11_N2_S1;		always @(posedge clk) O11_N2_S1 <=     O11_N4_S0  +  O11_N6_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O11_N0_S2;		always @(posedge clk) O11_N0_S2 <=     O11_N0_S1  +  O11_N2_S1 ;
 assign conv_mac_11 = O11_N0_S2;

logic signed [31:0] conv_mac_12;
logic signed [31:0] O12_N0_S0;		always @(posedge clk) O12_N0_S0 <=     O12_I12_R0_C0_SM1   +  O12_I12_R0_C1_SM1  ;
 logic signed [31:0] O12_N2_S0;		always @(posedge clk) O12_N2_S0 <=     O12_I12_R0_C2_SM1   +  O12_I12_R1_C0_SM1  ;
 logic signed [31:0] O12_N4_S0;		always @(posedge clk) O12_N4_S0 <=     O12_I12_R1_C1_SM1   +  O12_I12_R1_C2_SM1  ;
 logic signed [31:0] O12_N6_S0;		always @(posedge clk) O12_N6_S0 <=     O12_I12_R2_C0_SM1   +  O12_I12_R2_C1_SM1  ;
 logic signed [31:0] O12_N8_S0;		always @(posedge clk) O12_N8_S0 <=     O12_I12_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O12_N0_S1;		always @(posedge clk) O12_N0_S1 <=     O12_N0_S0  +  O12_N2_S0 ;
 logic signed [31:0] O12_N2_S1;		always @(posedge clk) O12_N2_S1 <=     O12_N4_S0  +  O12_N6_S0 ;
 logic signed [31:0] O12_N4_S1;		always @(posedge clk) O12_N4_S1 <=     O12_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O12_N0_S2;		always @(posedge clk) O12_N0_S2 <=     O12_N0_S1  +  O12_N2_S1 ;
 logic signed [31:0] O12_N2_S2;		always @(posedge clk) O12_N2_S2 <=     O12_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O12_N0_S3;		always @(posedge clk) O12_N0_S3 <=     O12_N0_S2  +  O12_N2_S2 ;
 assign conv_mac_12 = O12_N0_S3;

logic signed [31:0] conv_mac_13;
logic signed [31:0] O13_N0_S0;		always @(posedge clk) O13_N0_S0 <=     O13_I13_R0_C0_SM1   +  O13_I13_R0_C1_SM1  ;
 logic signed [31:0] O13_N2_S0;		always @(posedge clk) O13_N2_S0 <=     O13_I13_R0_C2_SM1   +  O13_I13_R1_C0_SM1  ;
 logic signed [31:0] O13_N4_S0;		always @(posedge clk) O13_N4_S0 <=     O13_I13_R1_C1_SM1   +  O13_I13_R1_C2_SM1  ;
 logic signed [31:0] O13_N6_S0;		always @(posedge clk) O13_N6_S0 <=     O13_I13_R2_C0_SM1   +  O13_I13_R2_C1_SM1  ;
 logic signed [31:0] O13_N8_S0;		always @(posedge clk) O13_N8_S0 <=     O13_I13_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O13_N0_S1;		always @(posedge clk) O13_N0_S1 <=     O13_N0_S0  +  O13_N2_S0 ;
 logic signed [31:0] O13_N2_S1;		always @(posedge clk) O13_N2_S1 <=     O13_N4_S0  +  O13_N6_S0 ;
 logic signed [31:0] O13_N4_S1;		always @(posedge clk) O13_N4_S1 <=     O13_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O13_N0_S2;		always @(posedge clk) O13_N0_S2 <=     O13_N0_S1  +  O13_N2_S1 ;
 logic signed [31:0] O13_N2_S2;		always @(posedge clk) O13_N2_S2 <=     O13_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O13_N0_S3;		always @(posedge clk) O13_N0_S3 <=     O13_N0_S2  +  O13_N2_S2 ;
 assign conv_mac_13 = O13_N0_S3;

logic signed [31:0] conv_mac_14;
logic signed [31:0] O14_N0_S0;		always @(posedge clk) O14_N0_S0 <=     O14_I14_R0_C1_SM1   +  O14_I14_R0_C2_SM1  ;
 logic signed [31:0] O14_N2_S0;		always @(posedge clk) O14_N2_S0 <=     O14_I14_R1_C0_SM1   +  O14_I14_R1_C1_SM1  ;
 logic signed [31:0] O14_N4_S0;		always @(posedge clk) O14_N4_S0 <=     O14_I14_R1_C2_SM1   +  O14_I14_R2_C0_SM1  ;
 logic signed [31:0] O14_N6_S0;		always @(posedge clk) O14_N6_S0 <=     O14_I14_R2_C1_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O14_N0_S1;		always @(posedge clk) O14_N0_S1 <=     O14_N0_S0  +  O14_N2_S0 ;
 logic signed [31:0] O14_N2_S1;		always @(posedge clk) O14_N2_S1 <=     O14_N4_S0  +  O14_N6_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O14_N0_S2;		always @(posedge clk) O14_N0_S2 <=     O14_N0_S1  +  O14_N2_S1 ;
 assign conv_mac_14 = O14_N0_S2;

logic signed [31:0] conv_mac_15;
logic signed [31:0] O15_N0_S0;		always @(posedge clk) O15_N0_S0 <=     O15_I15_R0_C0_SM1   +  O15_I15_R0_C2_SM1  ;
 logic signed [31:0] O15_N2_S0;		always @(posedge clk) O15_N2_S0 <=     O15_I15_R1_C0_SM1   +  O15_I15_R1_C1_SM1  ;
 logic signed [31:0] O15_N4_S0;		always @(posedge clk) O15_N4_S0 <=     O15_I15_R1_C2_SM1   +  O15_I15_R2_C0_SM1  ;
 logic signed [31:0] O15_N6_S0;		always @(posedge clk) O15_N6_S0 <=     O15_I15_R2_C1_SM1   +  O15_I15_R2_C2_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O15_N0_S1;		always @(posedge clk) O15_N0_S1 <=     O15_N0_S0  +  O15_N2_S0 ;
 logic signed [31:0] O15_N2_S1;		always @(posedge clk) O15_N2_S1 <=     O15_N4_S0  +  O15_N6_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O15_N0_S2;		always @(posedge clk) O15_N0_S2 <=     O15_N0_S1  +  O15_N2_S1 ;
 assign conv_mac_15 = O15_N0_S2;

logic signed [31:0] conv_mac_16;
logic signed [31:0] O16_N0_S0;		always @(posedge clk) O16_N0_S0 <=     O16_I16_R0_C0_SM1   +  O16_I16_R0_C1_SM1  ;
 logic signed [31:0] O16_N2_S0;		always @(posedge clk) O16_N2_S0 <=     O16_I16_R0_C2_SM1   +  O16_I16_R1_C0_SM1  ;
 logic signed [31:0] O16_N4_S0;		always @(posedge clk) O16_N4_S0 <=     O16_I16_R1_C1_SM1   +  O16_I16_R1_C2_SM1  ;
 logic signed [31:0] O16_N6_S0;		always @(posedge clk) O16_N6_S0 <=     O16_I16_R2_C1_SM1   +  O16_I16_R2_C2_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O16_N0_S1;		always @(posedge clk) O16_N0_S1 <=     O16_N0_S0  +  O16_N2_S0 ;
 logic signed [31:0] O16_N2_S1;		always @(posedge clk) O16_N2_S1 <=     O16_N4_S0  +  O16_N6_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O16_N0_S2;		always @(posedge clk) O16_N0_S2 <=     O16_N0_S1  +  O16_N2_S1 ;
 assign conv_mac_16 = O16_N0_S2;

logic signed [31:0] conv_mac_17;
logic signed [31:0] O17_N0_S0;		always @(posedge clk) O17_N0_S0 <=     O17_I17_R0_C0_SM1   +  O17_I17_R0_C1_SM1  ;
 logic signed [31:0] O17_N2_S0;		always @(posedge clk) O17_N2_S0 <=     O17_I17_R0_C2_SM1   +  O17_I17_R1_C0_SM1  ;
 logic signed [31:0] O17_N4_S0;		always @(posedge clk) O17_N4_S0 <=     O17_I17_R1_C1_SM1   +  O17_I17_R1_C2_SM1  ;
 logic signed [31:0] O17_N6_S0;		always @(posedge clk) O17_N6_S0 <=     O17_I17_R2_C0_SM1   +  O17_I17_R2_C1_SM1  ;
 logic signed [31:0] O17_N8_S0;		always @(posedge clk) O17_N8_S0 <=     O17_I17_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O17_N0_S1;		always @(posedge clk) O17_N0_S1 <=     O17_N0_S0  +  O17_N2_S0 ;
 logic signed [31:0] O17_N2_S1;		always @(posedge clk) O17_N2_S1 <=     O17_N4_S0  +  O17_N6_S0 ;
 logic signed [31:0] O17_N4_S1;		always @(posedge clk) O17_N4_S1 <=     O17_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O17_N0_S2;		always @(posedge clk) O17_N0_S2 <=     O17_N0_S1  +  O17_N2_S1 ;
 logic signed [31:0] O17_N2_S2;		always @(posedge clk) O17_N2_S2 <=     O17_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O17_N0_S3;		always @(posedge clk) O17_N0_S3 <=     O17_N0_S2  +  O17_N2_S2 ;
 assign conv_mac_17 = O17_N0_S3;

logic signed [31:0] conv_mac_18;
logic signed [31:0] O18_N0_S0;		always @(posedge clk) O18_N0_S0 <=     O18_I18_R0_C0_SM1   +  O18_I18_R0_C1_SM1  ;
 logic signed [31:0] O18_N2_S0;		always @(posedge clk) O18_N2_S0 <=     O18_I18_R0_C2_SM1   +  O18_I18_R1_C0_SM1  ;
 logic signed [31:0] O18_N4_S0;		always @(posedge clk) O18_N4_S0 <=     O18_I18_R1_C1_SM1   +  O18_I18_R1_C2_SM1  ;
 logic signed [31:0] O18_N6_S0;		always @(posedge clk) O18_N6_S0 <=     O18_I18_R2_C0_SM1   +  O18_I18_R2_C1_SM1  ;
 logic signed [31:0] O18_N8_S0;		always @(posedge clk) O18_N8_S0 <=     O18_I18_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O18_N0_S1;		always @(posedge clk) O18_N0_S1 <=     O18_N0_S0  +  O18_N2_S0 ;
 logic signed [31:0] O18_N2_S1;		always @(posedge clk) O18_N2_S1 <=     O18_N4_S0  +  O18_N6_S0 ;
 logic signed [31:0] O18_N4_S1;		always @(posedge clk) O18_N4_S1 <=     O18_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O18_N0_S2;		always @(posedge clk) O18_N0_S2 <=     O18_N0_S1  +  O18_N2_S1 ;
 logic signed [31:0] O18_N2_S2;		always @(posedge clk) O18_N2_S2 <=     O18_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O18_N0_S3;		always @(posedge clk) O18_N0_S3 <=     O18_N0_S2  +  O18_N2_S2 ;
 assign conv_mac_18 = O18_N0_S3;

logic signed [31:0] conv_mac_19;
logic signed [31:0] O19_N0_S0;		always @(posedge clk) O19_N0_S0 <=     O19_I19_R0_C0_SM1   +  O19_I19_R0_C1_SM1  ;
 logic signed [31:0] O19_N2_S0;		always @(posedge clk) O19_N2_S0 <=     O19_I19_R0_C2_SM1   +  O19_I19_R1_C0_SM1  ;
 logic signed [31:0] O19_N4_S0;		always @(posedge clk) O19_N4_S0 <=     O19_I19_R1_C1_SM1   +  O19_I19_R1_C2_SM1  ;
 logic signed [31:0] O19_N6_S0;		always @(posedge clk) O19_N6_S0 <=     O19_I19_R2_C0_SM1   +  O19_I19_R2_C1_SM1  ;
 logic signed [31:0] O19_N8_S0;		always @(posedge clk) O19_N8_S0 <=     O19_I19_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O19_N0_S1;		always @(posedge clk) O19_N0_S1 <=     O19_N0_S0  +  O19_N2_S0 ;
 logic signed [31:0] O19_N2_S1;		always @(posedge clk) O19_N2_S1 <=     O19_N4_S0  +  O19_N6_S0 ;
 logic signed [31:0] O19_N4_S1;		always @(posedge clk) O19_N4_S1 <=     O19_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O19_N0_S2;		always @(posedge clk) O19_N0_S2 <=     O19_N0_S1  +  O19_N2_S1 ;
 logic signed [31:0] O19_N2_S2;		always @(posedge clk) O19_N2_S2 <=     O19_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O19_N0_S3;		always @(posedge clk) O19_N0_S3 <=     O19_N0_S2  +  O19_N2_S2 ;
 assign conv_mac_19 = O19_N0_S3;

logic signed [31:0] conv_mac_20;
logic signed [31:0] O20_N0_S0;		always @(posedge clk) O20_N0_S0 <=     O20_I20_R0_C0_SM1   +  O20_I20_R0_C1_SM1  ;
 logic signed [31:0] O20_N2_S0;		always @(posedge clk) O20_N2_S0 <=     O20_I20_R0_C2_SM1   +  O20_I20_R1_C0_SM1  ;
 logic signed [31:0] O20_N4_S0;		always @(posedge clk) O20_N4_S0 <=     O20_I20_R1_C1_SM1   +  O20_I20_R1_C2_SM1  ;
 logic signed [31:0] O20_N6_S0;		always @(posedge clk) O20_N6_S0 <=     O20_I20_R2_C0_SM1   +  O20_I20_R2_C1_SM1  ;
 logic signed [31:0] O20_N8_S0;		always @(posedge clk) O20_N8_S0 <=     O20_I20_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O20_N0_S1;		always @(posedge clk) O20_N0_S1 <=     O20_N0_S0  +  O20_N2_S0 ;
 logic signed [31:0] O20_N2_S1;		always @(posedge clk) O20_N2_S1 <=     O20_N4_S0  +  O20_N6_S0 ;
 logic signed [31:0] O20_N4_S1;		always @(posedge clk) O20_N4_S1 <=     O20_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O20_N0_S2;		always @(posedge clk) O20_N0_S2 <=     O20_N0_S1  +  O20_N2_S1 ;
 logic signed [31:0] O20_N2_S2;		always @(posedge clk) O20_N2_S2 <=     O20_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O20_N0_S3;		always @(posedge clk) O20_N0_S3 <=     O20_N0_S2  +  O20_N2_S2 ;
 assign conv_mac_20 = O20_N0_S3;

logic signed [31:0] conv_mac_21;
logic signed [31:0] O21_N0_S0;		always @(posedge clk) O21_N0_S0 <=     O21_I21_R0_C0_SM1   +  O21_I21_R0_C1_SM1  ;
 logic signed [31:0] O21_N2_S0;		always @(posedge clk) O21_N2_S0 <=     O21_I21_R0_C2_SM1   +  O21_I21_R1_C0_SM1  ;
 logic signed [31:0] O21_N4_S0;		always @(posedge clk) O21_N4_S0 <=     O21_I21_R1_C1_SM1   +  O21_I21_R1_C2_SM1  ;
 logic signed [31:0] O21_N6_S0;		always @(posedge clk) O21_N6_S0 <=     O21_I21_R2_C0_SM1   +  O21_I21_R2_C1_SM1  ;
 logic signed [31:0] O21_N8_S0;		always @(posedge clk) O21_N8_S0 <=     O21_I21_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O21_N0_S1;		always @(posedge clk) O21_N0_S1 <=     O21_N0_S0  +  O21_N2_S0 ;
 logic signed [31:0] O21_N2_S1;		always @(posedge clk) O21_N2_S1 <=     O21_N4_S0  +  O21_N6_S0 ;
 logic signed [31:0] O21_N4_S1;		always @(posedge clk) O21_N4_S1 <=     O21_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O21_N0_S2;		always @(posedge clk) O21_N0_S2 <=     O21_N0_S1  +  O21_N2_S1 ;
 logic signed [31:0] O21_N2_S2;		always @(posedge clk) O21_N2_S2 <=     O21_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O21_N0_S3;		always @(posedge clk) O21_N0_S3 <=     O21_N0_S2  +  O21_N2_S2 ;
 assign conv_mac_21 = O21_N0_S3;

logic signed [31:0] conv_mac_22;
logic signed [31:0] O22_N0_S0;		always @(posedge clk) O22_N0_S0 <=     O22_I22_R0_C0_SM1   +  O22_I22_R0_C1_SM1  ;
 logic signed [31:0] O22_N2_S0;		always @(posedge clk) O22_N2_S0 <=     O22_I22_R0_C2_SM1   +  O22_I22_R1_C0_SM1  ;
 logic signed [31:0] O22_N4_S0;		always @(posedge clk) O22_N4_S0 <=     O22_I22_R1_C1_SM1   +  O22_I22_R1_C2_SM1  ;
 logic signed [31:0] O22_N6_S0;		always @(posedge clk) O22_N6_S0 <=     O22_I22_R2_C0_SM1   +  O22_I22_R2_C1_SM1  ;
 logic signed [31:0] O22_N8_S0;		always @(posedge clk) O22_N8_S0 <=     O22_I22_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O22_N0_S1;		always @(posedge clk) O22_N0_S1 <=     O22_N0_S0  +  O22_N2_S0 ;
 logic signed [31:0] O22_N2_S1;		always @(posedge clk) O22_N2_S1 <=     O22_N4_S0  +  O22_N6_S0 ;
 logic signed [31:0] O22_N4_S1;		always @(posedge clk) O22_N4_S1 <=     O22_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O22_N0_S2;		always @(posedge clk) O22_N0_S2 <=     O22_N0_S1  +  O22_N2_S1 ;
 logic signed [31:0] O22_N2_S2;		always @(posedge clk) O22_N2_S2 <=     O22_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O22_N0_S3;		always @(posedge clk) O22_N0_S3 <=     O22_N0_S2  +  O22_N2_S2 ;
 assign conv_mac_22 = O22_N0_S3;

logic signed [31:0] conv_mac_23;
logic signed [31:0] O23_N0_S0;		always @(posedge clk) O23_N0_S0 <=     O23_I23_R0_C0_SM1   +  O23_I23_R0_C1_SM1  ;
 logic signed [31:0] O23_N2_S0;		always @(posedge clk) O23_N2_S0 <=     O23_I23_R0_C2_SM1   +  O23_I23_R1_C0_SM1  ;
 logic signed [31:0] O23_N4_S0;		always @(posedge clk) O23_N4_S0 <=     O23_I23_R1_C1_SM1   +  O23_I23_R1_C2_SM1  ;
 logic signed [31:0] O23_N6_S0;		always @(posedge clk) O23_N6_S0 <=     O23_I23_R2_C0_SM1   +  O23_I23_R2_C1_SM1  ;
 logic signed [31:0] O23_N8_S0;		always @(posedge clk) O23_N8_S0 <=     O23_I23_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O23_N0_S1;		always @(posedge clk) O23_N0_S1 <=     O23_N0_S0  +  O23_N2_S0 ;
 logic signed [31:0] O23_N2_S1;		always @(posedge clk) O23_N2_S1 <=     O23_N4_S0  +  O23_N6_S0 ;
 logic signed [31:0] O23_N4_S1;		always @(posedge clk) O23_N4_S1 <=     O23_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O23_N0_S2;		always @(posedge clk) O23_N0_S2 <=     O23_N0_S1  +  O23_N2_S1 ;
 logic signed [31:0] O23_N2_S2;		always @(posedge clk) O23_N2_S2 <=     O23_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O23_N0_S3;		always @(posedge clk) O23_N0_S3 <=     O23_N0_S2  +  O23_N2_S2 ;
 assign conv_mac_23 = O23_N0_S3;

logic signed [31:0] conv_mac_24;
logic signed [31:0] O24_N0_S0;		always @(posedge clk) O24_N0_S0 <=     O24_I24_R0_C0_SM1   +  O24_I24_R0_C1_SM1  ;
 logic signed [31:0] O24_N2_S0;		always @(posedge clk) O24_N2_S0 <=     O24_I24_R0_C2_SM1   +  O24_I24_R1_C0_SM1  ;
 logic signed [31:0] O24_N4_S0;		always @(posedge clk) O24_N4_S0 <=     O24_I24_R1_C1_SM1   +  O24_I24_R1_C2_SM1  ;
 logic signed [31:0] O24_N6_S0;		always @(posedge clk) O24_N6_S0 <=     O24_I24_R2_C0_SM1   +  O24_I24_R2_C1_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O24_N0_S1;		always @(posedge clk) O24_N0_S1 <=     O24_N0_S0  +  O24_N2_S0 ;
 logic signed [31:0] O24_N2_S1;		always @(posedge clk) O24_N2_S1 <=     O24_N4_S0  +  O24_N6_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O24_N0_S2;		always @(posedge clk) O24_N0_S2 <=     O24_N0_S1  +  O24_N2_S1 ;
 assign conv_mac_24 = O24_N0_S2;

logic signed [31:0] conv_mac_25;
logic signed [31:0] O25_N0_S0;		always @(posedge clk) O25_N0_S0 <=     O25_I25_R0_C0_SM1   +  O25_I25_R0_C1_SM1  ;
 logic signed [31:0] O25_N2_S0;		always @(posedge clk) O25_N2_S0 <=     O25_I25_R0_C2_SM1   +  O25_I25_R1_C0_SM1  ;
 logic signed [31:0] O25_N4_S0;		always @(posedge clk) O25_N4_S0 <=     O25_I25_R1_C1_SM1   +  O25_I25_R1_C2_SM1  ;
 logic signed [31:0] O25_N6_S0;		always @(posedge clk) O25_N6_S0 <=     O25_I25_R2_C0_SM1   +  O25_I25_R2_C1_SM1  ;
 logic signed [31:0] O25_N8_S0;		always @(posedge clk) O25_N8_S0 <=     O25_I25_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O25_N0_S1;		always @(posedge clk) O25_N0_S1 <=     O25_N0_S0  +  O25_N2_S0 ;
 logic signed [31:0] O25_N2_S1;		always @(posedge clk) O25_N2_S1 <=     O25_N4_S0  +  O25_N6_S0 ;
 logic signed [31:0] O25_N4_S1;		always @(posedge clk) O25_N4_S1 <=     O25_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O25_N0_S2;		always @(posedge clk) O25_N0_S2 <=     O25_N0_S1  +  O25_N2_S1 ;
 logic signed [31:0] O25_N2_S2;		always @(posedge clk) O25_N2_S2 <=     O25_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O25_N0_S3;		always @(posedge clk) O25_N0_S3 <=     O25_N0_S2  +  O25_N2_S2 ;
 assign conv_mac_25 = O25_N0_S3;

logic signed [31:0] conv_mac_26;
logic signed [31:0] O26_N0_S0;		always @(posedge clk) O26_N0_S0 <=     O26_I26_R0_C0_SM1   +  O26_I26_R0_C1_SM1  ;
 logic signed [31:0] O26_N2_S0;		always @(posedge clk) O26_N2_S0 <=     O26_I26_R0_C2_SM1   +  O26_I26_R1_C0_SM1  ;
 logic signed [31:0] O26_N4_S0;		always @(posedge clk) O26_N4_S0 <=     O26_I26_R1_C1_SM1   +  O26_I26_R1_C2_SM1  ;
 logic signed [31:0] O26_N6_S0;		always @(posedge clk) O26_N6_S0 <=     O26_I26_R2_C0_SM1   +  O26_I26_R2_C1_SM1  ;
 logic signed [31:0] O26_N8_S0;		always @(posedge clk) O26_N8_S0 <=     O26_I26_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O26_N0_S1;		always @(posedge clk) O26_N0_S1 <=     O26_N0_S0  +  O26_N2_S0 ;
 logic signed [31:0] O26_N2_S1;		always @(posedge clk) O26_N2_S1 <=     O26_N4_S0  +  O26_N6_S0 ;
 logic signed [31:0] O26_N4_S1;		always @(posedge clk) O26_N4_S1 <=     O26_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O26_N0_S2;		always @(posedge clk) O26_N0_S2 <=     O26_N0_S1  +  O26_N2_S1 ;
 logic signed [31:0] O26_N2_S2;		always @(posedge clk) O26_N2_S2 <=     O26_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O26_N0_S3;		always @(posedge clk) O26_N0_S3 <=     O26_N0_S2  +  O26_N2_S2 ;
 assign conv_mac_26 = O26_N0_S3;

logic signed [31:0] conv_mac_27;
logic signed [31:0] O27_N0_S0;		always @(posedge clk) O27_N0_S0 <=     O27_I27_R0_C0_SM1   +  O27_I27_R0_C1_SM1  ;
 logic signed [31:0] O27_N2_S0;		always @(posedge clk) O27_N2_S0 <=     O27_I27_R0_C2_SM1   +  O27_I27_R1_C0_SM1  ;
 logic signed [31:0] O27_N4_S0;		always @(posedge clk) O27_N4_S0 <=     O27_I27_R1_C1_SM1   +  O27_I27_R1_C2_SM1  ;
 logic signed [31:0] O27_N6_S0;		always @(posedge clk) O27_N6_S0 <=     O27_I27_R2_C0_SM1   +  O27_I27_R2_C1_SM1  ;
 logic signed [31:0] O27_N8_S0;		always @(posedge clk) O27_N8_S0 <=     O27_I27_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O27_N0_S1;		always @(posedge clk) O27_N0_S1 <=     O27_N0_S0  +  O27_N2_S0 ;
 logic signed [31:0] O27_N2_S1;		always @(posedge clk) O27_N2_S1 <=     O27_N4_S0  +  O27_N6_S0 ;
 logic signed [31:0] O27_N4_S1;		always @(posedge clk) O27_N4_S1 <=     O27_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O27_N0_S2;		always @(posedge clk) O27_N0_S2 <=     O27_N0_S1  +  O27_N2_S1 ;
 logic signed [31:0] O27_N2_S2;		always @(posedge clk) O27_N2_S2 <=     O27_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O27_N0_S3;		always @(posedge clk) O27_N0_S3 <=     O27_N0_S2  +  O27_N2_S2 ;
 assign conv_mac_27 = O27_N0_S3;

logic signed [31:0] conv_mac_28;
logic signed [31:0] O28_N0_S0;		always @(posedge clk) O28_N0_S0 <=     O28_I28_R0_C0_SM1   +  O28_I28_R0_C1_SM1  ;
 logic signed [31:0] O28_N2_S0;		always @(posedge clk) O28_N2_S0 <=     O28_I28_R1_C0_SM1   +  O28_I28_R1_C1_SM1  ;
 logic signed [31:0] O28_N4_S0;		always @(posedge clk) O28_N4_S0 <=     O28_I28_R1_C2_SM1   +  O28_I28_R2_C0_SM1  ;
 logic signed [31:0] O28_N6_S0;		always @(posedge clk) O28_N6_S0 <=     O28_I28_R2_C1_SM1   +  O28_I28_R2_C2_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O28_N0_S1;		always @(posedge clk) O28_N0_S1 <=     O28_N0_S0  +  O28_N2_S0 ;
 logic signed [31:0] O28_N2_S1;		always @(posedge clk) O28_N2_S1 <=     O28_N4_S0  +  O28_N6_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O28_N0_S2;		always @(posedge clk) O28_N0_S2 <=     O28_N0_S1  +  O28_N2_S1 ;
 assign conv_mac_28 = O28_N0_S2;

logic signed [31:0] conv_mac_29;
logic signed [31:0] O29_N0_S0;		always @(posedge clk) O29_N0_S0 <=     O29_I29_R0_C0_SM1   +  O29_I29_R0_C1_SM1  ;
 logic signed [31:0] O29_N2_S0;		always @(posedge clk) O29_N2_S0 <=     O29_I29_R0_C2_SM1   +  O29_I29_R1_C0_SM1  ;
 logic signed [31:0] O29_N4_S0;		always @(posedge clk) O29_N4_S0 <=     O29_I29_R1_C1_SM1   +  O29_I29_R1_C2_SM1  ;
 logic signed [31:0] O29_N6_S0;		always @(posedge clk) O29_N6_S0 <=     O29_I29_R2_C0_SM1   +  O29_I29_R2_C1_SM1  ;
 logic signed [31:0] O29_N8_S0;		always @(posedge clk) O29_N8_S0 <=     O29_I29_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O29_N0_S1;		always @(posedge clk) O29_N0_S1 <=     O29_N0_S0  +  O29_N2_S0 ;
 logic signed [31:0] O29_N2_S1;		always @(posedge clk) O29_N2_S1 <=     O29_N4_S0  +  O29_N6_S0 ;
 logic signed [31:0] O29_N4_S1;		always @(posedge clk) O29_N4_S1 <=     O29_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O29_N0_S2;		always @(posedge clk) O29_N0_S2 <=     O29_N0_S1  +  O29_N2_S1 ;
 logic signed [31:0] O29_N2_S2;		always @(posedge clk) O29_N2_S2 <=     O29_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O29_N0_S3;		always @(posedge clk) O29_N0_S3 <=     O29_N0_S2  +  O29_N2_S2 ;
 assign conv_mac_29 = O29_N0_S3;

logic signed [31:0] conv_mac_30;
logic signed [31:0] O30_N0_S0;		always @(posedge clk) O30_N0_S0 <=     O30_I30_R0_C0_SM1   +  O30_I30_R0_C1_SM1  ;
 logic signed [31:0] O30_N2_S0;		always @(posedge clk) O30_N2_S0 <=     O30_I30_R0_C2_SM1   +  O30_I30_R1_C0_SM1  ;
 logic signed [31:0] O30_N4_S0;		always @(posedge clk) O30_N4_S0 <=     O30_I30_R1_C1_SM1   +  O30_I30_R1_C2_SM1  ;
 logic signed [31:0] O30_N6_S0;		always @(posedge clk) O30_N6_S0 <=     O30_I30_R2_C0_SM1   +  O30_I30_R2_C1_SM1  ;
 logic signed [31:0] O30_N8_S0;		always @(posedge clk) O30_N8_S0 <=     O30_I30_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O30_N0_S1;		always @(posedge clk) O30_N0_S1 <=     O30_N0_S0  +  O30_N2_S0 ;
 logic signed [31:0] O30_N2_S1;		always @(posedge clk) O30_N2_S1 <=     O30_N4_S0  +  O30_N6_S0 ;
 logic signed [31:0] O30_N4_S1;		always @(posedge clk) O30_N4_S1 <=     O30_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O30_N0_S2;		always @(posedge clk) O30_N0_S2 <=     O30_N0_S1  +  O30_N2_S1 ;
 logic signed [31:0] O30_N2_S2;		always @(posedge clk) O30_N2_S2 <=     O30_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O30_N0_S3;		always @(posedge clk) O30_N0_S3 <=     O30_N0_S2  +  O30_N2_S2 ;
 assign conv_mac_30 = O30_N0_S3;

logic signed [31:0] conv_mac_31;
logic signed [31:0] O31_N0_S0;		always @(posedge clk) O31_N0_S0 <=     O31_I31_R0_C0_SM1   +  O31_I31_R0_C1_SM1  ;
 logic signed [31:0] O31_N2_S0;		always @(posedge clk) O31_N2_S0 <=     O31_I31_R0_C2_SM1   +  O31_I31_R1_C0_SM1  ;
 logic signed [31:0] O31_N4_S0;		always @(posedge clk) O31_N4_S0 <=     O31_I31_R1_C1_SM1   +  O31_I31_R1_C2_SM1  ;
 logic signed [31:0] O31_N6_S0;		always @(posedge clk) O31_N6_S0 <=     O31_I31_R2_C0_SM1   +  O31_I31_R2_C1_SM1  ;
 logic signed [31:0] O31_N8_S0;		always @(posedge clk) O31_N8_S0 <=     O31_I31_R2_C2_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O31_N0_S1;		always @(posedge clk) O31_N0_S1 <=     O31_N0_S0  +  O31_N2_S0 ;
 logic signed [31:0] O31_N2_S1;		always @(posedge clk) O31_N2_S1 <=     O31_N4_S0  +  O31_N6_S0 ;
 logic signed [31:0] O31_N4_S1;		always @(posedge clk) O31_N4_S1 <=     O31_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O31_N0_S2;		always @(posedge clk) O31_N0_S2 <=     O31_N0_S1  +  O31_N2_S1 ;
 logic signed [31:0] O31_N2_S2;		always @(posedge clk) O31_N2_S2 <=     O31_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O31_N0_S3;		always @(posedge clk) O31_N0_S3 <=     O31_N0_S2  +  O31_N2_S2 ;
 assign conv_mac_31 = O31_N0_S3;

logic valid_D1;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D1<= 0 ;
	else valid_D1<=valid;
end
logic valid_D2;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D2<= 0 ;
	else valid_D2<=valid_D1;
end
logic valid_D3;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D3<= 0 ;
	else valid_D3<=valid_D2;
end
logic valid_D4;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D4<= 0 ;
	else valid_D4<=valid_D3;
end
logic valid_D5;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D5<= 0 ;
	else valid_D5<=valid_D4;
end
always_ff @(posedge clk) begin
	if (rstn == 0) ready <= 0 ;
	else ready <=valid_D5;
end
logic [31:0] bias_add_0;
assign bias_add_0 = conv_mac_0 - 4'd4;
logic [31:0] bias_add_1;
assign bias_add_1 = conv_mac_1;
logic [31:0] bias_add_2;
assign bias_add_2 = conv_mac_2 + 7'd49;
logic [31:0] bias_add_3;
assign bias_add_3 = conv_mac_3 + 7'd43;
logic [31:0] bias_add_4;
assign bias_add_4 = conv_mac_4 + 4'd5;
logic [31:0] bias_add_5;
assign bias_add_5 = conv_mac_5;
logic [31:0] bias_add_6;
assign bias_add_6 = conv_mac_6 - 3'd2;
logic [31:0] bias_add_7;
assign bias_add_7 = conv_mac_7 + 7'd38;
logic [31:0] bias_add_8;
assign bias_add_8 = conv_mac_8 - 3'd3;
logic [31:0] bias_add_9;
assign bias_add_9 = conv_mac_9 + 7'd38;
logic [31:0] bias_add_10;
assign bias_add_10 = conv_mac_10 - 4'd5;
logic [31:0] bias_add_11;
assign bias_add_11 = conv_mac_11 + 4'd5;
logic [31:0] bias_add_12;
assign bias_add_12 = conv_mac_12 - 4'd4;
logic [31:0] bias_add_13;
assign bias_add_13 = conv_mac_13 - 4'd4;
logic [31:0] bias_add_14;
assign bias_add_14 = conv_mac_14 + 6'd19;
logic [31:0] bias_add_15;
assign bias_add_15 = conv_mac_15 + 6'd31;
logic [31:0] bias_add_16;
assign bias_add_16 = conv_mac_16 - 5'd14;
logic [31:0] bias_add_17;
assign bias_add_17 = conv_mac_17 + 5'd8;
logic [31:0] bias_add_18;
assign bias_add_18 = conv_mac_18 + 6'd21;
logic [31:0] bias_add_19;
assign bias_add_19 = conv_mac_19 + 4'd5;
logic [31:0] bias_add_20;
assign bias_add_20 = conv_mac_20 + 7'd38;
logic [31:0] bias_add_21;
assign bias_add_21 = conv_mac_21 + 5'd15;
logic [31:0] bias_add_22;
assign bias_add_22 = conv_mac_22 + 3'd2;
logic [31:0] bias_add_23;
assign bias_add_23 = conv_mac_23 + 6'd17;
logic [31:0] bias_add_24;
assign bias_add_24 = conv_mac_24 + 5'd13;
logic [31:0] bias_add_25;
assign bias_add_25 = conv_mac_25 + 8'd67;
logic [31:0] bias_add_26;
assign bias_add_26 = conv_mac_26 + 7'd39;
logic [31:0] bias_add_27;
assign bias_add_27 = conv_mac_27 - 4'd7;
logic [31:0] bias_add_28;
assign bias_add_28 = conv_mac_28 - 6'd19;
logic [31:0] bias_add_29;
assign bias_add_29 = conv_mac_29 + 5'd15;
logic [31:0] bias_add_30;
assign bias_add_30 = conv_mac_30;
logic [31:0] bias_add_31;
assign bias_add_31 = conv_mac_31 + 7'd53;

logic [7:0] relu_0;
assign relu_0[7:0] = (bias_add_0[31]==0) ? ((bias_add_0<3'd6) ? {{bias_add_0[31],bias_add_0[10:4]}} :'d6) : '0;
logic [7:0] relu_1;
assign relu_1[7:0] = (bias_add_1[31]==0) ? ((bias_add_1<3'd6) ? {{bias_add_1[31],bias_add_1[10:4]}} :'d6) : '0;
logic [7:0] relu_2;
assign relu_2[7:0] = (bias_add_2[31]==0) ? ((bias_add_2<3'd6) ? {{bias_add_2[31],bias_add_2[10:4]}} :'d6) : '0;
logic [7:0] relu_3;
assign relu_3[7:0] = (bias_add_3[31]==0) ? ((bias_add_3<3'd6) ? {{bias_add_3[31],bias_add_3[10:4]}} :'d6) : '0;
logic [7:0] relu_4;
assign relu_4[7:0] = (bias_add_4[31]==0) ? ((bias_add_4<3'd6) ? {{bias_add_4[31],bias_add_4[10:4]}} :'d6) : '0;
logic [7:0] relu_5;
assign relu_5[7:0] = (bias_add_5[31]==0) ? ((bias_add_5<3'd6) ? {{bias_add_5[31],bias_add_5[10:4]}} :'d6) : '0;
logic [7:0] relu_6;
assign relu_6[7:0] = (bias_add_6[31]==0) ? ((bias_add_6<3'd6) ? {{bias_add_6[31],bias_add_6[10:4]}} :'d6) : '0;
logic [7:0] relu_7;
assign relu_7[7:0] = (bias_add_7[31]==0) ? ((bias_add_7<3'd6) ? {{bias_add_7[31],bias_add_7[10:4]}} :'d6) : '0;
logic [7:0] relu_8;
assign relu_8[7:0] = (bias_add_8[31]==0) ? ((bias_add_8<3'd6) ? {{bias_add_8[31],bias_add_8[10:4]}} :'d6) : '0;
logic [7:0] relu_9;
assign relu_9[7:0] = (bias_add_9[31]==0) ? ((bias_add_9<3'd6) ? {{bias_add_9[31],bias_add_9[10:4]}} :'d6) : '0;
logic [7:0] relu_10;
assign relu_10[7:0] = (bias_add_10[31]==0) ? ((bias_add_10<3'd6) ? {{bias_add_10[31],bias_add_10[10:4]}} :'d6) : '0;
logic [7:0] relu_11;
assign relu_11[7:0] = (bias_add_11[31]==0) ? ((bias_add_11<3'd6) ? {{bias_add_11[31],bias_add_11[10:4]}} :'d6) : '0;
logic [7:0] relu_12;
assign relu_12[7:0] = (bias_add_12[31]==0) ? ((bias_add_12<3'd6) ? {{bias_add_12[31],bias_add_12[10:4]}} :'d6) : '0;
logic [7:0] relu_13;
assign relu_13[7:0] = (bias_add_13[31]==0) ? ((bias_add_13<3'd6) ? {{bias_add_13[31],bias_add_13[10:4]}} :'d6) : '0;
logic [7:0] relu_14;
assign relu_14[7:0] = (bias_add_14[31]==0) ? ((bias_add_14<3'd6) ? {{bias_add_14[31],bias_add_14[10:4]}} :'d6) : '0;
logic [7:0] relu_15;
assign relu_15[7:0] = (bias_add_15[31]==0) ? ((bias_add_15<3'd6) ? {{bias_add_15[31],bias_add_15[10:4]}} :'d6) : '0;
logic [7:0] relu_16;
assign relu_16[7:0] = (bias_add_16[31]==0) ? ((bias_add_16<3'd6) ? {{bias_add_16[31],bias_add_16[10:4]}} :'d6) : '0;
logic [7:0] relu_17;
assign relu_17[7:0] = (bias_add_17[31]==0) ? ((bias_add_17<3'd6) ? {{bias_add_17[31],bias_add_17[10:4]}} :'d6) : '0;
logic [7:0] relu_18;
assign relu_18[7:0] = (bias_add_18[31]==0) ? ((bias_add_18<3'd6) ? {{bias_add_18[31],bias_add_18[10:4]}} :'d6) : '0;
logic [7:0] relu_19;
assign relu_19[7:0] = (bias_add_19[31]==0) ? ((bias_add_19<3'd6) ? {{bias_add_19[31],bias_add_19[10:4]}} :'d6) : '0;
logic [7:0] relu_20;
assign relu_20[7:0] = (bias_add_20[31]==0) ? ((bias_add_20<3'd6) ? {{bias_add_20[31],bias_add_20[10:4]}} :'d6) : '0;
logic [7:0] relu_21;
assign relu_21[7:0] = (bias_add_21[31]==0) ? ((bias_add_21<3'd6) ? {{bias_add_21[31],bias_add_21[10:4]}} :'d6) : '0;
logic [7:0] relu_22;
assign relu_22[7:0] = (bias_add_22[31]==0) ? ((bias_add_22<3'd6) ? {{bias_add_22[31],bias_add_22[10:4]}} :'d6) : '0;
logic [7:0] relu_23;
assign relu_23[7:0] = (bias_add_23[31]==0) ? ((bias_add_23<3'd6) ? {{bias_add_23[31],bias_add_23[10:4]}} :'d6) : '0;
logic [7:0] relu_24;
assign relu_24[7:0] = (bias_add_24[31]==0) ? ((bias_add_24<3'd6) ? {{bias_add_24[31],bias_add_24[10:4]}} :'d6) : '0;
logic [7:0] relu_25;
assign relu_25[7:0] = (bias_add_25[31]==0) ? ((bias_add_25<3'd6) ? {{bias_add_25[31],bias_add_25[10:4]}} :'d6) : '0;
logic [7:0] relu_26;
assign relu_26[7:0] = (bias_add_26[31]==0) ? ((bias_add_26<3'd6) ? {{bias_add_26[31],bias_add_26[10:4]}} :'d6) : '0;
logic [7:0] relu_27;
assign relu_27[7:0] = (bias_add_27[31]==0) ? ((bias_add_27<3'd6) ? {{bias_add_27[31],bias_add_27[10:4]}} :'d6) : '0;
logic [7:0] relu_28;
assign relu_28[7:0] = (bias_add_28[31]==0) ? ((bias_add_28<3'd6) ? {{bias_add_28[31],bias_add_28[10:4]}} :'d6) : '0;
logic [7:0] relu_29;
assign relu_29[7:0] = (bias_add_29[31]==0) ? ((bias_add_29<3'd6) ? {{bias_add_29[31],bias_add_29[10:4]}} :'d6) : '0;
logic [7:0] relu_30;
assign relu_30[7:0] = (bias_add_30[31]==0) ? ((bias_add_30<3'd6) ? {{bias_add_30[31],bias_add_30[10:4]}} :'d6) : '0;
logic [7:0] relu_31;
assign relu_31[7:0] = (bias_add_31[31]==0) ? ((bias_add_31<3'd6) ? {{bias_add_31[31],bias_add_31[10:4]}} :'d6) : '0;

assign output_act = {
	relu_31,
	relu_30,
	relu_29,
	relu_28,
	relu_27,
	relu_26,
	relu_25,
	relu_24,
	relu_23,
	relu_22,
	relu_21,
	relu_20,
	relu_19,
	relu_18,
	relu_17,
	relu_16,
	relu_15,
	relu_14,
	relu_13,
	relu_12,
	relu_11,
	relu_10,
	relu_9,
	relu_8,
	relu_7,
	relu_6,
	relu_5,
	relu_4,
	relu_3,
	relu_2,
	relu_1,
	relu_0
};

endmodule
module conv6_dw (
    input logic clk,
    input logic rstn,
    input logic valid,
    input logic [32*72-1:0] input_act,
    output logic [256-1:0] output_act,
    output logic ready
);
logic we;
logic [8:0] zero_number; 
assign zero_number = 9'd0; 
logic [32*72-1:0] input_act_ff;
genvar i;
generate
for (i=0;i<32;i++)
    begin: genblk_11
        always_ff @(posedge clk) begin
            if (rstn == 0) begin
                input_act_ff[(i+1)*72-1:i*72] <= '0;
            end
            else begin
                input_act_ff[(i+1)*72-1:i*72] <= input_act[(i+1)*72-1:i*72];
            end
        end
    end
endgenerate
logic [71:0] input_fmap_0;
assign input_fmap_0 = input_act_ff[71:0];
logic [71:0] input_fmap_1;
assign input_fmap_1 = input_act_ff[143:72];
logic [71:0] input_fmap_2;
assign input_fmap_2 = input_act_ff[215:144];
logic [71:0] input_fmap_3;
assign input_fmap_3 = input_act_ff[287:216];
logic [71:0] input_fmap_4;
assign input_fmap_4 = input_act_ff[359:288];
logic [71:0] input_fmap_5;
assign input_fmap_5 = input_act_ff[431:360];
logic [71:0] input_fmap_6;
assign input_fmap_6 = input_act_ff[503:432];
logic [71:0] input_fmap_7;
assign input_fmap_7 = input_act_ff[575:504];
logic [71:0] input_fmap_8;
assign input_fmap_8 = input_act_ff[647:576];
logic [71:0] input_fmap_9;
assign input_fmap_9 = input_act_ff[719:648];
logic [71:0] input_fmap_10;
assign input_fmap_10 = input_act_ff[791:720];
logic [71:0] input_fmap_11;
assign input_fmap_11 = input_act_ff[863:792];
logic [71:0] input_fmap_12;
assign input_fmap_12 = input_act_ff[935:864];
logic [71:0] input_fmap_13;
assign input_fmap_13 = input_act_ff[1007:936];
logic [71:0] input_fmap_14;
assign input_fmap_14 = input_act_ff[1079:1008];
logic [71:0] input_fmap_15;
assign input_fmap_15 = input_act_ff[1151:1080];
logic [71:0] input_fmap_16;
assign input_fmap_16 = input_act_ff[1223:1152];
logic [71:0] input_fmap_17;
assign input_fmap_17 = input_act_ff[1295:1224];
logic [71:0] input_fmap_18;
assign input_fmap_18 = input_act_ff[1367:1296];
logic [71:0] input_fmap_19;
assign input_fmap_19 = input_act_ff[1439:1368];
logic [71:0] input_fmap_20;
assign input_fmap_20 = input_act_ff[1511:1440];
logic [71:0] input_fmap_21;
assign input_fmap_21 = input_act_ff[1583:1512];
logic [71:0] input_fmap_22;
assign input_fmap_22 = input_act_ff[1655:1584];
logic [71:0] input_fmap_23;
assign input_fmap_23 = input_act_ff[1727:1656];
logic [71:0] input_fmap_24;
assign input_fmap_24 = input_act_ff[1799:1728];
logic [71:0] input_fmap_25;
assign input_fmap_25 = input_act_ff[1871:1800];
logic [71:0] input_fmap_26;
assign input_fmap_26 = input_act_ff[1943:1872];
logic [71:0] input_fmap_27;
assign input_fmap_27 = input_act_ff[2015:1944];
logic [71:0] input_fmap_28;
assign input_fmap_28 = input_act_ff[2087:2016];
logic [71:0] input_fmap_29;
assign input_fmap_29 = input_act_ff[2159:2088];
logic [71:0] input_fmap_30;
assign input_fmap_30 = input_act_ff[2231:2160];
logic [71:0] input_fmap_31;
assign input_fmap_31 = input_act_ff[2303:2232];

logic signed [31:0] conv_mac_0;
logic signed [63:0] chainout_0_O0; 
logic signed [63:0] O0_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O0(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd8),.bx(input_fmap_0[15:8]),.by(-9'sd7),.cx(input_fmap_0[23:16]),.cy(-9'sd4),.dx(input_fmap_0[31:24]),.dy(-9'sd11),.chainin(63'd0),.result(O0_N0_S1),.chainout(chainout_0_O0));
logic signed [63:0] chainout_2_O0; 
logic signed [63:0] O0_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O0(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[39:32]),.ay(-9'sd10),.bx(input_fmap_0[47:40]),.by(-9'sd6),.cx(input_fmap_0[55:48]),.cy(-9'sd5),.dx(input_fmap_0[63:56]),.dy(-9'sd5),.chainin(63'd0),.result(O0_N2_S1),.chainout(chainout_2_O0));
logic signed [63:0] chainout_4_O0; 
logic signed [63:0] O0_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O0(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[71:64]),.ay(-9'sd3),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O0_N4_S1),.chainout(chainout_4_O0));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O0_N0_S2;		always @(posedge clk) O0_N0_S2 <=     O0_N0_S1  +  O0_N2_S1 ;
 logic signed [21:0] O0_N2_S2;		always @(posedge clk) O0_N2_S2 <=     O0_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O0_N0_S3;		always @(posedge clk) O0_N0_S3 <=     O0_N0_S2  +  O0_N2_S2 ;
 assign conv_mac_0 = O0_N0_S3;

logic signed [31:0] conv_mac_1;
logic signed [63:0] chainout_0_O1; 
logic signed [63:0] O1_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O1(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay( 9'sd11),.bx(input_fmap_1[15:8]),.by( 9'sd10),.cx(input_fmap_1[23:16]),.cy( 9'sd2),.dx(input_fmap_1[31:24]),.dy( 9'sd18),.chainin(63'd0),.result(O1_N0_S1),.chainout(chainout_0_O1));
logic signed [63:0] chainout_2_O1; 
logic signed [63:0] O1_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O1(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[39:32]),.ay( 9'sd21),.bx(input_fmap_1[47:40]),.by( 9'sd4),.cx(input_fmap_1[55:48]),.cy( 9'sd10),.dx(input_fmap_1[63:56]),.dy( 9'sd10),.chainin(63'd0),.result(O1_N2_S1),.chainout(chainout_2_O1));
logic signed [63:0] chainout_4_O1; 
logic signed [63:0] O1_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O1(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[71:64]),.ay( 9'sd5),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O1_N4_S1),.chainout(chainout_4_O1));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O1_N0_S2;		always @(posedge clk) O1_N0_S2 <=     O1_N0_S1  +  O1_N2_S1 ;
 logic signed [21:0] O1_N2_S2;		always @(posedge clk) O1_N2_S2 <=     O1_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O1_N0_S3;		always @(posedge clk) O1_N0_S3 <=     O1_N0_S2  +  O1_N2_S2 ;
 assign conv_mac_1 = O1_N0_S3;

logic signed [31:0] conv_mac_2;
logic signed [63:0] chainout_0_O2; 
logic signed [63:0] O2_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O2(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_2[7:0]),.ay( 9'sd11),.bx(input_fmap_2[15:8]),.by( 9'sd11),.cx(input_fmap_2[23:16]),.cy( 9'sd5),.dx(input_fmap_2[31:24]),.dy( 9'sd12),.chainin(63'd0),.result(O2_N0_S1),.chainout(chainout_0_O2));
logic signed [63:0] chainout_2_O2; 
logic signed [63:0] O2_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O2(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_2[39:32]),.ay( 9'sd14),.bx(input_fmap_2[47:40]),.by( 9'sd7),.cx(input_fmap_2[55:48]),.cy( 9'sd7),.dx(input_fmap_2[63:56]),.dy( 9'sd5),.chainin(63'd0),.result(O2_N2_S1),.chainout(chainout_2_O2));
logic signed [63:0] chainout_4_O2; 
logic signed [63:0] O2_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O2(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_2[71:64]),.ay( 9'sd5),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O2_N4_S1),.chainout(chainout_4_O2));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O2_N0_S2;		always @(posedge clk) O2_N0_S2 <=     O2_N0_S1  +  O2_N2_S1 ;
 logic signed [21:0] O2_N2_S2;		always @(posedge clk) O2_N2_S2 <=     O2_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O2_N0_S3;		always @(posedge clk) O2_N0_S3 <=     O2_N0_S2  +  O2_N2_S2 ;
 assign conv_mac_2 = O2_N0_S3;

logic signed [31:0] conv_mac_3;
logic signed [63:0] chainout_0_O3; 
logic signed [63:0] O3_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O3(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_3[7:0]),.ay( 9'sd10),.bx(input_fmap_3[15:8]),.by( 9'sd11),.cx(input_fmap_3[23:16]),.cy( 9'sd7),.dx(input_fmap_3[31:24]),.dy( 9'sd9),.chainin(63'd0),.result(O3_N0_S1),.chainout(chainout_0_O3));
logic signed [63:0] chainout_2_O3; 
logic signed [63:0] O3_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O3(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_3[39:32]),.ay( 9'sd13),.bx(input_fmap_3[47:40]),.by( 9'sd7),.cx(input_fmap_3[55:48]),.cy( 9'sd4),.dx(input_fmap_3[63:56]),.dy( 9'sd7),.chainin(63'd0),.result(O3_N2_S1),.chainout(chainout_2_O3));
logic signed [63:0] chainout_4_O3; 
logic signed [63:0] O3_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O3(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_3[71:64]),.ay( 9'sd3),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O3_N4_S1),.chainout(chainout_4_O3));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O3_N0_S2;		always @(posedge clk) O3_N0_S2 <=     O3_N0_S1  +  O3_N2_S1 ;
 logic signed [21:0] O3_N2_S2;		always @(posedge clk) O3_N2_S2 <=     O3_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O3_N0_S3;		always @(posedge clk) O3_N0_S3 <=     O3_N0_S2  +  O3_N2_S2 ;
 assign conv_mac_3 = O3_N0_S3;

logic signed [31:0] conv_mac_4;
logic signed [63:0] chainout_0_O4; 
logic signed [63:0] O4_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O4(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_4[7:0]),.ay( 9'sd10),.bx(input_fmap_4[15:8]),.by(-9'sd1),.cx(input_fmap_4[23:16]),.cy(-9'sd6),.dx(input_fmap_4[31:24]),.dy( 9'sd14),.chainin(63'd0),.result(O4_N0_S1),.chainout(chainout_0_O4));
logic signed [63:0] chainout_2_O4; 
logic signed [63:0] O4_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O4(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_4[39:32]),.ay(-9'sd5),.bx(input_fmap_4[47:40]),.by(-9'sd9),.cx(input_fmap_4[55:48]),.cy( 9'sd7),.dx(input_fmap_4[63:56]),.dy(-9'sd3),.chainin(63'd0),.result(O4_N2_S1),.chainout(chainout_2_O4));
logic signed [63:0] chainout_4_O4; 
logic signed [63:0] O4_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O4(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_4[71:64]),.ay(-9'sd6),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O4_N4_S1),.chainout(chainout_4_O4));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O4_N0_S2;		always @(posedge clk) O4_N0_S2 <=     O4_N0_S1  +  O4_N2_S1 ;
 logic signed [21:0] O4_N2_S2;		always @(posedge clk) O4_N2_S2 <=     O4_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O4_N0_S3;		always @(posedge clk) O4_N0_S3 <=     O4_N0_S2  +  O4_N2_S2 ;
 assign conv_mac_4 = O4_N0_S3;

logic signed [31:0] conv_mac_5;
logic signed [63:0] chainout_0_O5; 
logic signed [63:0] O5_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O5(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_5[7:0]),.ay( 9'sd6),.bx(input_fmap_5[15:8]),.by( 9'sd10),.cx(input_fmap_5[23:16]),.cy( 9'sd3),.dx(input_fmap_5[31:24]),.dy( 9'sd9),.chainin(63'd0),.result(O5_N0_S1),.chainout(chainout_0_O5));
logic signed [63:0] chainout_2_O5; 
logic signed [63:0] O5_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O5(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_5[39:32]),.ay( 9'sd12),.bx(input_fmap_5[47:40]),.by( 9'sd7),.cx(input_fmap_5[55:48]),.cy( 9'sd3),.dx(input_fmap_5[63:56]),.dy( 9'sd4),.chainin(63'd0),.result(O5_N2_S1),.chainout(chainout_2_O5));
logic signed [63:0] chainout_4_O5; 
logic signed [63:0] O5_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O5(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_5[71:64]),.ay( 9'sd6),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O5_N4_S1),.chainout(chainout_4_O5));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O5_N0_S2;		always @(posedge clk) O5_N0_S2 <=     O5_N0_S1  +  O5_N2_S1 ;
 logic signed [21:0] O5_N2_S2;		always @(posedge clk) O5_N2_S2 <=     O5_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O5_N0_S3;		always @(posedge clk) O5_N0_S3 <=     O5_N0_S2  +  O5_N2_S2 ;
 assign conv_mac_5 = O5_N0_S3;

logic signed [31:0] conv_mac_6;
logic signed [63:0] chainout_0_O6; 
logic signed [63:0] O6_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O6(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_6[7:0]),.ay( 9'sd7),.bx(input_fmap_6[15:8]),.by( 9'sd11),.cx(input_fmap_6[23:16]),.cy( 9'sd7),.dx(input_fmap_6[31:24]),.dy( 9'sd7),.chainin(63'd0),.result(O6_N0_S1),.chainout(chainout_0_O6));
logic signed [63:0] chainout_2_O6; 
logic signed [63:0] O6_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O6(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_6[39:32]),.ay( 9'sd14),.bx(input_fmap_6[47:40]),.by( 9'sd11),.cx(input_fmap_6[55:48]),.cy( 9'sd3),.dx(input_fmap_6[63:56]),.dy( 9'sd7),.chainin(63'd0),.result(O6_N2_S1),.chainout(chainout_2_O6));
logic signed [63:0] chainout_4_O6; 
logic signed [63:0] O6_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O6(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_6[71:64]),.ay( 9'sd7),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O6_N4_S1),.chainout(chainout_4_O6));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O6_N0_S2;		always @(posedge clk) O6_N0_S2 <=     O6_N0_S1  +  O6_N2_S1 ;
 logic signed [21:0] O6_N2_S2;		always @(posedge clk) O6_N2_S2 <=     O6_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O6_N0_S3;		always @(posedge clk) O6_N0_S3 <=     O6_N0_S2  +  O6_N2_S2 ;
 assign conv_mac_6 = O6_N0_S3;

logic signed [31:0] conv_mac_7;
logic signed [63:0] chainout_0_O7; 
logic signed [63:0] O7_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O7(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_7[7:0]),.ay( 9'sd9),.bx(input_fmap_7[15:8]),.by( 9'sd11),.cx(input_fmap_7[23:16]),.cy( 9'sd4),.dx(input_fmap_7[31:24]),.dy( 9'sd13),.chainin(63'd0),.result(O7_N0_S1),.chainout(chainout_0_O7));
logic signed [63:0] chainout_2_O7; 
logic signed [63:0] O7_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O7(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_7[39:32]),.ay( 9'sd16),.bx(input_fmap_7[47:40]),.by( 9'sd9),.cx(input_fmap_7[55:48]),.cy( 9'sd5),.dx(input_fmap_7[63:56]),.dy( 9'sd10),.chainin(63'd0),.result(O7_N2_S1),.chainout(chainout_2_O7));
logic signed [63:0] chainout_4_O7; 
logic signed [63:0] O7_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O7(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_7[71:64]),.ay( 9'sd6),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O7_N4_S1),.chainout(chainout_4_O7));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O7_N0_S2;		always @(posedge clk) O7_N0_S2 <=     O7_N0_S1  +  O7_N2_S1 ;
 logic signed [21:0] O7_N2_S2;		always @(posedge clk) O7_N2_S2 <=     O7_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O7_N0_S3;		always @(posedge clk) O7_N0_S3 <=     O7_N0_S2  +  O7_N2_S2 ;
 assign conv_mac_7 = O7_N0_S3;

logic signed [31:0] conv_mac_8;
logic signed [63:0] chainout_0_O8; 
logic signed [63:0] O8_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O8(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_8[7:0]),.ay(-9'sd10),.bx(input_fmap_8[15:8]),.by( 9'sd7),.cx(input_fmap_8[23:16]),.cy( 9'sd5),.dx(input_fmap_8[31:24]),.dy(-9'sd14),.chainin(63'd0),.result(O8_N0_S1),.chainout(chainout_0_O8));
logic signed [63:0] chainout_2_O8; 
logic signed [63:0] O8_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O8(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_8[39:32]),.ay( 9'sd4),.bx(input_fmap_8[47:40]),.by( 9'sd8),.cx(input_fmap_8[55:48]),.cy(-9'sd10),.dx(input_fmap_8[63:56]),.dy(-9'sd1),.chainin(63'd0),.result(O8_N2_S1),.chainout(chainout_2_O8));
logic signed [63:0] chainout_4_O8; 
logic signed [63:0] O8_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O8(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_8[71:64]),.ay( 9'sd6),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O8_N4_S1),.chainout(chainout_4_O8));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O8_N0_S2;		always @(posedge clk) O8_N0_S2 <=     O8_N0_S1  +  O8_N2_S1 ;
 logic signed [21:0] O8_N2_S2;		always @(posedge clk) O8_N2_S2 <=     O8_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O8_N0_S3;		always @(posedge clk) O8_N0_S3 <=     O8_N0_S2  +  O8_N2_S2 ;
 assign conv_mac_8 = O8_N0_S3;

logic signed [31:0] conv_mac_9;
logic signed [63:0] chainout_0_O9; 
logic signed [63:0] O9_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O9(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_9[7:0]),.ay(-9'sd3),.bx(input_fmap_9[15:8]),.by( 9'sd12),.cx(input_fmap_9[23:16]),.cy( 9'sd8),.dx(input_fmap_9[31:24]),.dy( 9'sd2),.chainin(63'd0),.result(O9_N0_S1),.chainout(chainout_0_O9));
logic signed [63:0] chainout_2_O9; 
logic signed [63:0] O9_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O9(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_9[39:32]),.ay( 9'sd13),.bx(input_fmap_9[47:40]),.by( 9'sd13),.cx(input_fmap_9[55:48]),.cy( 9'sd3),.dx(input_fmap_9[63:56]),.dy( 9'sd7),.chainin(63'd0),.result(O9_N2_S1),.chainout(chainout_2_O9));
logic signed [63:0] chainout_4_O9; 
logic signed [63:0] O9_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O9(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_9[71:64]),.ay( 9'sd7),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O9_N4_S1),.chainout(chainout_4_O9));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O9_N0_S2;		always @(posedge clk) O9_N0_S2 <=     O9_N0_S1  +  O9_N2_S1 ;
 logic signed [21:0] O9_N2_S2;		always @(posedge clk) O9_N2_S2 <=     O9_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O9_N0_S3;		always @(posedge clk) O9_N0_S3 <=     O9_N0_S2  +  O9_N2_S2 ;
 assign conv_mac_9 = O9_N0_S3;

logic signed [31:0] conv_mac_10;
logic signed [63:0] chainout_0_O10; 
logic signed [63:0] O10_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O10(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_10[7:0]),.ay( 9'sd5),.bx(input_fmap_10[15:8]),.by( 9'sd11),.cx(input_fmap_10[23:16]),.cy( 9'sd8),.dx(input_fmap_10[31:24]),.dy( 9'sd9),.chainin(63'd0),.result(O10_N0_S1),.chainout(chainout_0_O10));
logic signed [63:0] chainout_2_O10; 
logic signed [63:0] O10_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O10(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_10[39:32]),.ay( 9'sd19),.bx(input_fmap_10[47:40]),.by( 9'sd9),.cx(input_fmap_10[55:48]),.cy( 9'sd4),.dx(input_fmap_10[63:56]),.dy( 9'sd8),.chainin(63'd0),.result(O10_N2_S1),.chainout(chainout_2_O10));
logic signed [63:0] chainout_4_O10; 
logic signed [63:0] O10_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O10(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_10[71:64]),.ay( 9'sd4),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O10_N4_S1),.chainout(chainout_4_O10));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O10_N0_S2;		always @(posedge clk) O10_N0_S2 <=     O10_N0_S1  +  O10_N2_S1 ;
 logic signed [21:0] O10_N2_S2;		always @(posedge clk) O10_N2_S2 <=     O10_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O10_N0_S3;		always @(posedge clk) O10_N0_S3 <=     O10_N0_S2  +  O10_N2_S2 ;
 assign conv_mac_10 = O10_N0_S3;

logic signed [31:0] conv_mac_11;
logic signed [63:0] chainout_0_O11; 
logic signed [63:0] O11_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O11(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_11[7:0]),.ay( 9'sd8),.bx(input_fmap_11[15:8]),.by( 9'sd11),.cx(input_fmap_11[23:16]),.cy( 9'sd6),.dx(input_fmap_11[31:24]),.dy( 9'sd10),.chainin(63'd0),.result(O11_N0_S1),.chainout(chainout_0_O11));
logic signed [63:0] chainout_2_O11; 
logic signed [63:0] O11_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O11(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_11[39:32]),.ay( 9'sd12),.bx(input_fmap_11[47:40]),.by( 9'sd8),.cx(input_fmap_11[55:48]),.cy( 9'sd6),.dx(input_fmap_11[63:56]),.dy( 9'sd4),.chainin(63'd0),.result(O11_N2_S1),.chainout(chainout_2_O11));
logic signed [63:0] chainout_4_O11; 
logic signed [63:0] O11_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O11(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_11[71:64]),.ay( 9'sd2),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O11_N4_S1),.chainout(chainout_4_O11));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O11_N0_S2;		always @(posedge clk) O11_N0_S2 <=     O11_N0_S1  +  O11_N2_S1 ;
 logic signed [21:0] O11_N2_S2;		always @(posedge clk) O11_N2_S2 <=     O11_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O11_N0_S3;		always @(posedge clk) O11_N0_S3 <=     O11_N0_S2  +  O11_N2_S2 ;
 assign conv_mac_11 = O11_N0_S3;

logic signed [31:0] conv_mac_12;
logic signed [63:0] chainout_0_O12; 
logic signed [63:0] O12_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O12(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_12[15:8]),.ay( 9'sd4),.bx(input_fmap_12[23:16]),.by( 9'sd5),.cx(input_fmap_12[31:24]),.cy( 9'sd4),.dx(input_fmap_12[39:32]),.dy( 9'sd9),.chainin(63'd0),.result(O12_N0_S1),.chainout(chainout_0_O12));
logic signed [63:0] chainout_2_O12; 
logic signed [63:0] O12_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O12(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_12[47:40]),.ay( 9'sd10),.bx(input_fmap_12[55:48]),.by( 9'sd4),.cx(input_fmap_12[63:56]),.cy( 9'sd10),.dx(input_fmap_12[71:64]),.dy( 9'sd8),.chainin(63'd0),.result(O12_N2_S1),.chainout(chainout_2_O12));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O12_N0_S2;		always @(posedge clk) O12_N0_S2 <=     O12_N0_S1  +  O12_N2_S1 ;
 assign conv_mac_12 = O12_N0_S2;

logic signed [31:0] conv_mac_13;
logic signed [63:0] chainout_0_O13; 
logic signed [63:0] O13_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O13(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_13[7:0]),.ay( 9'sd9),.bx(input_fmap_13[15:8]),.by( 9'sd9),.cx(input_fmap_13[23:16]),.cy( 9'sd5),.dx(input_fmap_13[31:24]),.dy( 9'sd11),.chainin(63'd0),.result(O13_N0_S1),.chainout(chainout_0_O13));
logic signed [63:0] chainout_2_O13; 
logic signed [63:0] O13_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O13(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_13[39:32]),.ay( 9'sd17),.bx(input_fmap_13[47:40]),.by( 9'sd6),.cx(input_fmap_13[55:48]),.cy( 9'sd6),.dx(input_fmap_13[63:56]),.dy( 9'sd8),.chainin(63'd0),.result(O13_N2_S1),.chainout(chainout_2_O13));
logic signed [63:0] chainout_4_O13; 
logic signed [63:0] O13_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O13(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_13[71:64]),.ay( 9'sd7),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O13_N4_S1),.chainout(chainout_4_O13));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O13_N0_S2;		always @(posedge clk) O13_N0_S2 <=     O13_N0_S1  +  O13_N2_S1 ;
 logic signed [21:0] O13_N2_S2;		always @(posedge clk) O13_N2_S2 <=     O13_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O13_N0_S3;		always @(posedge clk) O13_N0_S3 <=     O13_N0_S2  +  O13_N2_S2 ;
 assign conv_mac_13 = O13_N0_S3;

logic signed [31:0] conv_mac_14;
logic signed [63:0] chainout_0_O14; 
logic signed [63:0] O14_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O14(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_14[7:0]),.ay(-9'sd2),.bx(input_fmap_14[15:8]),.by(-9'sd7),.cx(input_fmap_14[23:16]),.cy(-9'sd7),.dx(input_fmap_14[31:24]),.dy(-9'sd5),.chainin(63'd0),.result(O14_N0_S1),.chainout(chainout_0_O14));
logic signed [63:0] chainout_2_O14; 
logic signed [63:0] O14_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O14(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_14[39:32]),.ay(-9'sd11),.bx(input_fmap_14[47:40]),.by(-9'sd11),.cx(input_fmap_14[55:48]),.cy(-9'sd4),.dx(input_fmap_14[63:56]),.dy(-9'sd8),.chainin(63'd0),.result(O14_N2_S1),.chainout(chainout_2_O14));
logic signed [63:0] chainout_4_O14; 
logic signed [63:0] O14_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O14(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_14[71:64]),.ay(-9'sd8),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O14_N4_S1),.chainout(chainout_4_O14));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O14_N0_S2;		always @(posedge clk) O14_N0_S2 <=     O14_N0_S1  +  O14_N2_S1 ;
 logic signed [21:0] O14_N2_S2;		always @(posedge clk) O14_N2_S2 <=     O14_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O14_N0_S3;		always @(posedge clk) O14_N0_S3 <=     O14_N0_S2  +  O14_N2_S2 ;
 assign conv_mac_14 = O14_N0_S3;

logic signed [31:0] conv_mac_15;
logic signed [63:0] chainout_0_O15; 
logic signed [63:0] O15_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O15(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_15[7:0]),.ay(-9'sd6),.bx(input_fmap_15[15:8]),.by(-9'sd7),.cx(input_fmap_15[23:16]),.cy(-9'sd3),.dx(input_fmap_15[31:24]),.dy(-9'sd8),.chainin(63'd0),.result(O15_N0_S1),.chainout(chainout_0_O15));
logic signed [63:0] chainout_2_O15; 
logic signed [63:0] O15_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O15(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_15[39:32]),.ay(-9'sd11),.bx(input_fmap_15[47:40]),.by(-9'sd6),.cx(input_fmap_15[55:48]),.cy(-9'sd4),.dx(input_fmap_15[63:56]),.dy(-9'sd5),.chainin(63'd0),.result(O15_N2_S1),.chainout(chainout_2_O15));
logic signed [63:0] chainout_4_O15; 
logic signed [63:0] O15_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O15(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_15[71:64]),.ay(-9'sd4),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O15_N4_S1),.chainout(chainout_4_O15));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O15_N0_S2;		always @(posedge clk) O15_N0_S2 <=     O15_N0_S1  +  O15_N2_S1 ;
 logic signed [21:0] O15_N2_S2;		always @(posedge clk) O15_N2_S2 <=     O15_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O15_N0_S3;		always @(posedge clk) O15_N0_S3 <=     O15_N0_S2  +  O15_N2_S2 ;
 assign conv_mac_15 = O15_N0_S3;

logic signed [31:0] conv_mac_16;
logic signed [63:0] chainout_0_O16; 
logic signed [63:0] O16_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O16(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_16[7:0]),.ay( 9'sd7),.bx(input_fmap_16[15:8]),.by( 9'sd8),.cx(input_fmap_16[23:16]),.cy( 9'sd4),.dx(input_fmap_16[31:24]),.dy( 9'sd8),.chainin(63'd0),.result(O16_N0_S1),.chainout(chainout_0_O16));
logic signed [63:0] chainout_2_O16; 
logic signed [63:0] O16_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O16(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_16[39:32]),.ay( 9'sd13),.bx(input_fmap_16[47:40]),.by( 9'sd8),.cx(input_fmap_16[55:48]),.cy( 9'sd5),.dx(input_fmap_16[63:56]),.dy( 9'sd6),.chainin(63'd0),.result(O16_N2_S1),.chainout(chainout_2_O16));
logic signed [63:0] chainout_4_O16; 
logic signed [63:0] O16_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O16(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_16[71:64]),.ay( 9'sd4),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O16_N4_S1),.chainout(chainout_4_O16));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O16_N0_S2;		always @(posedge clk) O16_N0_S2 <=     O16_N0_S1  +  O16_N2_S1 ;
 logic signed [21:0] O16_N2_S2;		always @(posedge clk) O16_N2_S2 <=     O16_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O16_N0_S3;		always @(posedge clk) O16_N0_S3 <=     O16_N0_S2  +  O16_N2_S2 ;
 assign conv_mac_16 = O16_N0_S3;

logic signed [31:0] conv_mac_17;
logic signed [63:0] chainout_0_O17; 
logic signed [63:0] O17_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O17(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_17[7:0]),.ay( 9'sd10),.bx(input_fmap_17[15:8]),.by( 9'sd11),.cx(input_fmap_17[23:16]),.cy( 9'sd5),.dx(input_fmap_17[31:24]),.dy( 9'sd12),.chainin(63'd0),.result(O17_N0_S1),.chainout(chainout_0_O17));
logic signed [63:0] chainout_2_O17; 
logic signed [63:0] O17_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O17(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_17[39:32]),.ay( 9'sd14),.bx(input_fmap_17[47:40]),.by( 9'sd4),.cx(input_fmap_17[55:48]),.cy( 9'sd8),.dx(input_fmap_17[63:56]),.dy( 9'sd7),.chainin(63'd0),.result(O17_N2_S1),.chainout(chainout_2_O17));
logic signed [63:0] chainout_4_O17; 
logic signed [63:0] O17_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O17(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_17[71:64]),.ay( 9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O17_N4_S1),.chainout(chainout_4_O17));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O17_N0_S2;		always @(posedge clk) O17_N0_S2 <=     O17_N0_S1  +  O17_N2_S1 ;
 logic signed [21:0] O17_N2_S2;		always @(posedge clk) O17_N2_S2 <=     O17_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O17_N0_S3;		always @(posedge clk) O17_N0_S3 <=     O17_N0_S2  +  O17_N2_S2 ;
 assign conv_mac_17 = O17_N0_S3;

logic signed [31:0] conv_mac_18;
logic signed [63:0] chainout_0_O18; 
logic signed [63:0] O18_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O18(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_18[7:0]),.ay(-9'sd5),.bx(input_fmap_18[15:8]),.by(-9'sd10),.cx(input_fmap_18[23:16]),.cy(-9'sd5),.dx(input_fmap_18[31:24]),.dy(-9'sd9),.chainin(63'd0),.result(O18_N0_S1),.chainout(chainout_0_O18));
logic signed [63:0] chainout_2_O18; 
logic signed [63:0] O18_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O18(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_18[39:32]),.ay(-9'sd13),.bx(input_fmap_18[47:40]),.by(-9'sd5),.cx(input_fmap_18[55:48]),.cy(-9'sd4),.dx(input_fmap_18[63:56]),.dy(-9'sd6),.chainin(63'd0),.result(O18_N2_S1),.chainout(chainout_2_O18));
logic signed [63:0] chainout_4_O18; 
logic signed [63:0] O18_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O18(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_18[71:64]),.ay(-9'sd4),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O18_N4_S1),.chainout(chainout_4_O18));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O18_N0_S2;		always @(posedge clk) O18_N0_S2 <=     O18_N0_S1  +  O18_N2_S1 ;
 logic signed [21:0] O18_N2_S2;		always @(posedge clk) O18_N2_S2 <=     O18_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O18_N0_S3;		always @(posedge clk) O18_N0_S3 <=     O18_N0_S2  +  O18_N2_S2 ;
 assign conv_mac_18 = O18_N0_S3;

logic signed [31:0] conv_mac_19;
logic signed [63:0] chainout_0_O19; 
logic signed [63:0] O19_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O19(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_19[7:0]),.ay(-9'sd8),.bx(input_fmap_19[15:8]),.by(-9'sd9),.cx(input_fmap_19[23:16]),.cy(-9'sd5),.dx(input_fmap_19[31:24]),.dy(-9'sd11),.chainin(63'd0),.result(O19_N0_S1),.chainout(chainout_0_O19));
logic signed [63:0] chainout_2_O19; 
logic signed [63:0] O19_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O19(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_19[39:32]),.ay(-9'sd11),.bx(input_fmap_19[55:48]),.by(-9'sd6),.cx(input_fmap_19[63:56]),.cy(-9'sd1),.dx(input_fmap_19[71:64]),.dy(-9'sd3),.chainin(63'd0),.result(O19_N2_S1),.chainout(chainout_2_O19));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O19_N0_S2;		always @(posedge clk) O19_N0_S2 <=     O19_N0_S1  +  O19_N2_S1 ;
 assign conv_mac_19 = O19_N0_S2;

logic signed [31:0] conv_mac_20;
logic signed [63:0] chainout_0_O20; 
logic signed [63:0] O20_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O20(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_20[7:0]),.ay(-9'sd10),.bx(input_fmap_20[15:8]),.by(-9'sd11),.cx(input_fmap_20[23:16]),.cy(-9'sd3),.dx(input_fmap_20[31:24]),.dy(-9'sd9),.chainin(63'd0),.result(O20_N0_S1),.chainout(chainout_0_O20));
logic signed [63:0] chainout_2_O20; 
logic signed [63:0] O20_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O20(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_20[39:32]),.ay(-9'sd12),.bx(input_fmap_20[47:40]),.by(-9'sd4),.cx(input_fmap_20[55:48]),.cy(-9'sd5),.dx(input_fmap_20[63:56]),.dy(-9'sd4),.chainin(63'd0),.result(O20_N2_S1),.chainout(chainout_2_O20));
logic signed [63:0] chainout_4_O20; 
logic signed [63:0] O20_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O20(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_20[71:64]),.ay(-9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O20_N4_S1),.chainout(chainout_4_O20));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O20_N0_S2;		always @(posedge clk) O20_N0_S2 <=     O20_N0_S1  +  O20_N2_S1 ;
 logic signed [21:0] O20_N2_S2;		always @(posedge clk) O20_N2_S2 <=     O20_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O20_N0_S3;		always @(posedge clk) O20_N0_S3 <=     O20_N0_S2  +  O20_N2_S2 ;
 assign conv_mac_20 = O20_N0_S3;

logic signed [31:0] conv_mac_21;
logic signed [63:0] chainout_0_O21; 
logic signed [63:0] O21_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O21(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_21[7:0]),.ay(-9'sd6),.bx(input_fmap_21[15:8]),.by(-9'sd7),.cx(input_fmap_21[23:16]),.cy(-9'sd4),.dx(input_fmap_21[31:24]),.dy(-9'sd8),.chainin(63'd0),.result(O21_N0_S1),.chainout(chainout_0_O21));
logic signed [63:0] chainout_2_O21; 
logic signed [63:0] O21_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O21(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_21[39:32]),.ay(-9'sd13),.bx(input_fmap_21[47:40]),.by(-9'sd6),.cx(input_fmap_21[55:48]),.cy(-9'sd3),.dx(input_fmap_21[63:56]),.dy(-9'sd7),.chainin(63'd0),.result(O21_N2_S1),.chainout(chainout_2_O21));
logic signed [63:0] chainout_4_O21; 
logic signed [63:0] O21_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O21(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_21[71:64]),.ay(-9'sd2),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O21_N4_S1),.chainout(chainout_4_O21));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O21_N0_S2;		always @(posedge clk) O21_N0_S2 <=     O21_N0_S1  +  O21_N2_S1 ;
 logic signed [21:0] O21_N2_S2;		always @(posedge clk) O21_N2_S2 <=     O21_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O21_N0_S3;		always @(posedge clk) O21_N0_S3 <=     O21_N0_S2  +  O21_N2_S2 ;
 assign conv_mac_21 = O21_N0_S3;

logic signed [31:0] conv_mac_22;
logic signed [63:0] chainout_0_O22; 
logic signed [63:0] O22_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O22(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_22[7:0]),.ay(-9'sd6),.bx(input_fmap_22[15:8]),.by(-9'sd7),.cx(input_fmap_22[23:16]),.cy(-9'sd4),.dx(input_fmap_22[31:24]),.dy(-9'sd10),.chainin(63'd0),.result(O22_N0_S1),.chainout(chainout_0_O22));
logic signed [63:0] chainout_2_O22; 
logic signed [63:0] O22_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O22(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_22[39:32]),.ay(-9'sd11),.bx(input_fmap_22[47:40]),.by(-9'sd5),.cx(input_fmap_22[55:48]),.cy(-9'sd4),.dx(input_fmap_22[63:56]),.dy(-9'sd5),.chainin(63'd0),.result(O22_N2_S1),.chainout(chainout_2_O22));
logic signed [63:0] chainout_4_O22; 
logic signed [63:0] O22_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O22(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_22[71:64]),.ay(-9'sd3),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O22_N4_S1),.chainout(chainout_4_O22));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O22_N0_S2;		always @(posedge clk) O22_N0_S2 <=     O22_N0_S1  +  O22_N2_S1 ;
 logic signed [21:0] O22_N2_S2;		always @(posedge clk) O22_N2_S2 <=     O22_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O22_N0_S3;		always @(posedge clk) O22_N0_S3 <=     O22_N0_S2  +  O22_N2_S2 ;
 assign conv_mac_22 = O22_N0_S3;

logic signed [31:0] conv_mac_23;
logic signed [63:0] chainout_0_O23; 
logic signed [63:0] O23_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O23(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_23[7:0]),.ay( 9'sd11),.bx(input_fmap_23[15:8]),.by( 9'sd11),.cx(input_fmap_23[23:16]),.cy( 9'sd6),.dx(input_fmap_23[31:24]),.dy( 9'sd13),.chainin(63'd0),.result(O23_N0_S1),.chainout(chainout_0_O23));
logic signed [63:0] chainout_2_O23; 
logic signed [63:0] O23_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O23(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_23[39:32]),.ay( 9'sd20),.bx(input_fmap_23[47:40]),.by( 9'sd9),.cx(input_fmap_23[55:48]),.cy( 9'sd6),.dx(input_fmap_23[63:56]),.dy( 9'sd8),.chainin(63'd0),.result(O23_N2_S1),.chainout(chainout_2_O23));
logic signed [63:0] chainout_4_O23; 
logic signed [63:0] O23_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O23(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_23[71:64]),.ay( 9'sd6),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O23_N4_S1),.chainout(chainout_4_O23));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O23_N0_S2;		always @(posedge clk) O23_N0_S2 <=     O23_N0_S1  +  O23_N2_S1 ;
 logic signed [21:0] O23_N2_S2;		always @(posedge clk) O23_N2_S2 <=     O23_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O23_N0_S3;		always @(posedge clk) O23_N0_S3 <=     O23_N0_S2  +  O23_N2_S2 ;
 assign conv_mac_23 = O23_N0_S3;

logic signed [31:0] conv_mac_24;
logic signed [63:0] chainout_0_O24; 
logic signed [63:0] O24_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O24(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_24[7:0]),.ay(-9'sd4),.bx(input_fmap_24[15:8]),.by(-9'sd10),.cx(input_fmap_24[23:16]),.cy(-9'sd6),.dx(input_fmap_24[31:24]),.dy(-9'sd7),.chainin(63'd0),.result(O24_N0_S1),.chainout(chainout_0_O24));
logic signed [63:0] chainout_2_O24; 
logic signed [63:0] O24_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O24(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_24[39:32]),.ay(-9'sd11),.bx(input_fmap_24[47:40]),.by(-9'sd8),.cx(input_fmap_24[55:48]),.cy(-9'sd2),.dx(input_fmap_24[63:56]),.dy(-9'sd5),.chainin(63'd0),.result(O24_N2_S1),.chainout(chainout_2_O24));
logic signed [63:0] chainout_4_O24; 
logic signed [63:0] O24_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O24(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_24[71:64]),.ay(-9'sd4),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O24_N4_S1),.chainout(chainout_4_O24));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O24_N0_S2;		always @(posedge clk) O24_N0_S2 <=     O24_N0_S1  +  O24_N2_S1 ;
 logic signed [21:0] O24_N2_S2;		always @(posedge clk) O24_N2_S2 <=     O24_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O24_N0_S3;		always @(posedge clk) O24_N0_S3 <=     O24_N0_S2  +  O24_N2_S2 ;
 assign conv_mac_24 = O24_N0_S3;

logic signed [31:0] conv_mac_25;
logic signed [63:0] chainout_0_O25; 
logic signed [63:0] O25_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O25(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_25[7:0]),.ay(-9'sd10),.bx(input_fmap_25[15:8]),.by(-9'sd14),.cx(input_fmap_25[23:16]),.cy(-9'sd4),.dx(input_fmap_25[31:24]),.dy(-9'sd12),.chainin(63'd0),.result(O25_N0_S1),.chainout(chainout_0_O25));
logic signed [63:0] chainout_2_O25; 
logic signed [63:0] O25_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O25(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_25[39:32]),.ay(-9'sd15),.bx(input_fmap_25[47:40]),.by(-9'sd6),.cx(input_fmap_25[55:48]),.cy(-9'sd3),.dx(input_fmap_25[63:56]),.dy(-9'sd6),.chainin(63'd0),.result(O25_N2_S1),.chainout(chainout_2_O25));
logic signed [63:0] chainout_4_O25; 
logic signed [63:0] O25_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O25(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_25[71:64]),.ay(-9'sd4),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O25_N4_S1),.chainout(chainout_4_O25));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O25_N0_S2;		always @(posedge clk) O25_N0_S2 <=     O25_N0_S1  +  O25_N2_S1 ;
 logic signed [21:0] O25_N2_S2;		always @(posedge clk) O25_N2_S2 <=     O25_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O25_N0_S3;		always @(posedge clk) O25_N0_S3 <=     O25_N0_S2  +  O25_N2_S2 ;
 assign conv_mac_25 = O25_N0_S3;

logic signed [31:0] conv_mac_26;
logic signed [63:0] chainout_0_O26; 
logic signed [63:0] O26_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O26(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_26[7:0]),.ay( 9'sd8),.bx(input_fmap_26[15:8]),.by( 9'sd13),.cx(input_fmap_26[23:16]),.cy( 9'sd6),.dx(input_fmap_26[31:24]),.dy( 9'sd10),.chainin(63'd0),.result(O26_N0_S1),.chainout(chainout_0_O26));
logic signed [63:0] chainout_2_O26; 
logic signed [63:0] O26_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O26(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_26[39:32]),.ay( 9'sd17),.bx(input_fmap_26[47:40]),.by( 9'sd5),.cx(input_fmap_26[55:48]),.cy( 9'sd3),.dx(input_fmap_26[63:56]),.dy( 9'sd9),.chainin(63'd0),.result(O26_N2_S1),.chainout(chainout_2_O26));
logic signed [63:0] chainout_4_O26; 
logic signed [63:0] O26_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O26(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_26[71:64]),.ay( 9'sd4),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O26_N4_S1),.chainout(chainout_4_O26));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O26_N0_S2;		always @(posedge clk) O26_N0_S2 <=     O26_N0_S1  +  O26_N2_S1 ;
 logic signed [21:0] O26_N2_S2;		always @(posedge clk) O26_N2_S2 <=     O26_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O26_N0_S3;		always @(posedge clk) O26_N0_S3 <=     O26_N0_S2  +  O26_N2_S2 ;
 assign conv_mac_26 = O26_N0_S3;

logic signed [31:0] conv_mac_27;
logic signed [63:0] chainout_0_O27; 
logic signed [63:0] O27_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O27(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_27[7:0]),.ay( 9'sd7),.bx(input_fmap_27[15:8]),.by( 9'sd10),.cx(input_fmap_27[23:16]),.cy( 9'sd5),.dx(input_fmap_27[31:24]),.dy( 9'sd11),.chainin(63'd0),.result(O27_N0_S1),.chainout(chainout_0_O27));
logic signed [63:0] chainout_2_O27; 
logic signed [63:0] O27_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O27(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_27[39:32]),.ay( 9'sd17),.bx(input_fmap_27[47:40]),.by( 9'sd5),.cx(input_fmap_27[55:48]),.cy( 9'sd5),.dx(input_fmap_27[63:56]),.dy( 9'sd6),.chainin(63'd0),.result(O27_N2_S1),.chainout(chainout_2_O27));
logic signed [63:0] chainout_4_O27; 
logic signed [63:0] O27_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O27(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_27[71:64]),.ay( 9'sd2),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O27_N4_S1),.chainout(chainout_4_O27));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O27_N0_S2;		always @(posedge clk) O27_N0_S2 <=     O27_N0_S1  +  O27_N2_S1 ;
 logic signed [21:0] O27_N2_S2;		always @(posedge clk) O27_N2_S2 <=     O27_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O27_N0_S3;		always @(posedge clk) O27_N0_S3 <=     O27_N0_S2  +  O27_N2_S2 ;
 assign conv_mac_27 = O27_N0_S3;

logic signed [31:0] conv_mac_28;
logic signed [63:0] chainout_0_O28; 
logic signed [63:0] O28_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O28(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_28[7:0]),.ay( 9'sd8),.bx(input_fmap_28[15:8]),.by( 9'sd10),.cx(input_fmap_28[23:16]),.cy( 9'sd6),.dx(input_fmap_28[31:24]),.dy( 9'sd12),.chainin(63'd0),.result(O28_N0_S1),.chainout(chainout_0_O28));
logic signed [63:0] chainout_2_O28; 
logic signed [63:0] O28_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O28(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_28[39:32]),.ay( 9'sd14),.bx(input_fmap_28[47:40]),.by( 9'sd7),.cx(input_fmap_28[55:48]),.cy( 9'sd5),.dx(input_fmap_28[63:56]),.dy( 9'sd7),.chainin(63'd0),.result(O28_N2_S1),.chainout(chainout_2_O28));
logic signed [63:0] chainout_4_O28; 
logic signed [63:0] O28_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O28(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_28[71:64]),.ay( 9'sd3),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O28_N4_S1),.chainout(chainout_4_O28));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O28_N0_S2;		always @(posedge clk) O28_N0_S2 <=     O28_N0_S1  +  O28_N2_S1 ;
 logic signed [21:0] O28_N2_S2;		always @(posedge clk) O28_N2_S2 <=     O28_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O28_N0_S3;		always @(posedge clk) O28_N0_S3 <=     O28_N0_S2  +  O28_N2_S2 ;
 assign conv_mac_28 = O28_N0_S3;

logic signed [31:0] conv_mac_29;
logic signed [63:0] chainout_0_O29; 
logic signed [63:0] O29_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O29(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_29[7:0]),.ay( 9'sd7),.bx(input_fmap_29[15:8]),.by( 9'sd8),.cx(input_fmap_29[23:16]),.cy( 9'sd6),.dx(input_fmap_29[31:24]),.dy( 9'sd8),.chainin(63'd0),.result(O29_N0_S1),.chainout(chainout_0_O29));
logic signed [63:0] chainout_2_O29; 
logic signed [63:0] O29_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O29(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_29[39:32]),.ay( 9'sd9),.bx(input_fmap_29[47:40]),.by( 9'sd7),.cx(input_fmap_29[55:48]),.cy( 9'sd4),.dx(input_fmap_29[63:56]),.dy( 9'sd6),.chainin(63'd0),.result(O29_N2_S1),.chainout(chainout_2_O29));
logic signed [63:0] chainout_4_O29; 
logic signed [63:0] O29_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O29(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_29[71:64]),.ay( 9'sd2),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O29_N4_S1),.chainout(chainout_4_O29));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O29_N0_S2;		always @(posedge clk) O29_N0_S2 <=     O29_N0_S1  +  O29_N2_S1 ;
 logic signed [21:0] O29_N2_S2;		always @(posedge clk) O29_N2_S2 <=     O29_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O29_N0_S3;		always @(posedge clk) O29_N0_S3 <=     O29_N0_S2  +  O29_N2_S2 ;
 assign conv_mac_29 = O29_N0_S3;

logic signed [31:0] conv_mac_30;
logic signed [63:0] chainout_0_O30; 
logic signed [63:0] O30_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O30(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_30[7:0]),.ay( 9'sd9),.bx(input_fmap_30[15:8]),.by( 9'sd9),.cx(input_fmap_30[23:16]),.cy( 9'sd3),.dx(input_fmap_30[31:24]),.dy( 9'sd11),.chainin(63'd0),.result(O30_N0_S1),.chainout(chainout_0_O30));
logic signed [63:0] chainout_2_O30; 
logic signed [63:0] O30_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O30(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_30[39:32]),.ay( 9'sd15),.bx(input_fmap_30[47:40]),.by( 9'sd5),.cx(input_fmap_30[55:48]),.cy( 9'sd6),.dx(input_fmap_30[63:56]),.dy( 9'sd9),.chainin(63'd0),.result(O30_N2_S1),.chainout(chainout_2_O30));
logic signed [63:0] chainout_4_O30; 
logic signed [63:0] O30_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O30(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_30[71:64]),.ay( 9'sd5),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O30_N4_S1),.chainout(chainout_4_O30));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O30_N0_S2;		always @(posedge clk) O30_N0_S2 <=     O30_N0_S1  +  O30_N2_S1 ;
 logic signed [21:0] O30_N2_S2;		always @(posedge clk) O30_N2_S2 <=     O30_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O30_N0_S3;		always @(posedge clk) O30_N0_S3 <=     O30_N0_S2  +  O30_N2_S2 ;
 assign conv_mac_30 = O30_N0_S3;

logic signed [31:0] conv_mac_31;
logic signed [63:0] chainout_0_O31; 
logic signed [63:0] O31_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O31(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_31[7:0]),.ay( 9'sd8),.bx(input_fmap_31[15:8]),.by( 9'sd12),.cx(input_fmap_31[23:16]),.cy( 9'sd5),.dx(input_fmap_31[31:24]),.dy( 9'sd10),.chainin(63'd0),.result(O31_N0_S1),.chainout(chainout_0_O31));
logic signed [63:0] chainout_2_O31; 
logic signed [63:0] O31_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O31(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_31[39:32]),.ay( 9'sd18),.bx(input_fmap_31[47:40]),.by( 9'sd5),.cx(input_fmap_31[55:48]),.cy( 9'sd5),.dx(input_fmap_31[63:56]),.dy( 9'sd7),.chainin(63'd0),.result(O31_N2_S1),.chainout(chainout_2_O31));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O31_N0_S2;		always @(posedge clk) O31_N0_S2 <=     O31_N0_S1  +  O31_N2_S1 ;
 assign conv_mac_31 = O31_N0_S2;

logic valid_D1;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D1<= 0 ;
	else valid_D1<=valid;
end
logic valid_D2;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D2<= 0 ;
	else valid_D2<=valid_D1;
end
logic valid_D3;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D3<= 0 ;
	else valid_D3<=valid_D2;
end
logic valid_D4;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D4<= 0 ;
	else valid_D4<=valid_D3;
end
always_ff @(posedge clk) begin
	if (rstn == 0) ready <= 0 ;
	else ready <=valid_D4;
end
logic [31:0] bias_add_0;
assign bias_add_0 = conv_mac_0 + 7'd49;
logic [31:0] bias_add_1;
assign bias_add_1 = conv_mac_1 + 6'd22;
logic [31:0] bias_add_2;
assign bias_add_2 = conv_mac_2 + 3'd2;
logic [31:0] bias_add_3;
assign bias_add_3 = conv_mac_3 + 5'd9;
logic [31:0] bias_add_4;
assign bias_add_4 = conv_mac_4 - 5'd9;
logic [31:0] bias_add_5;
assign bias_add_5 = conv_mac_5 + 3'd3;
logic [31:0] bias_add_6;
assign bias_add_6 = conv_mac_6 + 5'd10;
logic [31:0] bias_add_7;
assign bias_add_7 = conv_mac_7 + 4'd4;
logic [31:0] bias_add_8;
assign bias_add_8 = conv_mac_8;
logic [31:0] bias_add_9;
assign bias_add_9 = conv_mac_9 - 2'd1;
logic [31:0] bias_add_10;
assign bias_add_10 = conv_mac_10 + 5'd9;
logic [31:0] bias_add_11;
assign bias_add_11 = conv_mac_11 + 4'd7;
logic [31:0] bias_add_12;
assign bias_add_12 = conv_mac_12;
logic [31:0] bias_add_13;
assign bias_add_13 = conv_mac_13 + 6'd18;
logic [31:0] bias_add_14;
assign bias_add_14 = conv_mac_14 + 6'd18;
logic [31:0] bias_add_15;
assign bias_add_15 = conv_mac_15 + 6'd27;
logic [31:0] bias_add_16;
assign bias_add_16 = conv_mac_16 + 5'd9;
logic [31:0] bias_add_17;
assign bias_add_17 = conv_mac_17 + 5'd13;
logic [31:0] bias_add_18;
assign bias_add_18 = conv_mac_18 + 8'd68;
logic [31:0] bias_add_19;
assign bias_add_19 = conv_mac_19 + 8'd87;
logic [31:0] bias_add_20;
assign bias_add_20 = conv_mac_20 + 6'd28;
logic [31:0] bias_add_21;
assign bias_add_21 = conv_mac_21 + 7'd36;
logic [31:0] bias_add_22;
assign bias_add_22 = conv_mac_22 + 6'd16;
logic [31:0] bias_add_23;
assign bias_add_23 = conv_mac_23 + 5'd14;
logic [31:0] bias_add_24;
assign bias_add_24 = conv_mac_24 + 6'd16;
logic [31:0] bias_add_25;
assign bias_add_25 = conv_mac_25 + 8'd86;
logic [31:0] bias_add_26;
assign bias_add_26 = conv_mac_26 + 6'd18;
logic [31:0] bias_add_27;
assign bias_add_27 = conv_mac_27 + 5'd13;
logic [31:0] bias_add_28;
assign bias_add_28 = conv_mac_28 + 5'd11;
logic [31:0] bias_add_29;
assign bias_add_29 = conv_mac_29 - 5'd13;
logic [31:0] bias_add_30;
assign bias_add_30 = conv_mac_30 + 5'd15;
logic [31:0] bias_add_31;
assign bias_add_31 = conv_mac_31 - 4'd5;

logic [7:0] relu_0;
assign relu_0[7:0] = (bias_add_0[31]==0) ? ((bias_add_0<3'd6) ? {{bias_add_0[31],bias_add_0[10:4]}} :'d6) : '0;
logic [7:0] relu_1;
assign relu_1[7:0] = (bias_add_1[31]==0) ? ((bias_add_1<3'd6) ? {{bias_add_1[31],bias_add_1[10:4]}} :'d6) : '0;
logic [7:0] relu_2;
assign relu_2[7:0] = (bias_add_2[31]==0) ? ((bias_add_2<3'd6) ? {{bias_add_2[31],bias_add_2[10:4]}} :'d6) : '0;
logic [7:0] relu_3;
assign relu_3[7:0] = (bias_add_3[31]==0) ? ((bias_add_3<3'd6) ? {{bias_add_3[31],bias_add_3[10:4]}} :'d6) : '0;
logic [7:0] relu_4;
assign relu_4[7:0] = (bias_add_4[31]==0) ? ((bias_add_4<3'd6) ? {{bias_add_4[31],bias_add_4[10:4]}} :'d6) : '0;
logic [7:0] relu_5;
assign relu_5[7:0] = (bias_add_5[31]==0) ? ((bias_add_5<3'd6) ? {{bias_add_5[31],bias_add_5[10:4]}} :'d6) : '0;
logic [7:0] relu_6;
assign relu_6[7:0] = (bias_add_6[31]==0) ? ((bias_add_6<3'd6) ? {{bias_add_6[31],bias_add_6[10:4]}} :'d6) : '0;
logic [7:0] relu_7;
assign relu_7[7:0] = (bias_add_7[31]==0) ? ((bias_add_7<3'd6) ? {{bias_add_7[31],bias_add_7[10:4]}} :'d6) : '0;
logic [7:0] relu_8;
assign relu_8[7:0] = (bias_add_8[31]==0) ? ((bias_add_8<3'd6) ? {{bias_add_8[31],bias_add_8[10:4]}} :'d6) : '0;
logic [7:0] relu_9;
assign relu_9[7:0] = (bias_add_9[31]==0) ? ((bias_add_9<3'd6) ? {{bias_add_9[31],bias_add_9[10:4]}} :'d6) : '0;
logic [7:0] relu_10;
assign relu_10[7:0] = (bias_add_10[31]==0) ? ((bias_add_10<3'd6) ? {{bias_add_10[31],bias_add_10[10:4]}} :'d6) : '0;
logic [7:0] relu_11;
assign relu_11[7:0] = (bias_add_11[31]==0) ? ((bias_add_11<3'd6) ? {{bias_add_11[31],bias_add_11[10:4]}} :'d6) : '0;
logic [7:0] relu_12;
assign relu_12[7:0] = (bias_add_12[31]==0) ? ((bias_add_12<3'd6) ? {{bias_add_12[31],bias_add_12[10:4]}} :'d6) : '0;
logic [7:0] relu_13;
assign relu_13[7:0] = (bias_add_13[31]==0) ? ((bias_add_13<3'd6) ? {{bias_add_13[31],bias_add_13[10:4]}} :'d6) : '0;
logic [7:0] relu_14;
assign relu_14[7:0] = (bias_add_14[31]==0) ? ((bias_add_14<3'd6) ? {{bias_add_14[31],bias_add_14[10:4]}} :'d6) : '0;
logic [7:0] relu_15;
assign relu_15[7:0] = (bias_add_15[31]==0) ? ((bias_add_15<3'd6) ? {{bias_add_15[31],bias_add_15[10:4]}} :'d6) : '0;
logic [7:0] relu_16;
assign relu_16[7:0] = (bias_add_16[31]==0) ? ((bias_add_16<3'd6) ? {{bias_add_16[31],bias_add_16[10:4]}} :'d6) : '0;
logic [7:0] relu_17;
assign relu_17[7:0] = (bias_add_17[31]==0) ? ((bias_add_17<3'd6) ? {{bias_add_17[31],bias_add_17[10:4]}} :'d6) : '0;
logic [7:0] relu_18;
assign relu_18[7:0] = (bias_add_18[31]==0) ? ((bias_add_18<3'd6) ? {{bias_add_18[31],bias_add_18[10:4]}} :'d6) : '0;
logic [7:0] relu_19;
assign relu_19[7:0] = (bias_add_19[31]==0) ? ((bias_add_19<3'd6) ? {{bias_add_19[31],bias_add_19[10:4]}} :'d6) : '0;
logic [7:0] relu_20;
assign relu_20[7:0] = (bias_add_20[31]==0) ? ((bias_add_20<3'd6) ? {{bias_add_20[31],bias_add_20[10:4]}} :'d6) : '0;
logic [7:0] relu_21;
assign relu_21[7:0] = (bias_add_21[31]==0) ? ((bias_add_21<3'd6) ? {{bias_add_21[31],bias_add_21[10:4]}} :'d6) : '0;
logic [7:0] relu_22;
assign relu_22[7:0] = (bias_add_22[31]==0) ? ((bias_add_22<3'd6) ? {{bias_add_22[31],bias_add_22[10:4]}} :'d6) : '0;
logic [7:0] relu_23;
assign relu_23[7:0] = (bias_add_23[31]==0) ? ((bias_add_23<3'd6) ? {{bias_add_23[31],bias_add_23[10:4]}} :'d6) : '0;
logic [7:0] relu_24;
assign relu_24[7:0] = (bias_add_24[31]==0) ? ((bias_add_24<3'd6) ? {{bias_add_24[31],bias_add_24[10:4]}} :'d6) : '0;
logic [7:0] relu_25;
assign relu_25[7:0] = (bias_add_25[31]==0) ? ((bias_add_25<3'd6) ? {{bias_add_25[31],bias_add_25[10:4]}} :'d6) : '0;
logic [7:0] relu_26;
assign relu_26[7:0] = (bias_add_26[31]==0) ? ((bias_add_26<3'd6) ? {{bias_add_26[31],bias_add_26[10:4]}} :'d6) : '0;
logic [7:0] relu_27;
assign relu_27[7:0] = (bias_add_27[31]==0) ? ((bias_add_27<3'd6) ? {{bias_add_27[31],bias_add_27[10:4]}} :'d6) : '0;
logic [7:0] relu_28;
assign relu_28[7:0] = (bias_add_28[31]==0) ? ((bias_add_28<3'd6) ? {{bias_add_28[31],bias_add_28[10:4]}} :'d6) : '0;
logic [7:0] relu_29;
assign relu_29[7:0] = (bias_add_29[31]==0) ? ((bias_add_29<3'd6) ? {{bias_add_29[31],bias_add_29[10:4]}} :'d6) : '0;
logic [7:0] relu_30;
assign relu_30[7:0] = (bias_add_30[31]==0) ? ((bias_add_30<3'd6) ? {{bias_add_30[31],bias_add_30[10:4]}} :'d6) : '0;
logic [7:0] relu_31;
assign relu_31[7:0] = (bias_add_31[31]==0) ? ((bias_add_31<3'd6) ? {{bias_add_31[31],bias_add_31[10:4]}} :'d6) : '0;

assign output_act = {
	relu_31,
	relu_30,
	relu_29,
	relu_28,
	relu_27,
	relu_26,
	relu_25,
	relu_24,
	relu_23,
	relu_22,
	relu_21,
	relu_20,
	relu_19,
	relu_18,
	relu_17,
	relu_16,
	relu_15,
	relu_14,
	relu_13,
	relu_12,
	relu_11,
	relu_10,
	relu_9,
	relu_8,
	relu_7,
	relu_6,
	relu_5,
	relu_4,
	relu_3,
	relu_2,
	relu_1,
	relu_0
};

endmodule
module conv7_dw (
    input logic clk,
    input logic rstn,
    input logic valid,
    input logic [64*72-1:0] input_act,
    output logic [512-1:0] output_act,
    output logic ready
);
logic we;
logic [8:0] zero_number; 
assign zero_number = 9'd0; 
logic [64*72-1:0] input_act_ff;
genvar i;
generate
for (i=0;i<64;i++)
    begin: genblk_12
        always_ff @(posedge clk) begin
            if (rstn == 0) begin
                input_act_ff[(i+1)*72-1:i*72] <= '0;
            end
            else begin
                input_act_ff[(i+1)*72-1:i*72] <= input_act[(i+1)*72-1:i*72];
            end
        end
    end
endgenerate
logic [71:0] input_fmap_0;
assign input_fmap_0 = input_act_ff[71:0];
logic [71:0] input_fmap_1;
assign input_fmap_1 = input_act_ff[143:72];
logic [71:0] input_fmap_2;
assign input_fmap_2 = input_act_ff[215:144];
logic [71:0] input_fmap_3;
assign input_fmap_3 = input_act_ff[287:216];
logic [71:0] input_fmap_4;
assign input_fmap_4 = input_act_ff[359:288];
logic [71:0] input_fmap_5;
assign input_fmap_5 = input_act_ff[431:360];
logic [71:0] input_fmap_6;
assign input_fmap_6 = input_act_ff[503:432];
logic [71:0] input_fmap_7;
assign input_fmap_7 = input_act_ff[575:504];
logic [71:0] input_fmap_8;
assign input_fmap_8 = input_act_ff[647:576];
logic [71:0] input_fmap_9;
assign input_fmap_9 = input_act_ff[719:648];
logic [71:0] input_fmap_10;
assign input_fmap_10 = input_act_ff[791:720];
logic [71:0] input_fmap_11;
assign input_fmap_11 = input_act_ff[863:792];
logic [71:0] input_fmap_12;
assign input_fmap_12 = input_act_ff[935:864];
logic [71:0] input_fmap_13;
assign input_fmap_13 = input_act_ff[1007:936];
logic [71:0] input_fmap_14;
assign input_fmap_14 = input_act_ff[1079:1008];
logic [71:0] input_fmap_15;
assign input_fmap_15 = input_act_ff[1151:1080];
logic [71:0] input_fmap_16;
assign input_fmap_16 = input_act_ff[1223:1152];
logic [71:0] input_fmap_17;
assign input_fmap_17 = input_act_ff[1295:1224];
logic [71:0] input_fmap_18;
assign input_fmap_18 = input_act_ff[1367:1296];
logic [71:0] input_fmap_19;
assign input_fmap_19 = input_act_ff[1439:1368];
logic [71:0] input_fmap_20;
assign input_fmap_20 = input_act_ff[1511:1440];
logic [71:0] input_fmap_21;
assign input_fmap_21 = input_act_ff[1583:1512];
logic [71:0] input_fmap_22;
assign input_fmap_22 = input_act_ff[1655:1584];
logic [71:0] input_fmap_23;
assign input_fmap_23 = input_act_ff[1727:1656];
logic [71:0] input_fmap_24;
assign input_fmap_24 = input_act_ff[1799:1728];
logic [71:0] input_fmap_25;
assign input_fmap_25 = input_act_ff[1871:1800];
logic [71:0] input_fmap_26;
assign input_fmap_26 = input_act_ff[1943:1872];
logic [71:0] input_fmap_27;
assign input_fmap_27 = input_act_ff[2015:1944];
logic [71:0] input_fmap_28;
assign input_fmap_28 = input_act_ff[2087:2016];
logic [71:0] input_fmap_29;
assign input_fmap_29 = input_act_ff[2159:2088];
logic [71:0] input_fmap_30;
assign input_fmap_30 = input_act_ff[2231:2160];
logic [71:0] input_fmap_31;
assign input_fmap_31 = input_act_ff[2303:2232];
logic [71:0] input_fmap_32;
assign input_fmap_32 = input_act_ff[2375:2304];
logic [71:0] input_fmap_33;
assign input_fmap_33 = input_act_ff[2447:2376];
logic [71:0] input_fmap_34;
assign input_fmap_34 = input_act_ff[2519:2448];
logic [71:0] input_fmap_35;
assign input_fmap_35 = input_act_ff[2591:2520];
logic [71:0] input_fmap_36;
assign input_fmap_36 = input_act_ff[2663:2592];
logic [71:0] input_fmap_37;
assign input_fmap_37 = input_act_ff[2735:2664];
logic [71:0] input_fmap_38;
assign input_fmap_38 = input_act_ff[2807:2736];
logic [71:0] input_fmap_39;
assign input_fmap_39 = input_act_ff[2879:2808];
logic [71:0] input_fmap_40;
assign input_fmap_40 = input_act_ff[2951:2880];
logic [71:0] input_fmap_41;
assign input_fmap_41 = input_act_ff[3023:2952];
logic [71:0] input_fmap_42;
assign input_fmap_42 = input_act_ff[3095:3024];
logic [71:0] input_fmap_43;
assign input_fmap_43 = input_act_ff[3167:3096];
logic [71:0] input_fmap_44;
assign input_fmap_44 = input_act_ff[3239:3168];
logic [71:0] input_fmap_45;
assign input_fmap_45 = input_act_ff[3311:3240];
logic [71:0] input_fmap_46;
assign input_fmap_46 = input_act_ff[3383:3312];
logic [71:0] input_fmap_47;
assign input_fmap_47 = input_act_ff[3455:3384];
logic [71:0] input_fmap_48;
assign input_fmap_48 = input_act_ff[3527:3456];
logic [71:0] input_fmap_49;
assign input_fmap_49 = input_act_ff[3599:3528];
logic [71:0] input_fmap_50;
assign input_fmap_50 = input_act_ff[3671:3600];
logic [71:0] input_fmap_51;
assign input_fmap_51 = input_act_ff[3743:3672];
logic [71:0] input_fmap_52;
assign input_fmap_52 = input_act_ff[3815:3744];
logic [71:0] input_fmap_53;
assign input_fmap_53 = input_act_ff[3887:3816];
logic [71:0] input_fmap_54;
assign input_fmap_54 = input_act_ff[3959:3888];
logic [71:0] input_fmap_55;
assign input_fmap_55 = input_act_ff[4031:3960];
logic [71:0] input_fmap_56;
assign input_fmap_56 = input_act_ff[4103:4032];
logic [71:0] input_fmap_57;
assign input_fmap_57 = input_act_ff[4175:4104];
logic [71:0] input_fmap_58;
assign input_fmap_58 = input_act_ff[4247:4176];
logic [71:0] input_fmap_59;
assign input_fmap_59 = input_act_ff[4319:4248];
logic [71:0] input_fmap_60;
assign input_fmap_60 = input_act_ff[4391:4320];
logic [71:0] input_fmap_61;
assign input_fmap_61 = input_act_ff[4463:4392];
logic [71:0] input_fmap_62;
assign input_fmap_62 = input_act_ff[4535:4464];
logic [71:0] input_fmap_63;
assign input_fmap_63 = input_act_ff[4607:4536];

logic signed [31:0] conv_mac_0;
logic signed [63:0] chainout_0_O0; 
logic signed [63:0] O0_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O0(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd2),.bx(input_fmap_0[15:8]),.by(-9'sd5),.cx(input_fmap_0[23:16]),.cy(-9'sd1),.dx(input_fmap_0[31:24]),.dy(-9'sd10),.chainin(63'd0),.result(O0_N0_S1),.chainout(chainout_0_O0));
logic signed [63:0] chainout_2_O0; 
logic signed [63:0] O0_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O0(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[39:32]),.ay(-9'sd4),.bx(input_fmap_0[47:40]),.by(-9'sd7),.cx(input_fmap_0[55:48]),.cy(-9'sd5),.dx(input_fmap_0[63:56]),.dy(-9'sd5),.chainin(63'd0),.result(O0_N2_S1),.chainout(chainout_2_O0));
logic signed [63:0] chainout_4_O0; 
logic signed [63:0] O0_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O0(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[71:64]),.ay(-9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O0_N4_S1),.chainout(chainout_4_O0));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O0_N0_S2;		always @(posedge clk) O0_N0_S2 <=     O0_N0_S1  +  O0_N2_S1 ;
 logic signed [21:0] O0_N2_S2;		always @(posedge clk) O0_N2_S2 <=     O0_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O0_N0_S3;		always @(posedge clk) O0_N0_S3 <=     O0_N0_S2  +  O0_N2_S2 ;
 assign conv_mac_0 = O0_N0_S3;

logic signed [31:0] conv_mac_1;
logic signed [63:0] chainout_0_O1; 
logic signed [63:0] O1_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O1(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay(-9'sd3),.bx(input_fmap_1[15:8]),.by(-9'sd16),.cx(input_fmap_1[23:16]),.cy(-9'sd1),.dx(input_fmap_1[31:24]),.dy( 9'sd8),.chainin(63'd0),.result(O1_N0_S1),.chainout(chainout_0_O1));
logic signed [63:0] chainout_2_O1; 
logic signed [63:0] O1_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O1(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[39:32]),.ay( 9'sd31),.bx(input_fmap_1[47:40]),.by(-9'sd22),.cx(input_fmap_1[55:48]),.cy( 9'sd3),.dx(input_fmap_1[63:56]),.dy( 9'sd4),.chainin(63'd0),.result(O1_N2_S1),.chainout(chainout_2_O1));
logic signed [63:0] chainout_4_O1; 
logic signed [63:0] O1_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O1(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[71:64]),.ay(-9'sd12),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O1_N4_S1),.chainout(chainout_4_O1));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O1_N0_S2;		always @(posedge clk) O1_N0_S2 <=     O1_N0_S1  +  O1_N2_S1 ;
 logic signed [21:0] O1_N2_S2;		always @(posedge clk) O1_N2_S2 <=     O1_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O1_N0_S3;		always @(posedge clk) O1_N0_S3 <=     O1_N0_S2  +  O1_N2_S2 ;
 assign conv_mac_1 = O1_N0_S3;

logic signed [31:0] conv_mac_2;
logic signed [63:0] chainout_0_O2; 
logic signed [63:0] O2_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O2(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_2[7:0]),.ay( 9'sd2),.bx(input_fmap_2[15:8]),.by(-9'sd14),.cx(input_fmap_2[23:16]),.cy(-9'sd2),.dx(input_fmap_2[31:24]),.dy(-9'sd5),.chainin(63'd0),.result(O2_N0_S1),.chainout(chainout_0_O2));
logic signed [63:0] chainout_2_O2; 
logic signed [63:0] O2_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O2(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_2[39:32]),.ay( 9'sd39),.bx(input_fmap_2[47:40]),.by(-9'sd8),.cx(input_fmap_2[55:48]),.cy(-9'sd15),.dx(input_fmap_2[63:56]),.dy( 9'sd4),.chainin(63'd0),.result(O2_N2_S1),.chainout(chainout_2_O2));
logic signed [63:0] chainout_4_O2; 
logic signed [63:0] O2_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O2(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_2[71:64]),.ay( 9'sd3),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O2_N4_S1),.chainout(chainout_4_O2));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O2_N0_S2;		always @(posedge clk) O2_N0_S2 <=     O2_N0_S1  +  O2_N2_S1 ;
 logic signed [21:0] O2_N2_S2;		always @(posedge clk) O2_N2_S2 <=     O2_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O2_N0_S3;		always @(posedge clk) O2_N0_S3 <=     O2_N0_S2  +  O2_N2_S2 ;
 assign conv_mac_2 = O2_N0_S3;

logic signed [31:0] conv_mac_3;
logic signed [63:0] chainout_0_O3; 
logic signed [63:0] O3_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O3(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_3[7:0]),.ay( 9'sd7),.bx(input_fmap_3[15:8]),.by( 9'sd15),.cx(input_fmap_3[31:24]),.cy( 9'sd14),.dx(input_fmap_3[39:32]),.dy(-9'sd1),.chainin(63'd0),.result(O3_N0_S1),.chainout(chainout_0_O3));
logic signed [63:0] chainout_2_O3; 
logic signed [63:0] O3_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O3(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_3[47:40]),.ay(-9'sd8),.bx(input_fmap_3[63:56]),.by(-9'sd11),.cx(input_fmap_3[71:64]),.cy(-9'sd7),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O3_N2_S1),.chainout(chainout_2_O3));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O3_N0_S2;		always @(posedge clk) O3_N0_S2 <=     O3_N0_S1  +  O3_N2_S1 ;
 assign conv_mac_3 = O3_N0_S2;

logic signed [31:0] conv_mac_4;
logic signed [63:0] chainout_0_O4; 
logic signed [63:0] O4_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O4(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_4[7:0]),.ay(-9'sd2),.bx(input_fmap_4[15:8]),.by(-9'sd12),.cx(input_fmap_4[23:16]),.cy(-9'sd9),.dx(input_fmap_4[31:24]),.dy(-9'sd6),.chainin(63'd0),.result(O4_N0_S1),.chainout(chainout_0_O4));
logic signed [63:0] chainout_2_O4; 
logic signed [63:0] O4_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O4(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_4[39:32]),.ay( 9'sd37),.bx(input_fmap_4[47:40]),.by( 9'sd3),.cx(input_fmap_4[55:48]),.cy(-9'sd6),.dx(input_fmap_4[63:56]),.dy( 9'sd10),.chainin(63'd0),.result(O4_N2_S1),.chainout(chainout_2_O4));
logic signed [63:0] chainout_4_O4; 
logic signed [63:0] O4_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O4(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_4[71:64]),.ay(-9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O4_N4_S1),.chainout(chainout_4_O4));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O4_N0_S2;		always @(posedge clk) O4_N0_S2 <=     O4_N0_S1  +  O4_N2_S1 ;
 logic signed [21:0] O4_N2_S2;		always @(posedge clk) O4_N2_S2 <=     O4_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O4_N0_S3;		always @(posedge clk) O4_N0_S3 <=     O4_N0_S2  +  O4_N2_S2 ;
 assign conv_mac_4 = O4_N0_S3;

logic signed [31:0] conv_mac_5;
logic signed [63:0] chainout_0_O5; 
logic signed [63:0] O5_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O5(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_5[15:8]),.ay( 9'sd4),.bx(input_fmap_5[23:16]),.by(-9'sd9),.cx(input_fmap_5[31:24]),.cy( 9'sd15),.dx(input_fmap_5[39:32]),.dy( 9'sd28),.chainin(63'd0),.result(O5_N0_S1),.chainout(chainout_0_O5));
logic signed [63:0] chainout_2_O5; 
logic signed [63:0] O5_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O5(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_5[47:40]),.ay(-9'sd17),.bx(input_fmap_5[55:48]),.by(-9'sd4),.cx(input_fmap_5[71:64]),.cy(-9'sd5),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O5_N2_S1),.chainout(chainout_2_O5));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O5_N0_S2;		always @(posedge clk) O5_N0_S2 <=     O5_N0_S1  +  O5_N2_S1 ;
 assign conv_mac_5 = O5_N0_S2;

logic signed [31:0] conv_mac_6;
logic signed [63:0] chainout_0_O6; 
logic signed [63:0] O6_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O6(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_6[7:0]),.ay(-9'sd10),.bx(input_fmap_6[15:8]),.by(-9'sd16),.cx(input_fmap_6[23:16]),.cy(-9'sd1),.dx(input_fmap_6[31:24]),.dy( 9'sd12),.chainin(63'd0),.result(O6_N0_S1),.chainout(chainout_0_O6));
logic signed [63:0] chainout_2_O6; 
logic signed [63:0] O6_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O6(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_6[39:32]),.ay( 9'sd22),.bx(input_fmap_6[47:40]),.by(-9'sd9),.cx(input_fmap_6[55:48]),.cy(-9'sd4),.dx(input_fmap_6[63:56]),.dy( 9'sd3),.chainin(63'd0),.result(O6_N2_S1),.chainout(chainout_2_O6));
logic signed [63:0] chainout_4_O6; 
logic signed [63:0] O6_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O6(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_6[71:64]),.ay(-9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O6_N4_S1),.chainout(chainout_4_O6));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O6_N0_S2;		always @(posedge clk) O6_N0_S2 <=     O6_N0_S1  +  O6_N2_S1 ;
 logic signed [21:0] O6_N2_S2;		always @(posedge clk) O6_N2_S2 <=     O6_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O6_N0_S3;		always @(posedge clk) O6_N0_S3 <=     O6_N0_S2  +  O6_N2_S2 ;
 assign conv_mac_6 = O6_N0_S3;

logic signed [31:0] conv_mac_7;
logic signed [63:0] chainout_0_O7; 
logic signed [63:0] O7_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O7(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_7[7:0]),.ay(-9'sd4),.bx(input_fmap_7[15:8]),.by(-9'sd9),.cx(input_fmap_7[23:16]),.cy( 9'sd3),.dx(input_fmap_7[31:24]),.dy(-9'sd6),.chainin(63'd0),.result(O7_N0_S1),.chainout(chainout_0_O7));
logic signed [63:0] chainout_2_O7; 
logic signed [63:0] O7_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O7(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_7[39:32]),.ay(-9'sd16),.bx(input_fmap_7[47:40]),.by( 9'sd2),.cx(input_fmap_7[55:48]),.cy(-9'sd1),.dx(input_fmap_7[63:56]),.dy(-9'sd6),.chainin(63'd0),.result(O7_N2_S1),.chainout(chainout_2_O7));
logic signed [63:0] chainout_4_O7; 
logic signed [63:0] O7_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O7(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_7[71:64]),.ay(-9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O7_N4_S1),.chainout(chainout_4_O7));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O7_N0_S2;		always @(posedge clk) O7_N0_S2 <=     O7_N0_S1  +  O7_N2_S1 ;
 logic signed [21:0] O7_N2_S2;		always @(posedge clk) O7_N2_S2 <=     O7_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O7_N0_S3;		always @(posedge clk) O7_N0_S3 <=     O7_N0_S2  +  O7_N2_S2 ;
 assign conv_mac_7 = O7_N0_S3;

logic signed [31:0] conv_mac_8;
logic signed [63:0] chainout_0_O8; 
logic signed [63:0] O8_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O8(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_8[7:0]),.ay( 9'sd3),.bx(input_fmap_8[15:8]),.by( 9'sd11),.cx(input_fmap_8[23:16]),.cy( 9'sd7),.dx(input_fmap_8[31:24]),.dy(-9'sd7),.chainin(63'd0),.result(O8_N0_S1),.chainout(chainout_0_O8));
logic signed [63:0] chainout_2_O8; 
logic signed [63:0] O8_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O8(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_8[39:32]),.ay(-9'sd25),.bx(input_fmap_8[47:40]),.by( 9'sd13),.cx(input_fmap_8[55:48]),.cy(-9'sd2),.dx(input_fmap_8[63:56]),.dy(-9'sd10),.chainin(63'd0),.result(O8_N2_S1),.chainout(chainout_2_O8));
logic signed [63:0] chainout_4_O8; 
logic signed [63:0] O8_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O8(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_8[71:64]),.ay(-9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O8_N4_S1),.chainout(chainout_4_O8));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O8_N0_S2;		always @(posedge clk) O8_N0_S2 <=     O8_N0_S1  +  O8_N2_S1 ;
 logic signed [21:0] O8_N2_S2;		always @(posedge clk) O8_N2_S2 <=     O8_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O8_N0_S3;		always @(posedge clk) O8_N0_S3 <=     O8_N0_S2  +  O8_N2_S2 ;
 assign conv_mac_8 = O8_N0_S3;

logic signed [31:0] conv_mac_9;
logic signed [63:0] chainout_0_O9; 
logic signed [63:0] O9_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O9(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_9[7:0]),.ay( 9'sd6),.bx(input_fmap_9[15:8]),.by(-9'sd4),.cx(input_fmap_9[23:16]),.cy(-9'sd6),.dx(input_fmap_9[31:24]),.dy( 9'sd22),.chainin(63'd0),.result(O9_N0_S1),.chainout(chainout_0_O9));
logic signed [63:0] chainout_2_O9; 
logic signed [63:0] O9_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O9(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_9[39:32]),.ay(-9'sd4),.bx(input_fmap_9[47:40]),.by(-9'sd7),.cx(input_fmap_9[55:48]),.cy( 9'sd4),.dx(input_fmap_9[63:56]),.dy(-9'sd8),.chainin(63'd0),.result(O9_N2_S1),.chainout(chainout_2_O9));
logic signed [63:0] chainout_4_O9; 
logic signed [63:0] O9_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O9(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_9[71:64]),.ay(-9'sd7),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O9_N4_S1),.chainout(chainout_4_O9));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O9_N0_S2;		always @(posedge clk) O9_N0_S2 <=     O9_N0_S1  +  O9_N2_S1 ;
 logic signed [21:0] O9_N2_S2;		always @(posedge clk) O9_N2_S2 <=     O9_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O9_N0_S3;		always @(posedge clk) O9_N0_S3 <=     O9_N0_S2  +  O9_N2_S2 ;
 assign conv_mac_9 = O9_N0_S3;

logic signed [31:0] conv_mac_10;
logic signed [63:0] chainout_0_O10; 
logic signed [63:0] O10_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O10(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_10[7:0]),.ay(-9'sd1),.bx(input_fmap_10[15:8]),.by( 9'sd8),.cx(input_fmap_10[23:16]),.cy( 9'sd2),.dx(input_fmap_10[31:24]),.dy( 9'sd6),.chainin(63'd0),.result(O10_N0_S1),.chainout(chainout_0_O10));
logic signed [63:0] chainout_2_O10; 
logic signed [63:0] O10_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O10(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_10[39:32]),.ay( 9'sd18),.bx(input_fmap_10[47:40]),.by( 9'sd5),.cx(input_fmap_10[55:48]),.cy(-9'sd4),.dx(input_fmap_10[63:56]),.dy(-9'sd1),.chainin(63'd0),.result(O10_N2_S1),.chainout(chainout_2_O10));
logic signed [63:0] chainout_4_O10; 
logic signed [63:0] O10_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O10(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_10[71:64]),.ay(-9'sd2),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O10_N4_S1),.chainout(chainout_4_O10));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O10_N0_S2;		always @(posedge clk) O10_N0_S2 <=     O10_N0_S1  +  O10_N2_S1 ;
 logic signed [21:0] O10_N2_S2;		always @(posedge clk) O10_N2_S2 <=     O10_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O10_N0_S3;		always @(posedge clk) O10_N0_S3 <=     O10_N0_S2  +  O10_N2_S2 ;
 assign conv_mac_10 = O10_N0_S3;

logic signed [31:0] conv_mac_11;
logic signed [63:0] chainout_0_O11; 
logic signed [63:0] O11_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O11(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_11[7:0]),.ay( 9'sd2),.bx(input_fmap_11[15:8]),.by( 9'sd2),.cx(input_fmap_11[23:16]),.cy(-9'sd11),.dx(input_fmap_11[31:24]),.dy( 9'sd14),.chainin(63'd0),.result(O11_N0_S1),.chainout(chainout_0_O11));
logic signed [63:0] chainout_2_O11; 
logic signed [63:0] O11_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O11(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_11[39:32]),.ay( 9'sd23),.bx(input_fmap_11[47:40]),.by( 9'sd3),.cx(input_fmap_11[55:48]),.cy( 9'sd3),.dx(input_fmap_11[63:56]),.dy( 9'sd7),.chainin(63'd0),.result(O11_N2_S1),.chainout(chainout_2_O11));
logic signed [63:0] chainout_4_O11; 
logic signed [63:0] O11_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O11(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_11[71:64]),.ay(-9'sd10),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O11_N4_S1),.chainout(chainout_4_O11));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O11_N0_S2;		always @(posedge clk) O11_N0_S2 <=     O11_N0_S1  +  O11_N2_S1 ;
 logic signed [21:0] O11_N2_S2;		always @(posedge clk) O11_N2_S2 <=     O11_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O11_N0_S3;		always @(posedge clk) O11_N0_S3 <=     O11_N0_S2  +  O11_N2_S2 ;
 assign conv_mac_11 = O11_N0_S3;

logic signed [31:0] conv_mac_12;
logic signed [63:0] chainout_0_O12; 
logic signed [63:0] O12_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O12(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_12[7:0]),.ay( 9'sd12),.bx(input_fmap_12[15:8]),.by(-9'sd7),.cx(input_fmap_12[23:16]),.cy(-9'sd5),.dx(input_fmap_12[31:24]),.dy( 9'sd25),.chainin(63'd0),.result(O12_N0_S1),.chainout(chainout_0_O12));
logic signed [63:0] chainout_2_O12; 
logic signed [63:0] O12_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O12(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_12[39:32]),.ay(-9'sd22),.bx(input_fmap_12[47:40]),.by(-9'sd3),.cx(input_fmap_12[55:48]),.cy( 9'sd8),.dx(input_fmap_12[71:64]),.dy(-9'sd6),.chainin(63'd0),.result(O12_N2_S1),.chainout(chainout_2_O12));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O12_N0_S2;		always @(posedge clk) O12_N0_S2 <=     O12_N0_S1  +  O12_N2_S1 ;
 assign conv_mac_12 = O12_N0_S2;

logic signed [31:0] conv_mac_13;
logic signed [63:0] chainout_0_O13; 
logic signed [63:0] O13_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O13(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_13[7:0]),.ay(-9'sd14),.bx(input_fmap_13[15:8]),.by(-9'sd8),.cx(input_fmap_13[31:24]),.cy(-9'sd13),.dx(input_fmap_13[39:32]),.dy(-9'sd9),.chainin(63'd0),.result(O13_N0_S1),.chainout(chainout_0_O13));
logic signed [63:0] chainout_2_O13; 
logic signed [63:0] O13_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O13(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_13[47:40]),.ay( 9'sd14),.bx(input_fmap_13[63:56]),.by( 9'sd3),.cx(input_fmap_13[71:64]),.cy( 9'sd10),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O13_N2_S1),.chainout(chainout_2_O13));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O13_N0_S2;		always @(posedge clk) O13_N0_S2 <=     O13_N0_S1  +  O13_N2_S1 ;
 assign conv_mac_13 = O13_N0_S2;

logic signed [31:0] conv_mac_14;
logic signed [63:0] chainout_0_O14; 
logic signed [63:0] O14_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O14(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_14[7:0]),.ay(-9'sd3),.bx(input_fmap_14[15:8]),.by(-9'sd1),.cx(input_fmap_14[23:16]),.cy(-9'sd1),.dx(input_fmap_14[31:24]),.dy( 9'sd5),.chainin(63'd0),.result(O14_N0_S1),.chainout(chainout_0_O14));
logic signed [63:0] chainout_2_O14; 
logic signed [63:0] O14_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O14(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_14[39:32]),.ay(-9'sd19),.bx(input_fmap_14[47:40]),.by( 9'sd5),.cx(input_fmap_14[55:48]),.cy( 9'sd6),.dx(input_fmap_14[63:56]),.dy(-9'sd5),.chainin(63'd0),.result(O14_N2_S1),.chainout(chainout_2_O14));
logic signed [63:0] chainout_4_O14; 
logic signed [63:0] O14_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O14(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_14[71:64]),.ay(-9'sd3),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O14_N4_S1),.chainout(chainout_4_O14));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O14_N0_S2;		always @(posedge clk) O14_N0_S2 <=     O14_N0_S1  +  O14_N2_S1 ;
 logic signed [21:0] O14_N2_S2;		always @(posedge clk) O14_N2_S2 <=     O14_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O14_N0_S3;		always @(posedge clk) O14_N0_S3 <=     O14_N0_S2  +  O14_N2_S2 ;
 assign conv_mac_14 = O14_N0_S3;

logic signed [31:0] conv_mac_15;
logic signed [63:0] chainout_0_O15; 
logic signed [63:0] O15_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O15(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_15[7:0]),.ay(-9'sd2),.bx(input_fmap_15[15:8]),.by(-9'sd2),.cx(input_fmap_15[23:16]),.cy( 9'sd1),.dx(input_fmap_15[31:24]),.dy(-9'sd6),.chainin(63'd0),.result(O15_N0_S1),.chainout(chainout_0_O15));
logic signed [63:0] chainout_2_O15; 
logic signed [63:0] O15_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O15(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_15[39:32]),.ay(-9'sd23),.bx(input_fmap_15[47:40]),.by( 9'sd5),.cx(input_fmap_15[55:48]),.cy(-9'sd5),.dx(input_fmap_15[63:56]),.dy( 9'sd3),.chainin(63'd0),.result(O15_N2_S1),.chainout(chainout_2_O15));
logic signed [63:0] chainout_4_O15; 
logic signed [63:0] O15_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O15(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_15[71:64]),.ay( 9'sd6),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O15_N4_S1),.chainout(chainout_4_O15));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O15_N0_S2;		always @(posedge clk) O15_N0_S2 <=     O15_N0_S1  +  O15_N2_S1 ;
 logic signed [21:0] O15_N2_S2;		always @(posedge clk) O15_N2_S2 <=     O15_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O15_N0_S3;		always @(posedge clk) O15_N0_S3 <=     O15_N0_S2  +  O15_N2_S2 ;
 assign conv_mac_15 = O15_N0_S3;

logic signed [31:0] conv_mac_16;
logic signed [63:0] chainout_0_O16; 
logic signed [63:0] O16_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O16(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_16[7:0]),.ay(-9'sd5),.bx(input_fmap_16[15:8]),.by(-9'sd4),.cx(input_fmap_16[23:16]),.cy( 9'sd8),.dx(input_fmap_16[31:24]),.dy(-9'sd18),.chainin(63'd0),.result(O16_N0_S1),.chainout(chainout_0_O16));
logic signed [63:0] chainout_2_O16; 
logic signed [63:0] O16_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O16(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_16[39:32]),.ay(-9'sd6),.bx(input_fmap_16[47:40]),.by( 9'sd22),.cx(input_fmap_16[55:48]),.cy(-9'sd7),.dx(input_fmap_16[71:64]),.dy( 9'sd7),.chainin(63'd0),.result(O16_N2_S1),.chainout(chainout_2_O16));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O16_N0_S2;		always @(posedge clk) O16_N0_S2 <=     O16_N0_S1  +  O16_N2_S1 ;
 assign conv_mac_16 = O16_N0_S2;

logic signed [31:0] conv_mac_17;
logic signed [63:0] chainout_0_O17; 
logic signed [63:0] O17_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O17(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_17[7:0]),.ay( 9'sd3),.bx(input_fmap_17[15:8]),.by(-9'sd5),.cx(input_fmap_17[23:16]),.cy( 9'sd2),.dx(input_fmap_17[31:24]),.dy( 9'sd1),.chainin(63'd0),.result(O17_N0_S1),.chainout(chainout_0_O17));
logic signed [63:0] chainout_2_O17; 
logic signed [63:0] O17_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O17(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_17[39:32]),.ay(-9'sd28),.bx(input_fmap_17[47:40]),.by( 9'sd2),.cx(input_fmap_17[55:48]),.cy( 9'sd1),.dx(input_fmap_17[63:56]),.dy(-9'sd1),.chainin(63'd0),.result(O17_N2_S1),.chainout(chainout_2_O17));
logic signed [63:0] chainout_4_O17; 
logic signed [63:0] O17_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O17(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_17[71:64]),.ay(-9'sd3),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O17_N4_S1),.chainout(chainout_4_O17));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O17_N0_S2;		always @(posedge clk) O17_N0_S2 <=     O17_N0_S1  +  O17_N2_S1 ;
 logic signed [21:0] O17_N2_S2;		always @(posedge clk) O17_N2_S2 <=     O17_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O17_N0_S3;		always @(posedge clk) O17_N0_S3 <=     O17_N0_S2  +  O17_N2_S2 ;
 assign conv_mac_17 = O17_N0_S3;

logic signed [31:0] conv_mac_18;
logic signed [63:0] chainout_0_O18; 
logic signed [63:0] O18_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O18(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_18[7:0]),.ay(-9'sd5),.bx(input_fmap_18[15:8]),.by(-9'sd2),.cx(input_fmap_18[23:16]),.cy( 9'sd2),.dx(input_fmap_18[31:24]),.dy(-9'sd1),.chainin(63'd0),.result(O18_N0_S1),.chainout(chainout_0_O18));
logic signed [63:0] chainout_2_O18; 
logic signed [63:0] O18_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O18(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_18[39:32]),.ay( 9'sd30),.bx(input_fmap_18[47:40]),.by(-9'sd4),.cx(input_fmap_18[55:48]),.cy( 9'sd2),.dx(input_fmap_18[63:56]),.dy( 9'sd2),.chainin(63'd0),.result(O18_N2_S1),.chainout(chainout_2_O18));
logic signed [63:0] chainout_4_O18; 
logic signed [63:0] O18_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O18(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_18[71:64]),.ay(-9'sd5),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O18_N4_S1),.chainout(chainout_4_O18));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O18_N0_S2;		always @(posedge clk) O18_N0_S2 <=     O18_N0_S1  +  O18_N2_S1 ;
 logic signed [21:0] O18_N2_S2;		always @(posedge clk) O18_N2_S2 <=     O18_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O18_N0_S3;		always @(posedge clk) O18_N0_S3 <=     O18_N0_S2  +  O18_N2_S2 ;
 assign conv_mac_18 = O18_N0_S3;

logic signed [31:0] conv_mac_19;
logic signed [63:0] chainout_0_O19; 
logic signed [63:0] O19_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O19(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_19[7:0]),.ay( 9'sd1),.bx(input_fmap_19[15:8]),.by(-9'sd9),.cx(input_fmap_19[23:16]),.cy(-9'sd2),.dx(input_fmap_19[31:24]),.dy(-9'sd7),.chainin(63'd0),.result(O19_N0_S1),.chainout(chainout_0_O19));
logic signed [63:0] chainout_2_O19; 
logic signed [63:0] O19_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O19(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_19[39:32]),.ay(-9'sd20),.bx(input_fmap_19[47:40]),.by( 9'sd6),.cx(input_fmap_19[63:56]),.cy( 9'sd8),.dx(input_fmap_19[71:64]),.dy( 9'sd2),.chainin(63'd0),.result(O19_N2_S1),.chainout(chainout_2_O19));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O19_N0_S2;		always @(posedge clk) O19_N0_S2 <=     O19_N0_S1  +  O19_N2_S1 ;
 assign conv_mac_19 = O19_N0_S2;

logic signed [31:0] conv_mac_20;
logic signed [63:0] chainout_0_O20; 
logic signed [63:0] O20_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O20(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_20[7:0]),.ay(-9'sd7),.bx(input_fmap_20[15:8]),.by(-9'sd16),.cx(input_fmap_20[23:16]),.cy(-9'sd4),.dx(input_fmap_20[31:24]),.dy( 9'sd5),.chainin(63'd0),.result(O20_N0_S1),.chainout(chainout_0_O20));
logic signed [63:0] chainout_2_O20; 
logic signed [63:0] O20_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O20(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_20[39:32]),.ay( 9'sd37),.bx(input_fmap_20[47:40]),.by(-9'sd5),.cx(input_fmap_20[55:48]),.cy( 9'sd2),.dx(input_fmap_20[63:56]),.dy( 9'sd10),.chainin(63'd0),.result(O20_N2_S1),.chainout(chainout_2_O20));
logic signed [63:0] chainout_4_O20; 
logic signed [63:0] O20_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O20(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_20[71:64]),.ay(-9'sd3),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O20_N4_S1),.chainout(chainout_4_O20));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O20_N0_S2;		always @(posedge clk) O20_N0_S2 <=     O20_N0_S1  +  O20_N2_S1 ;
 logic signed [21:0] O20_N2_S2;		always @(posedge clk) O20_N2_S2 <=     O20_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O20_N0_S3;		always @(posedge clk) O20_N0_S3 <=     O20_N0_S2  +  O20_N2_S2 ;
 assign conv_mac_20 = O20_N0_S3;

logic signed [31:0] conv_mac_21;
logic signed [63:0] chainout_0_O21; 
logic signed [63:0] O21_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O21(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_21[7:0]),.ay(-9'sd7),.bx(input_fmap_21[15:8]),.by( 9'sd9),.cx(input_fmap_21[23:16]),.cy(-9'sd1),.dx(input_fmap_21[31:24]),.dy(-9'sd4),.chainin(63'd0),.result(O21_N0_S1),.chainout(chainout_0_O21));
logic signed [63:0] chainout_2_O21; 
logic signed [63:0] O21_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O21(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_21[39:32]),.ay( 9'sd35),.bx(input_fmap_21[47:40]),.by(-9'sd1),.cx(input_fmap_21[55:48]),.cy(-9'sd10),.dx(input_fmap_21[63:56]),.dy(-9'sd17),.chainin(63'd0),.result(O21_N2_S1),.chainout(chainout_2_O21));
logic signed [63:0] chainout_4_O21; 
logic signed [63:0] O21_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O21(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_21[71:64]),.ay(-9'sd6),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O21_N4_S1),.chainout(chainout_4_O21));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O21_N0_S2;		always @(posedge clk) O21_N0_S2 <=     O21_N0_S1  +  O21_N2_S1 ;
 logic signed [21:0] O21_N2_S2;		always @(posedge clk) O21_N2_S2 <=     O21_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O21_N0_S3;		always @(posedge clk) O21_N0_S3 <=     O21_N0_S2  +  O21_N2_S2 ;
 assign conv_mac_21 = O21_N0_S3;

logic signed [31:0] conv_mac_22;
logic signed [63:0] chainout_0_O22; 
logic signed [63:0] O22_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O22(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_22[7:0]),.ay(-9'sd1),.bx(input_fmap_22[15:8]),.by(-9'sd8),.cx(input_fmap_22[23:16]),.cy( 9'sd1),.dx(input_fmap_22[31:24]),.dy( 9'sd3),.chainin(63'd0),.result(O22_N0_S1),.chainout(chainout_0_O22));
logic signed [63:0] chainout_2_O22; 
logic signed [63:0] O22_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O22(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_22[39:32]),.ay(-9'sd18),.bx(input_fmap_22[47:40]),.by(-9'sd5),.cx(input_fmap_22[55:48]),.cy( 9'sd8),.dx(input_fmap_22[63:56]),.dy( 9'sd5),.chainin(63'd0),.result(O22_N2_S1),.chainout(chainout_2_O22));
logic signed [63:0] chainout_4_O22; 
logic signed [63:0] O22_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O22(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_22[71:64]),.ay( 9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O22_N4_S1),.chainout(chainout_4_O22));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O22_N0_S2;		always @(posedge clk) O22_N0_S2 <=     O22_N0_S1  +  O22_N2_S1 ;
 logic signed [21:0] O22_N2_S2;		always @(posedge clk) O22_N2_S2 <=     O22_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O22_N0_S3;		always @(posedge clk) O22_N0_S3 <=     O22_N0_S2  +  O22_N2_S2 ;
 assign conv_mac_22 = O22_N0_S3;

logic signed [31:0] conv_mac_23;
logic signed [63:0] chainout_0_O23; 
logic signed [63:0] O23_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O23(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_23[7:0]),.ay( 9'sd10),.bx(input_fmap_23[15:8]),.by( 9'sd24),.cx(input_fmap_23[23:16]),.cy( 9'sd8),.dx(input_fmap_23[31:24]),.dy(-9'sd5),.chainin(63'd0),.result(O23_N0_S1),.chainout(chainout_0_O23));
logic signed [63:0] chainout_2_O23; 
logic signed [63:0] O23_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O23(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_23[39:32]),.ay(-9'sd7),.bx(input_fmap_23[47:40]),.by(-9'sd11),.cx(input_fmap_23[55:48]),.cy(-9'sd4),.dx(input_fmap_23[63:56]),.dy(-9'sd13),.chainin(63'd0),.result(O23_N2_S1),.chainout(chainout_2_O23));
logic signed [63:0] chainout_4_O23; 
logic signed [63:0] O23_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O23(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_23[71:64]),.ay(-9'sd5),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O23_N4_S1),.chainout(chainout_4_O23));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O23_N0_S2;		always @(posedge clk) O23_N0_S2 <=     O23_N0_S1  +  O23_N2_S1 ;
 logic signed [21:0] O23_N2_S2;		always @(posedge clk) O23_N2_S2 <=     O23_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O23_N0_S3;		always @(posedge clk) O23_N0_S3 <=     O23_N0_S2  +  O23_N2_S2 ;
 assign conv_mac_23 = O23_N0_S3;

logic signed [31:0] conv_mac_24;
logic signed [63:0] chainout_0_O24; 
logic signed [63:0] O24_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O24(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_24[7:0]),.ay(-9'sd17),.bx(input_fmap_24[15:8]),.by( 9'sd51),.cx(input_fmap_24[23:16]),.cy( 9'sd5),.dx(input_fmap_24[31:24]),.dy(-9'sd4),.chainin(63'd0),.result(O24_N0_S1),.chainout(chainout_0_O24));
logic signed [63:0] chainout_2_O24; 
logic signed [63:0] O24_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O24(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_24[39:32]),.ay(-9'sd1),.bx(input_fmap_24[47:40]),.by(-9'sd1),.cx(input_fmap_24[55:48]),.cy(-9'sd4),.dx(input_fmap_24[63:56]),.dy(-9'sd10),.chainin(63'd0),.result(O24_N2_S1),.chainout(chainout_2_O24));
logic signed [63:0] chainout_4_O24; 
logic signed [63:0] O24_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O24(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_24[71:64]),.ay(-9'sd5),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O24_N4_S1),.chainout(chainout_4_O24));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O24_N0_S2;		always @(posedge clk) O24_N0_S2 <=     O24_N0_S1  +  O24_N2_S1 ;
 logic signed [21:0] O24_N2_S2;		always @(posedge clk) O24_N2_S2 <=     O24_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O24_N0_S3;		always @(posedge clk) O24_N0_S3 <=     O24_N0_S2  +  O24_N2_S2 ;
 assign conv_mac_24 = O24_N0_S3;

logic signed [31:0] conv_mac_25;
logic signed [63:0] chainout_0_O25; 
logic signed [63:0] O25_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O25(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_25[7:0]),.ay( 9'sd11),.bx(input_fmap_25[15:8]),.by(-9'sd8),.cx(input_fmap_25[23:16]),.cy(-9'sd4),.dx(input_fmap_25[31:24]),.dy( 9'sd33),.chainin(63'd0),.result(O25_N0_S1),.chainout(chainout_0_O25));
logic signed [63:0] chainout_2_O25; 
logic signed [63:0] O25_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O25(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_25[39:32]),.ay(-9'sd9),.bx(input_fmap_25[47:40]),.by(-9'sd21),.cx(input_fmap_25[55:48]),.cy( 9'sd7),.dx(input_fmap_25[63:56]),.dy(-9'sd4),.chainin(63'd0),.result(O25_N2_S1),.chainout(chainout_2_O25));
logic signed [63:0] chainout_4_O25; 
logic signed [63:0] O25_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O25(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_25[71:64]),.ay(-9'sd5),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O25_N4_S1),.chainout(chainout_4_O25));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O25_N0_S2;		always @(posedge clk) O25_N0_S2 <=     O25_N0_S1  +  O25_N2_S1 ;
 logic signed [21:0] O25_N2_S2;		always @(posedge clk) O25_N2_S2 <=     O25_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O25_N0_S3;		always @(posedge clk) O25_N0_S3 <=     O25_N0_S2  +  O25_N2_S2 ;
 assign conv_mac_25 = O25_N0_S3;

logic signed [31:0] conv_mac_26;
logic signed [63:0] chainout_0_O26; 
logic signed [63:0] O26_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O26(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_26[7:0]),.ay( 9'sd7),.bx(input_fmap_26[15:8]),.by(-9'sd8),.cx(input_fmap_26[23:16]),.cy(-9'sd2),.dx(input_fmap_26[31:24]),.dy( 9'sd32),.chainin(63'd0),.result(O26_N0_S1),.chainout(chainout_0_O26));
logic signed [63:0] chainout_2_O26; 
logic signed [63:0] O26_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O26(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_26[39:32]),.ay(-9'sd4),.bx(input_fmap_26[47:40]),.by(-9'sd26),.cx(input_fmap_26[55:48]),.cy( 9'sd5),.dx(input_fmap_26[63:56]),.dy( 9'sd2),.chainin(63'd0),.result(O26_N2_S1),.chainout(chainout_2_O26));
logic signed [63:0] chainout_4_O26; 
logic signed [63:0] O26_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O26(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_26[71:64]),.ay(-9'sd6),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O26_N4_S1),.chainout(chainout_4_O26));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O26_N0_S2;		always @(posedge clk) O26_N0_S2 <=     O26_N0_S1  +  O26_N2_S1 ;
 logic signed [21:0] O26_N2_S2;		always @(posedge clk) O26_N2_S2 <=     O26_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O26_N0_S3;		always @(posedge clk) O26_N0_S3 <=     O26_N0_S2  +  O26_N2_S2 ;
 assign conv_mac_26 = O26_N0_S3;

logic signed [31:0] conv_mac_27;
logic signed [63:0] chainout_0_O27; 
logic signed [63:0] O27_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O27(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_27[15:8]),.ay( 9'sd1),.bx(input_fmap_27[23:16]),.by( 9'sd2),.cx(input_fmap_27[31:24]),.cy(-9'sd6),.dx(input_fmap_27[39:32]),.dy(-9'sd24),.chainin(63'd0),.result(O27_N0_S1),.chainout(chainout_0_O27));
logic signed [63:0] chainout_2_O27; 
logic signed [63:0] O27_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O27(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_27[55:48]),.ay(-9'sd3),.bx(input_fmap_27[71:64]),.by( 9'sd11),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O27_N2_S1),.chainout(chainout_2_O27));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O27_N0_S2;		always @(posedge clk) O27_N0_S2 <=     O27_N0_S1  +  O27_N2_S1 ;
 assign conv_mac_27 = O27_N0_S2;

logic signed [31:0] conv_mac_28;
logic signed [63:0] chainout_0_O28; 
logic signed [63:0] O28_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O28(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_28[7:0]),.ay(-9'sd3),.bx(input_fmap_28[15:8]),.by( 9'sd5),.cx(input_fmap_28[23:16]),.cy(-9'sd9),.dx(input_fmap_28[31:24]),.dy( 9'sd11),.chainin(63'd0),.result(O28_N0_S1),.chainout(chainout_0_O28));
logic signed [63:0] chainout_2_O28; 
logic signed [63:0] O28_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O28(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_28[39:32]),.ay( 9'sd19),.bx(input_fmap_28[47:40]),.by( 9'sd4),.cx(input_fmap_28[55:48]),.cy(-9'sd1),.dx(input_fmap_28[63:56]),.dy(-9'sd5),.chainin(63'd0),.result(O28_N2_S1),.chainout(chainout_2_O28));
logic signed [63:0] chainout_4_O28; 
logic signed [63:0] O28_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O28(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_28[71:64]),.ay(-9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O28_N4_S1),.chainout(chainout_4_O28));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O28_N0_S2;		always @(posedge clk) O28_N0_S2 <=     O28_N0_S1  +  O28_N2_S1 ;
 logic signed [21:0] O28_N2_S2;		always @(posedge clk) O28_N2_S2 <=     O28_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O28_N0_S3;		always @(posedge clk) O28_N0_S3 <=     O28_N0_S2  +  O28_N2_S2 ;
 assign conv_mac_28 = O28_N0_S3;

logic signed [31:0] conv_mac_29;
logic signed [63:0] chainout_0_O29; 
logic signed [63:0] O29_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O29(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_29[7:0]),.ay( 9'sd4),.bx(input_fmap_29[15:8]),.by( 9'sd29),.cx(input_fmap_29[23:16]),.cy( 9'sd8),.dx(input_fmap_29[31:24]),.dy(-9'sd8),.chainin(63'd0),.result(O29_N0_S1),.chainout(chainout_0_O29));
logic signed [63:0] chainout_2_O29; 
logic signed [63:0] O29_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O29(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_29[39:32]),.ay(-9'sd13),.bx(input_fmap_29[47:40]),.by(-9'sd2),.cx(input_fmap_29[55:48]),.cy(-9'sd3),.dx(input_fmap_29[63:56]),.dy(-9'sd15),.chainin(63'd0),.result(O29_N2_S1),.chainout(chainout_2_O29));
logic signed [63:0] chainout_4_O29; 
logic signed [63:0] O29_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O29(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_29[71:64]),.ay(-9'sd2),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O29_N4_S1),.chainout(chainout_4_O29));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O29_N0_S2;		always @(posedge clk) O29_N0_S2 <=     O29_N0_S1  +  O29_N2_S1 ;
 logic signed [21:0] O29_N2_S2;		always @(posedge clk) O29_N2_S2 <=     O29_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O29_N0_S3;		always @(posedge clk) O29_N0_S3 <=     O29_N0_S2  +  O29_N2_S2 ;
 assign conv_mac_29 = O29_N0_S3;

logic signed [31:0] conv_mac_30;
logic signed [63:0] chainout_0_O30; 
logic signed [63:0] O30_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O30(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_30[7:0]),.ay( 9'sd14),.bx(input_fmap_30[15:8]),.by( 9'sd24),.cx(input_fmap_30[23:16]),.cy( 9'sd9),.dx(input_fmap_30[31:24]),.dy(-9'sd17),.chainin(63'd0),.result(O30_N0_S1),.chainout(chainout_0_O30));
logic signed [63:0] chainout_2_O30; 
logic signed [63:0] O30_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O30(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_30[39:32]),.ay(-9'sd10),.bx(input_fmap_30[55:48]),.by(-9'sd3),.cx(input_fmap_30[63:56]),.cy(-9'sd11),.dx(input_fmap_30[71:64]),.dy(-9'sd4),.chainin(63'd0),.result(O30_N2_S1),.chainout(chainout_2_O30));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O30_N0_S2;		always @(posedge clk) O30_N0_S2 <=     O30_N0_S1  +  O30_N2_S1 ;
 assign conv_mac_30 = O30_N0_S2;

logic signed [31:0] conv_mac_31;
logic signed [63:0] chainout_0_O31; 
logic signed [63:0] O31_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O31(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_31[7:0]),.ay( 9'sd5),.bx(input_fmap_31[15:8]),.by(-9'sd6),.cx(input_fmap_31[23:16]),.cy( 9'sd5),.dx(input_fmap_31[31:24]),.dy( 9'sd2),.chainin(63'd0),.result(O31_N0_S1),.chainout(chainout_0_O31));
logic signed [63:0] chainout_2_O31; 
logic signed [63:0] O31_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O31(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_31[39:32]),.ay(-9'sd38),.bx(input_fmap_31[55:48]),.by( 9'sd5),.cx(input_fmap_31[63:56]),.cy( 9'sd9),.dx(input_fmap_31[71:64]),.dy( 9'sd2),.chainin(63'd0),.result(O31_N2_S1),.chainout(chainout_2_O31));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O31_N0_S2;		always @(posedge clk) O31_N0_S2 <=     O31_N0_S1  +  O31_N2_S1 ;
 assign conv_mac_31 = O31_N0_S2;

logic signed [31:0] conv_mac_32;
logic signed [63:0] chainout_0_O32; 
logic signed [63:0] O32_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O32(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_32[7:0]),.ay(-9'sd3),.bx(input_fmap_32[15:8]),.by(-9'sd2),.cx(input_fmap_32[23:16]),.cy( 9'sd1),.dx(input_fmap_32[31:24]),.dy( 9'sd4),.chainin(63'd0),.result(O32_N0_S1),.chainout(chainout_0_O32));
logic signed [63:0] chainout_2_O32; 
logic signed [63:0] O32_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O32(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_32[39:32]),.ay( 9'sd4),.bx(input_fmap_32[47:40]),.by( 9'sd4),.cx(input_fmap_32[55:48]),.cy(-9'sd12),.dx(input_fmap_32[63:56]),.dy(-9'sd11),.chainin(63'd0),.result(O32_N2_S1),.chainout(chainout_2_O32));
logic signed [63:0] chainout_4_O32; 
logic signed [63:0] O32_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O32(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_32[71:64]),.ay(-9'sd9),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O32_N4_S1),.chainout(chainout_4_O32));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O32_N0_S2;		always @(posedge clk) O32_N0_S2 <=     O32_N0_S1  +  O32_N2_S1 ;
 logic signed [21:0] O32_N2_S2;		always @(posedge clk) O32_N2_S2 <=     O32_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O32_N0_S3;		always @(posedge clk) O32_N0_S3 <=     O32_N0_S2  +  O32_N2_S2 ;
 assign conv_mac_32 = O32_N0_S3;

logic signed [31:0] conv_mac_33;
logic signed [63:0] chainout_0_O33; 
logic signed [63:0] O33_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O33(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_33[7:0]),.ay( 9'sd9),.bx(input_fmap_33[15:8]),.by(-9'sd2),.cx(input_fmap_33[23:16]),.cy(-9'sd5),.dx(input_fmap_33[31:24]),.dy( 9'sd24),.chainin(63'd0),.result(O33_N0_S1),.chainout(chainout_0_O33));
logic signed [63:0] chainout_2_O33; 
logic signed [63:0] O33_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O33(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_33[39:32]),.ay( 9'sd7),.bx(input_fmap_33[47:40]),.by(-9'sd28),.cx(input_fmap_33[55:48]),.cy( 9'sd8),.dx(input_fmap_33[63:56]),.dy(-9'sd9),.chainin(63'd0),.result(O33_N2_S1),.chainout(chainout_2_O33));
logic signed [63:0] chainout_4_O33; 
logic signed [63:0] O33_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O33(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_33[71:64]),.ay(-9'sd3),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O33_N4_S1),.chainout(chainout_4_O33));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O33_N0_S2;		always @(posedge clk) O33_N0_S2 <=     O33_N0_S1  +  O33_N2_S1 ;
 logic signed [21:0] O33_N2_S2;		always @(posedge clk) O33_N2_S2 <=     O33_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O33_N0_S3;		always @(posedge clk) O33_N0_S3 <=     O33_N0_S2  +  O33_N2_S2 ;
 assign conv_mac_33 = O33_N0_S3;

logic signed [31:0] conv_mac_34;
logic signed [63:0] chainout_0_O34; 
logic signed [63:0] O34_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O34(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_34[7:0]),.ay(-9'sd4),.bx(input_fmap_34[15:8]),.by( 9'sd7),.cx(input_fmap_34[23:16]),.cy( 9'sd2),.dx(input_fmap_34[31:24]),.dy( 9'sd9),.chainin(63'd0),.result(O34_N0_S1),.chainout(chainout_0_O34));
logic signed [63:0] chainout_2_O34; 
logic signed [63:0] O34_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O34(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_34[39:32]),.ay( 9'sd20),.bx(input_fmap_34[47:40]),.by(-9'sd4),.cx(input_fmap_34[55:48]),.cy(-9'sd1),.dx(input_fmap_34[63:56]),.dy(-9'sd10),.chainin(63'd0),.result(O34_N2_S1),.chainout(chainout_2_O34));
logic signed [63:0] chainout_4_O34; 
logic signed [63:0] O34_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O34(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_34[71:64]),.ay(-9'sd2),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O34_N4_S1),.chainout(chainout_4_O34));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O34_N0_S2;		always @(posedge clk) O34_N0_S2 <=     O34_N0_S1  +  O34_N2_S1 ;
 logic signed [21:0] O34_N2_S2;		always @(posedge clk) O34_N2_S2 <=     O34_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O34_N0_S3;		always @(posedge clk) O34_N0_S3 <=     O34_N0_S2  +  O34_N2_S2 ;
 assign conv_mac_34 = O34_N0_S3;

logic signed [31:0] conv_mac_35;
logic signed [63:0] chainout_0_O35; 
logic signed [63:0] O35_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O35(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_35[7:0]),.ay( 9'sd1),.bx(input_fmap_35[15:8]),.by( 9'sd9),.cx(input_fmap_35[23:16]),.cy(-9'sd5),.dx(input_fmap_35[31:24]),.dy( 9'sd4),.chainin(63'd0),.result(O35_N0_S1),.chainout(chainout_0_O35));
logic signed [63:0] chainout_2_O35; 
logic signed [63:0] O35_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O35(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_35[39:32]),.ay( 9'sd25),.bx(input_fmap_35[47:40]),.by(-9'sd2),.cx(input_fmap_35[55:48]),.cy(-9'sd6),.dx(input_fmap_35[63:56]),.dy(-9'sd7),.chainin(63'd0),.result(O35_N2_S1),.chainout(chainout_2_O35));
logic signed [63:0] chainout_4_O35; 
logic signed [63:0] O35_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O35(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_35[71:64]),.ay(-9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O35_N4_S1),.chainout(chainout_4_O35));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O35_N0_S2;		always @(posedge clk) O35_N0_S2 <=     O35_N0_S1  +  O35_N2_S1 ;
 logic signed [21:0] O35_N2_S2;		always @(posedge clk) O35_N2_S2 <=     O35_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O35_N0_S3;		always @(posedge clk) O35_N0_S3 <=     O35_N0_S2  +  O35_N2_S2 ;
 assign conv_mac_35 = O35_N0_S3;

logic signed [31:0] conv_mac_36;
logic signed [63:0] chainout_0_O36; 
logic signed [63:0] O36_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O36(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_36[7:0]),.ay( 9'sd1),.bx(input_fmap_36[15:8]),.by(-9'sd7),.cx(input_fmap_36[23:16]),.cy(-9'sd3),.dx(input_fmap_36[31:24]),.dy(-9'sd5),.chainin(63'd0),.result(O36_N0_S1),.chainout(chainout_0_O36));
logic signed [63:0] chainout_2_O36; 
logic signed [63:0] O36_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O36(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_36[39:32]),.ay(-9'sd19),.bx(input_fmap_36[47:40]),.by(-9'sd4),.cx(input_fmap_36[55:48]),.cy( 9'sd5),.dx(input_fmap_36[63:56]),.dy( 9'sd25),.chainin(63'd0),.result(O36_N2_S1),.chainout(chainout_2_O36));
logic signed [63:0] chainout_4_O36; 
logic signed [63:0] O36_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O36(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_36[71:64]),.ay( 9'sd6),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O36_N4_S1),.chainout(chainout_4_O36));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O36_N0_S2;		always @(posedge clk) O36_N0_S2 <=     O36_N0_S1  +  O36_N2_S1 ;
 logic signed [21:0] O36_N2_S2;		always @(posedge clk) O36_N2_S2 <=     O36_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O36_N0_S3;		always @(posedge clk) O36_N0_S3 <=     O36_N0_S2  +  O36_N2_S2 ;
 assign conv_mac_36 = O36_N0_S3;

logic signed [31:0] conv_mac_37;
logic signed [63:0] chainout_0_O37; 
logic signed [63:0] O37_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O37(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_37[7:0]),.ay(-9'sd2),.bx(input_fmap_37[15:8]),.by(-9'sd16),.cx(input_fmap_37[23:16]),.cy(-9'sd3),.dx(input_fmap_37[31:24]),.dy(-9'sd5),.chainin(63'd0),.result(O37_N0_S1),.chainout(chainout_0_O37));
logic signed [63:0] chainout_2_O37; 
logic signed [63:0] O37_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O37(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_37[39:32]),.ay(-9'sd14),.bx(input_fmap_37[47:40]),.by(-9'sd1),.cx(input_fmap_37[55:48]),.cy( 9'sd2),.dx(input_fmap_37[63:56]),.dy( 9'sd30),.chainin(63'd0),.result(O37_N2_S1),.chainout(chainout_2_O37));
logic signed [63:0] chainout_4_O37; 
logic signed [63:0] O37_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O37(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_37[71:64]),.ay( 9'sd4),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O37_N4_S1),.chainout(chainout_4_O37));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O37_N0_S2;		always @(posedge clk) O37_N0_S2 <=     O37_N0_S1  +  O37_N2_S1 ;
 logic signed [21:0] O37_N2_S2;		always @(posedge clk) O37_N2_S2 <=     O37_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O37_N0_S3;		always @(posedge clk) O37_N0_S3 <=     O37_N0_S2  +  O37_N2_S2 ;
 assign conv_mac_37 = O37_N0_S3;

logic signed [31:0] conv_mac_38;
logic signed [63:0] chainout_0_O38; 
logic signed [63:0] O38_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O38(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_38[7:0]),.ay(-9'sd2),.bx(input_fmap_38[15:8]),.by(-9'sd27),.cx(input_fmap_38[23:16]),.cy(-9'sd2),.dx(input_fmap_38[31:24]),.dy( 9'sd1),.chainin(63'd0),.result(O38_N0_S1),.chainout(chainout_0_O38));
logic signed [63:0] chainout_2_O38; 
logic signed [63:0] O38_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O38(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_38[39:32]),.ay(-9'sd1),.bx(input_fmap_38[47:40]),.by( 9'sd5),.cx(input_fmap_38[55:48]),.cy( 9'sd3),.dx(input_fmap_38[63:56]),.dy( 9'sd20),.chainin(63'd0),.result(O38_N2_S1),.chainout(chainout_2_O38));
logic signed [63:0] chainout_4_O38; 
logic signed [63:0] O38_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O38(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_38[71:64]),.ay( 9'sd6),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O38_N4_S1),.chainout(chainout_4_O38));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O38_N0_S2;		always @(posedge clk) O38_N0_S2 <=     O38_N0_S1  +  O38_N2_S1 ;
 logic signed [21:0] O38_N2_S2;		always @(posedge clk) O38_N2_S2 <=     O38_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O38_N0_S3;		always @(posedge clk) O38_N0_S3 <=     O38_N0_S2  +  O38_N2_S2 ;
 assign conv_mac_38 = O38_N0_S3;

logic signed [31:0] conv_mac_39;
logic signed [63:0] chainout_0_O39; 
logic signed [63:0] O39_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O39(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_39[7:0]),.ay(-9'sd9),.bx(input_fmap_39[15:8]),.by( 9'sd2),.cx(input_fmap_39[23:16]),.cy( 9'sd6),.dx(input_fmap_39[31:24]),.dy(-9'sd20),.chainin(63'd0),.result(O39_N0_S1),.chainout(chainout_0_O39));
logic signed [63:0] chainout_2_O39; 
logic signed [63:0] O39_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O39(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_39[39:32]),.ay(-9'sd4),.bx(input_fmap_39[47:40]),.by( 9'sd26),.cx(input_fmap_39[55:48]),.cy(-9'sd7),.dx(input_fmap_39[63:56]),.dy(-9'sd5),.chainin(63'd0),.result(O39_N2_S1),.chainout(chainout_2_O39));
logic signed [63:0] chainout_4_O39; 
logic signed [63:0] O39_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O39(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_39[71:64]),.ay( 9'sd8),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O39_N4_S1),.chainout(chainout_4_O39));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O39_N0_S2;		always @(posedge clk) O39_N0_S2 <=     O39_N0_S1  +  O39_N2_S1 ;
 logic signed [21:0] O39_N2_S2;		always @(posedge clk) O39_N2_S2 <=     O39_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O39_N0_S3;		always @(posedge clk) O39_N0_S3 <=     O39_N0_S2  +  O39_N2_S2 ;
 assign conv_mac_39 = O39_N0_S3;

logic signed [31:0] conv_mac_40;
logic signed [63:0] chainout_0_O40; 
logic signed [63:0] O40_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O40(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_40[7:0]),.ay(-9'sd11),.bx(input_fmap_40[15:8]),.by(-9'sd5),.cx(input_fmap_40[23:16]),.cy( 9'sd12),.dx(input_fmap_40[31:24]),.dy(-9'sd26),.chainin(63'd0),.result(O40_N0_S1),.chainout(chainout_0_O40));
logic signed [63:0] chainout_2_O40; 
logic signed [63:0] O40_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O40(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_40[39:32]),.ay(-9'sd2),.bx(input_fmap_40[47:40]),.by( 9'sd27),.cx(input_fmap_40[55:48]),.cy(-9'sd4),.dx(input_fmap_40[63:56]),.dy(-9'sd3),.chainin(63'd0),.result(O40_N2_S1),.chainout(chainout_2_O40));
logic signed [63:0] chainout_4_O40; 
logic signed [63:0] O40_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O40(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_40[71:64]),.ay( 9'sd9),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O40_N4_S1),.chainout(chainout_4_O40));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O40_N0_S2;		always @(posedge clk) O40_N0_S2 <=     O40_N0_S1  +  O40_N2_S1 ;
 logic signed [21:0] O40_N2_S2;		always @(posedge clk) O40_N2_S2 <=     O40_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O40_N0_S3;		always @(posedge clk) O40_N0_S3 <=     O40_N0_S2  +  O40_N2_S2 ;
 assign conv_mac_40 = O40_N0_S3;

logic signed [31:0] conv_mac_41;
logic signed [63:0] chainout_0_O41; 
logic signed [63:0] O41_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O41(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_41[7:0]),.ay( 9'sd2),.bx(input_fmap_41[15:8]),.by(-9'sd1),.cx(input_fmap_41[23:16]),.cy( 9'sd2),.dx(input_fmap_41[31:24]),.dy( 9'sd1),.chainin(63'd0),.result(O41_N0_S1),.chainout(chainout_0_O41));
logic signed [63:0] chainout_2_O41; 
logic signed [63:0] O41_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O41(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_41[39:32]),.ay(-9'sd20),.bx(input_fmap_41[47:40]),.by( 9'sd5),.cx(input_fmap_41[55:48]),.cy(-9'sd11),.dx(input_fmap_41[63:56]),.dy(-9'sd2),.chainin(63'd0),.result(O41_N2_S1),.chainout(chainout_2_O41));
logic signed [63:0] chainout_4_O41; 
logic signed [63:0] O41_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O41(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_41[71:64]),.ay( 9'sd6),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O41_N4_S1),.chainout(chainout_4_O41));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O41_N0_S2;		always @(posedge clk) O41_N0_S2 <=     O41_N0_S1  +  O41_N2_S1 ;
 logic signed [21:0] O41_N2_S2;		always @(posedge clk) O41_N2_S2 <=     O41_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O41_N0_S3;		always @(posedge clk) O41_N0_S3 <=     O41_N0_S2  +  O41_N2_S2 ;
 assign conv_mac_41 = O41_N0_S3;

logic signed [31:0] conv_mac_42;
logic signed [63:0] chainout_0_O42; 
logic signed [63:0] O42_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O42(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_42[7:0]),.ay(-9'sd11),.bx(input_fmap_42[15:8]),.by(-9'sd6),.cx(input_fmap_42[23:16]),.cy(-9'sd6),.dx(input_fmap_42[31:24]),.dy(-9'sd7),.chainin(63'd0),.result(O42_N0_S1),.chainout(chainout_0_O42));
logic signed [63:0] chainout_2_O42; 
logic signed [63:0] O42_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O42(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_42[39:32]),.ay( 9'sd43),.bx(input_fmap_42[47:40]),.by(-9'sd11),.cx(input_fmap_42[55:48]),.cy(-9'sd3),.dx(input_fmap_42[63:56]),.dy(-9'sd4),.chainin(63'd0),.result(O42_N2_S1),.chainout(chainout_2_O42));
logic signed [63:0] chainout_4_O42; 
logic signed [63:0] O42_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O42(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_42[71:64]),.ay( 9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O42_N4_S1),.chainout(chainout_4_O42));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O42_N0_S2;		always @(posedge clk) O42_N0_S2 <=     O42_N0_S1  +  O42_N2_S1 ;
 logic signed [21:0] O42_N2_S2;		always @(posedge clk) O42_N2_S2 <=     O42_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O42_N0_S3;		always @(posedge clk) O42_N0_S3 <=     O42_N0_S2  +  O42_N2_S2 ;
 assign conv_mac_42 = O42_N0_S3;

logic signed [31:0] conv_mac_43;
logic signed [63:0] chainout_0_O43; 
logic signed [63:0] O43_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O43(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_43[7:0]),.ay(-9'sd10),.bx(input_fmap_43[15:8]),.by( 9'sd9),.cx(input_fmap_43[23:16]),.cy(-9'sd3),.dx(input_fmap_43[39:32]),.dy( 9'sd41),.chainin(63'd0),.result(O43_N0_S1),.chainout(chainout_0_O43));
logic signed [63:0] chainout_2_O43; 
logic signed [63:0] O43_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O43(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_43[47:40]),.ay(-9'sd5),.bx(input_fmap_43[55:48]),.by( 9'sd5),.cx(input_fmap_43[63:56]),.cy(-9'sd16),.dx(input_fmap_43[71:64]),.dy(-9'sd1),.chainin(63'd0),.result(O43_N2_S1),.chainout(chainout_2_O43));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O43_N0_S2;		always @(posedge clk) O43_N0_S2 <=     O43_N0_S1  +  O43_N2_S1 ;
 assign conv_mac_43 = O43_N0_S2;

logic signed [31:0] conv_mac_44;
logic signed [63:0] chainout_0_O44; 
logic signed [63:0] O44_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O44(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_44[7:0]),.ay( 9'sd2),.bx(input_fmap_44[15:8]),.by(-9'sd6),.cx(input_fmap_44[23:16]),.cy( 9'sd1),.dx(input_fmap_44[31:24]),.dy(-9'sd10),.chainin(63'd0),.result(O44_N0_S1),.chainout(chainout_0_O44));
logic signed [63:0] chainout_2_O44; 
logic signed [63:0] O44_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O44(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_44[39:32]),.ay(-9'sd15),.bx(input_fmap_44[47:40]),.by(-9'sd1),.cx(input_fmap_44[55:48]),.cy( 9'sd1),.dx(input_fmap_44[63:56]),.dy( 9'sd2),.chainin(63'd0),.result(O44_N2_S1),.chainout(chainout_2_O44));
logic signed [63:0] chainout_4_O44; 
logic signed [63:0] O44_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O44(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_44[71:64]),.ay( 9'sd3),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O44_N4_S1),.chainout(chainout_4_O44));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O44_N0_S2;		always @(posedge clk) O44_N0_S2 <=     O44_N0_S1  +  O44_N2_S1 ;
 logic signed [21:0] O44_N2_S2;		always @(posedge clk) O44_N2_S2 <=     O44_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O44_N0_S3;		always @(posedge clk) O44_N0_S3 <=     O44_N0_S2  +  O44_N2_S2 ;
 assign conv_mac_44 = O44_N0_S3;

logic signed [31:0] conv_mac_45;
logic signed [63:0] chainout_0_O45; 
logic signed [63:0] O45_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O45(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_45[7:0]),.ay(-9'sd2),.bx(input_fmap_45[15:8]),.by( 9'sd7),.cx(input_fmap_45[23:16]),.cy( 9'sd7),.dx(input_fmap_45[31:24]),.dy(-9'sd12),.chainin(63'd0),.result(O45_N0_S1),.chainout(chainout_0_O45));
logic signed [63:0] chainout_2_O45; 
logic signed [63:0] O45_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O45(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_45[39:32]),.ay(-9'sd1),.bx(input_fmap_45[47:40]),.by( 9'sd15),.cx(input_fmap_45[55:48]),.cy(-9'sd7),.dx(input_fmap_45[63:56]),.dy(-9'sd14),.chainin(63'd0),.result(O45_N2_S1),.chainout(chainout_2_O45));
logic signed [63:0] chainout_4_O45; 
logic signed [63:0] O45_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O45(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_45[71:64]),.ay( 9'sd3),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O45_N4_S1),.chainout(chainout_4_O45));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O45_N0_S2;		always @(posedge clk) O45_N0_S2 <=     O45_N0_S1  +  O45_N2_S1 ;
 logic signed [21:0] O45_N2_S2;		always @(posedge clk) O45_N2_S2 <=     O45_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O45_N0_S3;		always @(posedge clk) O45_N0_S3 <=     O45_N0_S2  +  O45_N2_S2 ;
 assign conv_mac_45 = O45_N0_S3;

logic signed [31:0] conv_mac_46;
logic signed [63:0] chainout_0_O46; 
logic signed [63:0] O46_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O46(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_46[7:0]),.ay(-9'sd1),.bx(input_fmap_46[15:8]),.by(-9'sd3),.cx(input_fmap_46[23:16]),.cy( 9'sd1),.dx(input_fmap_46[31:24]),.dy(-9'sd10),.chainin(63'd0),.result(O46_N0_S1),.chainout(chainout_0_O46));
logic signed [63:0] chainout_2_O46; 
logic signed [63:0] O46_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O46(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_46[39:32]),.ay( 9'sd66),.bx(input_fmap_46[47:40]),.by(-9'sd11),.cx(input_fmap_46[55:48]),.cy(-9'sd2),.dx(input_fmap_46[63:56]),.dy(-9'sd7),.chainin(63'd0),.result(O46_N2_S1),.chainout(chainout_2_O46));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O46_N0_S2;		always @(posedge clk) O46_N0_S2 <=     O46_N0_S1  +  O46_N2_S1 ;
 assign conv_mac_46 = O46_N0_S2;

logic signed [31:0] conv_mac_47;
logic signed [63:0] chainout_0_O47; 
logic signed [63:0] O47_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O47(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_47[7:0]),.ay(-9'sd6),.bx(input_fmap_47[23:16]),.by(-9'sd10),.cx(input_fmap_47[31:24]),.cy( 9'sd11),.dx(input_fmap_47[39:32]),.dy( 9'sd34),.chainin(63'd0),.result(O47_N0_S1),.chainout(chainout_0_O47));
logic signed [63:0] chainout_2_O47; 
logic signed [63:0] O47_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O47(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_47[47:40]),.ay(-9'sd7),.bx(input_fmap_47[55:48]),.by(-9'sd1),.cx(input_fmap_47[63:56]),.cy( 9'sd8),.dx(input_fmap_47[71:64]),.dy(-9'sd4),.chainin(63'd0),.result(O47_N2_S1),.chainout(chainout_2_O47));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O47_N0_S2;		always @(posedge clk) O47_N0_S2 <=     O47_N0_S1  +  O47_N2_S1 ;
 assign conv_mac_47 = O47_N0_S2;

logic signed [31:0] conv_mac_48;
logic signed [63:0] chainout_0_O48; 
logic signed [63:0] O48_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O48(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_48[7:0]),.ay(-9'sd9),.bx(input_fmap_48[15:8]),.by(-9'sd10),.cx(input_fmap_48[23:16]),.cy(-9'sd7),.dx(input_fmap_48[31:24]),.dy( 9'sd10),.chainin(63'd0),.result(O48_N0_S1),.chainout(chainout_0_O48));
logic signed [63:0] chainout_2_O48; 
logic signed [63:0] O48_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O48(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_48[39:32]),.ay( 9'sd27),.bx(input_fmap_48[47:40]),.by(-9'sd4),.cx(input_fmap_48[55:48]),.cy(-9'sd5),.dx(input_fmap_48[63:56]),.dy(-9'sd2),.chainin(63'd0),.result(O48_N2_S1),.chainout(chainout_2_O48));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O48_N0_S2;		always @(posedge clk) O48_N0_S2 <=     O48_N0_S1  +  O48_N2_S1 ;
 assign conv_mac_48 = O48_N0_S2;

logic signed [31:0] conv_mac_49;
logic signed [63:0] chainout_0_O49; 
logic signed [63:0] O49_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O49(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_49[7:0]),.ay( 9'sd10),.bx(input_fmap_49[15:8]),.by( 9'sd20),.cx(input_fmap_49[23:16]),.cy( 9'sd3),.dx(input_fmap_49[31:24]),.dy(-9'sd4),.chainin(63'd0),.result(O49_N0_S1),.chainout(chainout_0_O49));
logic signed [63:0] chainout_2_O49; 
logic signed [63:0] O49_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O49(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_49[47:40]),.ay(-9'sd5),.bx(input_fmap_49[55:48]),.by(-9'sd7),.cx(input_fmap_49[63:56]),.cy(-9'sd22),.dx(input_fmap_49[71:64]),.dy(-9'sd5),.chainin(63'd0),.result(O49_N2_S1),.chainout(chainout_2_O49));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O49_N0_S2;		always @(posedge clk) O49_N0_S2 <=     O49_N0_S1  +  O49_N2_S1 ;
 assign conv_mac_49 = O49_N0_S2;

logic signed [31:0] conv_mac_50;
logic signed [63:0] chainout_0_O50; 
logic signed [63:0] O50_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O50(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_50[7:0]),.ay(-9'sd2),.bx(input_fmap_50[15:8]),.by( 9'sd3),.cx(input_fmap_50[23:16]),.cy( 9'sd7),.dx(input_fmap_50[31:24]),.dy(-9'sd6),.chainin(63'd0),.result(O50_N0_S1),.chainout(chainout_0_O50));
logic signed [63:0] chainout_2_O50; 
logic signed [63:0] O50_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O50(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_50[39:32]),.ay(-9'sd21),.bx(input_fmap_50[47:40]),.by( 9'sd13),.cx(input_fmap_50[55:48]),.cy(-9'sd6),.dx(input_fmap_50[63:56]),.dy(-9'sd6),.chainin(63'd0),.result(O50_N2_S1),.chainout(chainout_2_O50));
logic signed [63:0] chainout_4_O50; 
logic signed [63:0] O50_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O50(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_50[71:64]),.ay( 9'sd10),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O50_N4_S1),.chainout(chainout_4_O50));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O50_N0_S2;		always @(posedge clk) O50_N0_S2 <=     O50_N0_S1  +  O50_N2_S1 ;
 logic signed [21:0] O50_N2_S2;		always @(posedge clk) O50_N2_S2 <=     O50_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O50_N0_S3;		always @(posedge clk) O50_N0_S3 <=     O50_N0_S2  +  O50_N2_S2 ;
 assign conv_mac_50 = O50_N0_S3;

logic signed [31:0] conv_mac_51;
logic signed [63:0] chainout_0_O51; 
logic signed [63:0] O51_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O51(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_51[7:0]),.ay( 9'sd2),.bx(input_fmap_51[23:16]),.by( 9'sd1),.cx(input_fmap_51[31:24]),.cy(-9'sd5),.dx(input_fmap_51[39:32]),.dy( 9'sd36),.chainin(63'd0),.result(O51_N0_S1),.chainout(chainout_0_O51));
logic signed [63:0] chainout_2_O51; 
logic signed [63:0] O51_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O51(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_51[47:40]),.ay(-9'sd7),.bx(input_fmap_51[55:48]),.by(-9'sd2),.cx(input_fmap_51[63:56]),.cy(-9'sd11),.dx(input_fmap_51[71:64]),.dy(-9'sd2),.chainin(63'd0),.result(O51_N2_S1),.chainout(chainout_2_O51));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O51_N0_S2;		always @(posedge clk) O51_N0_S2 <=     O51_N0_S1  +  O51_N2_S1 ;
 assign conv_mac_51 = O51_N0_S2;

logic signed [31:0] conv_mac_52;
logic signed [63:0] chainout_0_O52; 
logic signed [63:0] O52_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O52(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_52[7:0]),.ay(-9'sd5),.bx(input_fmap_52[15:8]),.by(-9'sd7),.cx(input_fmap_52[23:16]),.cy(-9'sd2),.dx(input_fmap_52[31:24]),.dy( 9'sd4),.chainin(63'd0),.result(O52_N0_S1),.chainout(chainout_0_O52));
logic signed [63:0] chainout_2_O52; 
logic signed [63:0] O52_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O52(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_52[39:32]),.ay( 9'sd39),.bx(input_fmap_52[47:40]),.by(-9'sd15),.cx(input_fmap_52[55:48]),.cy(-9'sd2),.dx(input_fmap_52[63:56]),.dy(-9'sd3),.chainin(63'd0),.result(O52_N2_S1),.chainout(chainout_2_O52));
logic signed [63:0] chainout_4_O52; 
logic signed [63:0] O52_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O52(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_52[71:64]),.ay( 9'sd2),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O52_N4_S1),.chainout(chainout_4_O52));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O52_N0_S2;		always @(posedge clk) O52_N0_S2 <=     O52_N0_S1  +  O52_N2_S1 ;
 logic signed [21:0] O52_N2_S2;		always @(posedge clk) O52_N2_S2 <=     O52_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O52_N0_S3;		always @(posedge clk) O52_N0_S3 <=     O52_N0_S2  +  O52_N2_S2 ;
 assign conv_mac_52 = O52_N0_S3;

logic signed [31:0] conv_mac_53;
logic signed [63:0] chainout_0_O53; 
logic signed [63:0] O53_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O53(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_53[7:0]),.ay( 9'sd12),.bx(input_fmap_53[15:8]),.by(-9'sd14),.cx(input_fmap_53[23:16]),.cy(-9'sd2),.dx(input_fmap_53[31:24]),.dy(-9'sd16),.chainin(63'd0),.result(O53_N0_S1),.chainout(chainout_0_O53));
logic signed [63:0] chainout_2_O53; 
logic signed [63:0] O53_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O53(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_53[39:32]),.ay( 9'sd42),.bx(input_fmap_53[47:40]),.by(-9'sd11),.cx(input_fmap_53[55:48]),.cy(-9'sd6),.dx(input_fmap_53[63:56]),.dy(-9'sd3),.chainin(63'd0),.result(O53_N2_S1),.chainout(chainout_2_O53));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O53_N0_S2;		always @(posedge clk) O53_N0_S2 <=     O53_N0_S1  +  O53_N2_S1 ;
 assign conv_mac_53 = O53_N0_S2;

logic signed [31:0] conv_mac_54;
logic signed [63:0] chainout_0_O54; 
logic signed [63:0] O54_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O54(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_54[7:0]),.ay( 9'sd7),.bx(input_fmap_54[15:8]),.by( 9'sd11),.cx(input_fmap_54[23:16]),.cy(-9'sd5),.dx(input_fmap_54[31:24]),.dy( 9'sd15),.chainin(63'd0),.result(O54_N0_S1),.chainout(chainout_0_O54));
logic signed [63:0] chainout_2_O54; 
logic signed [63:0] O54_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O54(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_54[39:32]),.ay(-9'sd5),.bx(input_fmap_54[47:40]),.by(-9'sd14),.cx(input_fmap_54[55:48]),.cy( 9'sd4),.dx(input_fmap_54[63:56]),.dy(-9'sd7),.chainin(63'd0),.result(O54_N2_S1),.chainout(chainout_2_O54));
logic signed [63:0] chainout_4_O54; 
logic signed [63:0] O54_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O54(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_54[71:64]),.ay(-9'sd9),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O54_N4_S1),.chainout(chainout_4_O54));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O54_N0_S2;		always @(posedge clk) O54_N0_S2 <=     O54_N0_S1  +  O54_N2_S1 ;
 logic signed [21:0] O54_N2_S2;		always @(posedge clk) O54_N2_S2 <=     O54_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O54_N0_S3;		always @(posedge clk) O54_N0_S3 <=     O54_N0_S2  +  O54_N2_S2 ;
 assign conv_mac_54 = O54_N0_S3;

logic signed [31:0] conv_mac_55;
logic signed [63:0] chainout_0_O55; 
logic signed [63:0] O55_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O55(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_55[15:8]),.ay(-9'sd9),.bx(input_fmap_55[23:16]),.by(-9'sd6),.cx(input_fmap_55[31:24]),.cy(-9'sd10),.dx(input_fmap_55[39:32]),.dy(-9'sd13),.chainin(63'd0),.result(O55_N0_S1),.chainout(chainout_0_O55));
logic signed [63:0] chainout_2_O55; 
logic signed [63:0] O55_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O55(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_55[47:40]),.ay( 9'sd2),.bx(input_fmap_55[55:48]),.by( 9'sd1),.cx(input_fmap_55[63:56]),.cy( 9'sd14),.dx(input_fmap_55[71:64]),.dy( 9'sd7),.chainin(63'd0),.result(O55_N2_S1),.chainout(chainout_2_O55));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O55_N0_S2;		always @(posedge clk) O55_N0_S2 <=     O55_N0_S1  +  O55_N2_S1 ;
 assign conv_mac_55 = O55_N0_S2;

logic signed [31:0] conv_mac_56;
logic signed [63:0] chainout_0_O56; 
logic signed [63:0] O56_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O56(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_56[7:0]),.ay( 9'sd5),.bx(input_fmap_56[15:8]),.by( 9'sd11),.cx(input_fmap_56[23:16]),.cy( 9'sd1),.dx(input_fmap_56[31:24]),.dy(-9'sd9),.chainin(63'd0),.result(O56_N0_S1),.chainout(chainout_0_O56));
logic signed [63:0] chainout_2_O56; 
logic signed [63:0] O56_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O56(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_56[39:32]),.ay(-9'sd30),.bx(input_fmap_56[47:40]),.by( 9'sd5),.cx(input_fmap_56[63:56]),.cy(-9'sd6),.dx(input_fmap_56[71:64]),.dy( 9'sd1),.chainin(63'd0),.result(O56_N2_S1),.chainout(chainout_2_O56));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O56_N0_S2;		always @(posedge clk) O56_N0_S2 <=     O56_N0_S1  +  O56_N2_S1 ;
 assign conv_mac_56 = O56_N0_S2;

logic signed [31:0] conv_mac_57;
logic signed [63:0] chainout_0_O57; 
logic signed [63:0] O57_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O57(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_57[7:0]),.ay( 9'sd4),.bx(input_fmap_57[15:8]),.by( 9'sd13),.cx(input_fmap_57[23:16]),.cy(-9'sd2),.dx(input_fmap_57[31:24]),.dy( 9'sd4),.chainin(63'd0),.result(O57_N0_S1),.chainout(chainout_0_O57));
logic signed [63:0] chainout_2_O57; 
logic signed [63:0] O57_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O57(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_57[39:32]),.ay( 9'sd26),.bx(input_fmap_57[47:40]),.by(-9'sd2),.cx(input_fmap_57[55:48]),.cy(-9'sd12),.dx(input_fmap_57[63:56]),.dy(-9'sd22),.chainin(63'd0),.result(O57_N2_S1),.chainout(chainout_2_O57));
logic signed [63:0] chainout_4_O57; 
logic signed [63:0] O57_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O57(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_57[71:64]),.ay(-9'sd9),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O57_N4_S1),.chainout(chainout_4_O57));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O57_N0_S2;		always @(posedge clk) O57_N0_S2 <=     O57_N0_S1  +  O57_N2_S1 ;
 logic signed [21:0] O57_N2_S2;		always @(posedge clk) O57_N2_S2 <=     O57_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O57_N0_S3;		always @(posedge clk) O57_N0_S3 <=     O57_N0_S2  +  O57_N2_S2 ;
 assign conv_mac_57 = O57_N0_S3;

logic signed [31:0] conv_mac_58;
logic signed [63:0] chainout_0_O58; 
logic signed [63:0] O58_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O58(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_58[7:0]),.ay( 9'sd1),.bx(input_fmap_58[15:8]),.by(-9'sd7),.cx(input_fmap_58[23:16]),.cy(-9'sd2),.dx(input_fmap_58[31:24]),.dy( 9'sd1),.chainin(63'd0),.result(O58_N0_S1),.chainout(chainout_0_O58));
logic signed [63:0] chainout_2_O58; 
logic signed [63:0] O58_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O58(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_58[39:32]),.ay(-9'sd23),.bx(input_fmap_58[47:40]),.by( 9'sd9),.cx(input_fmap_58[55:48]),.cy( 9'sd2),.dx(input_fmap_58[63:56]),.dy( 9'sd28),.chainin(63'd0),.result(O58_N2_S1),.chainout(chainout_2_O58));
logic signed [63:0] chainout_4_O58; 
logic signed [63:0] O58_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O58(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_58[71:64]),.ay(-9'sd5),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O58_N4_S1),.chainout(chainout_4_O58));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O58_N0_S2;		always @(posedge clk) O58_N0_S2 <=     O58_N0_S1  +  O58_N2_S1 ;
 logic signed [21:0] O58_N2_S2;		always @(posedge clk) O58_N2_S2 <=     O58_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O58_N0_S3;		always @(posedge clk) O58_N0_S3 <=     O58_N0_S2  +  O58_N2_S2 ;
 assign conv_mac_58 = O58_N0_S3;

logic signed [31:0] conv_mac_59;
logic signed [63:0] chainout_0_O59; 
logic signed [63:0] O59_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O59(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_59[7:0]),.ay(-9'sd3),.bx(input_fmap_59[15:8]),.by(-9'sd8),.cx(input_fmap_59[23:16]),.cy(-9'sd3),.dx(input_fmap_59[31:24]),.dy( 9'sd25),.chainin(63'd0),.result(O59_N0_S1),.chainout(chainout_0_O59));
logic signed [63:0] chainout_2_O59; 
logic signed [63:0] O59_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O59(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_59[39:32]),.ay( 9'sd5),.bx(input_fmap_59[47:40]),.by(-9'sd13),.cx(input_fmap_59[55:48]),.cy(-9'sd2),.dx(input_fmap_59[63:56]),.dy( 9'sd9),.chainin(63'd0),.result(O59_N2_S1),.chainout(chainout_2_O59));
logic signed [63:0] chainout_4_O59; 
logic signed [63:0] O59_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O59(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_59[71:64]),.ay(-9'sd3),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O59_N4_S1),.chainout(chainout_4_O59));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O59_N0_S2;		always @(posedge clk) O59_N0_S2 <=     O59_N0_S1  +  O59_N2_S1 ;
 logic signed [21:0] O59_N2_S2;		always @(posedge clk) O59_N2_S2 <=     O59_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O59_N0_S3;		always @(posedge clk) O59_N0_S3 <=     O59_N0_S2  +  O59_N2_S2 ;
 assign conv_mac_59 = O59_N0_S3;

logic signed [31:0] conv_mac_60;
logic signed [63:0] chainout_0_O60; 
logic signed [63:0] O60_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O60(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_60[7:0]),.ay(-9'sd5),.bx(input_fmap_60[15:8]),.by(-9'sd5),.cx(input_fmap_60[23:16]),.cy( 9'sd6),.dx(input_fmap_60[31:24]),.dy(-9'sd21),.chainin(63'd0),.result(O60_N0_S1),.chainout(chainout_0_O60));
logic signed [63:0] chainout_2_O60; 
logic signed [63:0] O60_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O60(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_60[39:32]),.ay( 9'sd1),.bx(input_fmap_60[47:40]),.by( 9'sd19),.cx(input_fmap_60[55:48]),.cy(-9'sd7),.dx(input_fmap_60[63:56]),.dy( 9'sd6),.chainin(63'd0),.result(O60_N2_S1),.chainout(chainout_2_O60));
logic signed [63:0] chainout_4_O60; 
logic signed [63:0] O60_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O60(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_60[71:64]),.ay( 9'sd3),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O60_N4_S1),.chainout(chainout_4_O60));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O60_N0_S2;		always @(posedge clk) O60_N0_S2 <=     O60_N0_S1  +  O60_N2_S1 ;
 logic signed [21:0] O60_N2_S2;		always @(posedge clk) O60_N2_S2 <=     O60_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O60_N0_S3;		always @(posedge clk) O60_N0_S3 <=     O60_N0_S2  +  O60_N2_S2 ;
 assign conv_mac_60 = O60_N0_S3;

logic signed [31:0] conv_mac_61;
logic signed [63:0] chainout_0_O61; 
logic signed [63:0] O61_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O61(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_61[7:0]),.ay(-9'sd6),.bx(input_fmap_61[15:8]),.by(-9'sd15),.cx(input_fmap_61[23:16]),.cy(-9'sd8),.dx(input_fmap_61[31:24]),.dy(-9'sd3),.chainin(63'd0),.result(O61_N0_S1),.chainout(chainout_0_O61));
logic signed [63:0] chainout_2_O61; 
logic signed [63:0] O61_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O61(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_61[39:32]),.ay( 9'sd56),.bx(input_fmap_61[47:40]),.by( 9'sd4),.cx(input_fmap_61[55:48]),.cy( 9'sd3),.dx(input_fmap_61[63:56]),.dy(-9'sd5),.chainin(63'd0),.result(O61_N2_S1),.chainout(chainout_2_O61));
logic signed [63:0] chainout_4_O61; 
logic signed [63:0] O61_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O61(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_61[71:64]),.ay(-9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O61_N4_S1),.chainout(chainout_4_O61));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O61_N0_S2;		always @(posedge clk) O61_N0_S2 <=     O61_N0_S1  +  O61_N2_S1 ;
 logic signed [21:0] O61_N2_S2;		always @(posedge clk) O61_N2_S2 <=     O61_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O61_N0_S3;		always @(posedge clk) O61_N0_S3 <=     O61_N0_S2  +  O61_N2_S2 ;
 assign conv_mac_61 = O61_N0_S3;

logic signed [31:0] conv_mac_62;
logic signed [63:0] chainout_0_O62; 
logic signed [63:0] O62_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O62(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_62[7:0]),.ay(-9'sd1),.bx(input_fmap_62[15:8]),.by(-9'sd7),.cx(input_fmap_62[23:16]),.cy(-9'sd3),.dx(input_fmap_62[31:24]),.dy( 9'sd2),.chainin(63'd0),.result(O62_N0_S1),.chainout(chainout_0_O62));
logic signed [63:0] chainout_2_O62; 
logic signed [63:0] O62_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O62(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_62[39:32]),.ay( 9'sd25),.bx(input_fmap_62[47:40]),.by( 9'sd5),.cx(input_fmap_62[55:48]),.cy(-9'sd1),.dx(input_fmap_62[63:56]),.dy( 9'sd6),.chainin(63'd0),.result(O62_N2_S1),.chainout(chainout_2_O62));
logic signed [63:0] chainout_4_O62; 
logic signed [63:0] O62_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O62(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_62[71:64]),.ay(-9'sd2),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O62_N4_S1),.chainout(chainout_4_O62));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O62_N0_S2;		always @(posedge clk) O62_N0_S2 <=     O62_N0_S1  +  O62_N2_S1 ;
 logic signed [21:0] O62_N2_S2;		always @(posedge clk) O62_N2_S2 <=     O62_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O62_N0_S3;		always @(posedge clk) O62_N0_S3 <=     O62_N0_S2  +  O62_N2_S2 ;
 assign conv_mac_62 = O62_N0_S3;

logic signed [31:0] conv_mac_63;
logic signed [63:0] chainout_0_O63; 
logic signed [63:0] O63_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O63(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_63[7:0]),.ay( 9'sd10),.bx(input_fmap_63[15:8]),.by( 9'sd33),.cx(input_fmap_63[23:16]),.cy( 9'sd5),.dx(input_fmap_63[31:24]),.dy(-9'sd1),.chainin(63'd0),.result(O63_N0_S1),.chainout(chainout_0_O63));
logic signed [63:0] chainout_2_O63; 
logic signed [63:0] O63_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O63(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_63[39:32]),.ay(-9'sd20),.bx(input_fmap_63[47:40]),.by(-9'sd8),.cx(input_fmap_63[55:48]),.cy(-9'sd9),.dx(input_fmap_63[63:56]),.dy(-9'sd15),.chainin(63'd0),.result(O63_N2_S1),.chainout(chainout_2_O63));
logic signed [63:0] chainout_4_O63; 
logic signed [63:0] O63_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O63(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_63[71:64]),.ay( 9'sd3),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O63_N4_S1),.chainout(chainout_4_O63));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O63_N0_S2;		always @(posedge clk) O63_N0_S2 <=     O63_N0_S1  +  O63_N2_S1 ;
 logic signed [21:0] O63_N2_S2;		always @(posedge clk) O63_N2_S2 <=     O63_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O63_N0_S3;		always @(posedge clk) O63_N0_S3 <=     O63_N0_S2  +  O63_N2_S2 ;
 assign conv_mac_63 = O63_N0_S3;

logic valid_D1;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D1<= 0 ;
	else valid_D1<=valid;
end
logic valid_D2;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D2<= 0 ;
	else valid_D2<=valid_D1;
end
logic valid_D3;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D3<= 0 ;
	else valid_D3<=valid_D2;
end
logic valid_D4;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D4<= 0 ;
	else valid_D4<=valid_D3;
end
always_ff @(posedge clk) begin
	if (rstn == 0) ready <= 0 ;
	else ready <=valid_D4;
end
logic [31:0] bias_add_0;
assign bias_add_0 = conv_mac_0 + 6'd20;
logic [31:0] bias_add_1;
assign bias_add_1 = conv_mac_1 + 4'd5;
logic [31:0] bias_add_2;
assign bias_add_2 = conv_mac_2;
logic [31:0] bias_add_3;
assign bias_add_3 = conv_mac_3 - 5'd8;
logic [31:0] bias_add_4;
assign bias_add_4 = conv_mac_4 + 6'd19;
logic [31:0] bias_add_5;
assign bias_add_5 = conv_mac_5;
logic [31:0] bias_add_6;
assign bias_add_6 = conv_mac_6 + 4'd6;
logic [31:0] bias_add_7;
assign bias_add_7 = conv_mac_7 + 7'd33;
logic [31:0] bias_add_8;
assign bias_add_8 = conv_mac_8 + 6'd17;
logic [31:0] bias_add_9;
assign bias_add_9 = conv_mac_9;
logic [31:0] bias_add_10;
assign bias_add_10 = conv_mac_10 - 4'd6;
logic [31:0] bias_add_11;
assign bias_add_11 = conv_mac_11 + 2'd1;
logic [31:0] bias_add_12;
assign bias_add_12 = conv_mac_12 - 2'd1;
logic [31:0] bias_add_13;
assign bias_add_13 = conv_mac_13 + 6'd20;
logic [31:0] bias_add_14;
assign bias_add_14 = conv_mac_14 + 6'd20;
logic [31:0] bias_add_15;
assign bias_add_15 = conv_mac_15 + 6'd29;
logic [31:0] bias_add_16;
assign bias_add_16 = conv_mac_16;
logic [31:0] bias_add_17;
assign bias_add_17 = conv_mac_17 + 7'd56;
logic [31:0] bias_add_18;
assign bias_add_18 = conv_mac_18 - 4'd5;
logic [31:0] bias_add_19;
assign bias_add_19 = conv_mac_19 + 6'd30;
logic [31:0] bias_add_20;
assign bias_add_20 = conv_mac_20 + 5'd8;
logic [31:0] bias_add_21;
assign bias_add_21 = conv_mac_21 + 4'd7;
logic [31:0] bias_add_22;
assign bias_add_22 = conv_mac_22 + 7'd40;
logic [31:0] bias_add_23;
assign bias_add_23 = conv_mac_23 - 4'd5;
logic [31:0] bias_add_24;
assign bias_add_24 = conv_mac_24 + 5'd13;
logic [31:0] bias_add_25;
assign bias_add_25 = conv_mac_25 - 3'd2;
logic [31:0] bias_add_26;
assign bias_add_26 = conv_mac_26 - 2'd1;
logic [31:0] bias_add_27;
assign bias_add_27 = conv_mac_27 + 7'd43;
logic [31:0] bias_add_28;
assign bias_add_28 = conv_mac_28 - 3'd3;
logic [31:0] bias_add_29;
assign bias_add_29 = conv_mac_29 + 4'd5;
logic [31:0] bias_add_30;
assign bias_add_30 = conv_mac_30 - 3'd2;
logic [31:0] bias_add_31;
assign bias_add_31 = conv_mac_31 + 7'd54;
logic [31:0] bias_add_32;
assign bias_add_32 = conv_mac_32 + 6'd28;
logic [31:0] bias_add_33;
assign bias_add_33 = conv_mac_33 - 3'd2;
logic [31:0] bias_add_34;
assign bias_add_34 = conv_mac_34 - 3'd3;
logic [31:0] bias_add_35;
assign bias_add_35 = conv_mac_35 + 4'd7;
logic [31:0] bias_add_36;
assign bias_add_36 = conv_mac_36;
logic [31:0] bias_add_37;
assign bias_add_37 = conv_mac_37 - 2'd1;
logic [31:0] bias_add_38;
assign bias_add_38 = conv_mac_38 - 4'd4;
logic [31:0] bias_add_39;
assign bias_add_39 = conv_mac_39 - 4'd4;
logic [31:0] bias_add_40;
assign bias_add_40 = conv_mac_40 - 2'd1;
logic [31:0] bias_add_41;
assign bias_add_41 = conv_mac_41 + 6'd31;
logic [31:0] bias_add_42;
assign bias_add_42 = conv_mac_42 + 5'd11;
logic [31:0] bias_add_43;
assign bias_add_43 = conv_mac_43 + 4'd4;
logic [31:0] bias_add_44;
assign bias_add_44 = conv_mac_44 + 6'd28;
logic [31:0] bias_add_45;
assign bias_add_45 = conv_mac_45;
logic [31:0] bias_add_46;
assign bias_add_46 = conv_mac_46 + 6'd20;
logic [31:0] bias_add_47;
assign bias_add_47 = conv_mac_47 + 5'd8;
logic [31:0] bias_add_48;
assign bias_add_48 = conv_mac_48 - 3'd2;
logic [31:0] bias_add_49;
assign bias_add_49 = conv_mac_49 + 5'd9;
logic [31:0] bias_add_50;
assign bias_add_50 = conv_mac_50 + 5'd13;
logic [31:0] bias_add_51;
assign bias_add_51 = conv_mac_51 + 6'd17;
logic [31:0] bias_add_52;
assign bias_add_52 = conv_mac_52 + 5'd10;
logic [31:0] bias_add_53;
assign bias_add_53 = conv_mac_53 - 2'd1;
logic [31:0] bias_add_54;
assign bias_add_54 = conv_mac_54 + 2'd1;
logic [31:0] bias_add_55;
assign bias_add_55 = conv_mac_55 + 6'd20;
logic [31:0] bias_add_56;
assign bias_add_56 = conv_mac_56 + 7'd34;
logic [31:0] bias_add_57;
assign bias_add_57 = conv_mac_57 + 2'd1;
logic [31:0] bias_add_58;
assign bias_add_58 = conv_mac_58 - 3'd3;
logic [31:0] bias_add_59;
assign bias_add_59 = conv_mac_59 - 5'd9;
logic [31:0] bias_add_60;
assign bias_add_60 = conv_mac_60 - 3'd2;
logic [31:0] bias_add_61;
assign bias_add_61 = conv_mac_61 + 6'd23;
logic [31:0] bias_add_62;
assign bias_add_62 = conv_mac_62 - 4'd7;
logic [31:0] bias_add_63;
assign bias_add_63 = conv_mac_63 + 4'd6;

logic [7:0] relu_0;
assign relu_0[7:0] = (bias_add_0[31]==0) ? ((bias_add_0<3'd6) ? {{bias_add_0[31],bias_add_0[10:4]}} :'d6) : '0;
logic [7:0] relu_1;
assign relu_1[7:0] = (bias_add_1[31]==0) ? ((bias_add_1<3'd6) ? {{bias_add_1[31],bias_add_1[10:4]}} :'d6) : '0;
logic [7:0] relu_2;
assign relu_2[7:0] = (bias_add_2[31]==0) ? ((bias_add_2<3'd6) ? {{bias_add_2[31],bias_add_2[10:4]}} :'d6) : '0;
logic [7:0] relu_3;
assign relu_3[7:0] = (bias_add_3[31]==0) ? ((bias_add_3<3'd6) ? {{bias_add_3[31],bias_add_3[10:4]}} :'d6) : '0;
logic [7:0] relu_4;
assign relu_4[7:0] = (bias_add_4[31]==0) ? ((bias_add_4<3'd6) ? {{bias_add_4[31],bias_add_4[10:4]}} :'d6) : '0;
logic [7:0] relu_5;
assign relu_5[7:0] = (bias_add_5[31]==0) ? ((bias_add_5<3'd6) ? {{bias_add_5[31],bias_add_5[10:4]}} :'d6) : '0;
logic [7:0] relu_6;
assign relu_6[7:0] = (bias_add_6[31]==0) ? ((bias_add_6<3'd6) ? {{bias_add_6[31],bias_add_6[10:4]}} :'d6) : '0;
logic [7:0] relu_7;
assign relu_7[7:0] = (bias_add_7[31]==0) ? ((bias_add_7<3'd6) ? {{bias_add_7[31],bias_add_7[10:4]}} :'d6) : '0;
logic [7:0] relu_8;
assign relu_8[7:0] = (bias_add_8[31]==0) ? ((bias_add_8<3'd6) ? {{bias_add_8[31],bias_add_8[10:4]}} :'d6) : '0;
logic [7:0] relu_9;
assign relu_9[7:0] = (bias_add_9[31]==0) ? ((bias_add_9<3'd6) ? {{bias_add_9[31],bias_add_9[10:4]}} :'d6) : '0;
logic [7:0] relu_10;
assign relu_10[7:0] = (bias_add_10[31]==0) ? ((bias_add_10<3'd6) ? {{bias_add_10[31],bias_add_10[10:4]}} :'d6) : '0;
logic [7:0] relu_11;
assign relu_11[7:0] = (bias_add_11[31]==0) ? ((bias_add_11<3'd6) ? {{bias_add_11[31],bias_add_11[10:4]}} :'d6) : '0;
logic [7:0] relu_12;
assign relu_12[7:0] = (bias_add_12[31]==0) ? ((bias_add_12<3'd6) ? {{bias_add_12[31],bias_add_12[10:4]}} :'d6) : '0;
logic [7:0] relu_13;
assign relu_13[7:0] = (bias_add_13[31]==0) ? ((bias_add_13<3'd6) ? {{bias_add_13[31],bias_add_13[10:4]}} :'d6) : '0;
logic [7:0] relu_14;
assign relu_14[7:0] = (bias_add_14[31]==0) ? ((bias_add_14<3'd6) ? {{bias_add_14[31],bias_add_14[10:4]}} :'d6) : '0;
logic [7:0] relu_15;
assign relu_15[7:0] = (bias_add_15[31]==0) ? ((bias_add_15<3'd6) ? {{bias_add_15[31],bias_add_15[10:4]}} :'d6) : '0;
logic [7:0] relu_16;
assign relu_16[7:0] = (bias_add_16[31]==0) ? ((bias_add_16<3'd6) ? {{bias_add_16[31],bias_add_16[10:4]}} :'d6) : '0;
logic [7:0] relu_17;
assign relu_17[7:0] = (bias_add_17[31]==0) ? ((bias_add_17<3'd6) ? {{bias_add_17[31],bias_add_17[10:4]}} :'d6) : '0;
logic [7:0] relu_18;
assign relu_18[7:0] = (bias_add_18[31]==0) ? ((bias_add_18<3'd6) ? {{bias_add_18[31],bias_add_18[10:4]}} :'d6) : '0;
logic [7:0] relu_19;
assign relu_19[7:0] = (bias_add_19[31]==0) ? ((bias_add_19<3'd6) ? {{bias_add_19[31],bias_add_19[10:4]}} :'d6) : '0;
logic [7:0] relu_20;
assign relu_20[7:0] = (bias_add_20[31]==0) ? ((bias_add_20<3'd6) ? {{bias_add_20[31],bias_add_20[10:4]}} :'d6) : '0;
logic [7:0] relu_21;
assign relu_21[7:0] = (bias_add_21[31]==0) ? ((bias_add_21<3'd6) ? {{bias_add_21[31],bias_add_21[10:4]}} :'d6) : '0;
logic [7:0] relu_22;
assign relu_22[7:0] = (bias_add_22[31]==0) ? ((bias_add_22<3'd6) ? {{bias_add_22[31],bias_add_22[10:4]}} :'d6) : '0;
logic [7:0] relu_23;
assign relu_23[7:0] = (bias_add_23[31]==0) ? ((bias_add_23<3'd6) ? {{bias_add_23[31],bias_add_23[10:4]}} :'d6) : '0;
logic [7:0] relu_24;
assign relu_24[7:0] = (bias_add_24[31]==0) ? ((bias_add_24<3'd6) ? {{bias_add_24[31],bias_add_24[10:4]}} :'d6) : '0;
logic [7:0] relu_25;
assign relu_25[7:0] = (bias_add_25[31]==0) ? ((bias_add_25<3'd6) ? {{bias_add_25[31],bias_add_25[10:4]}} :'d6) : '0;
logic [7:0] relu_26;
assign relu_26[7:0] = (bias_add_26[31]==0) ? ((bias_add_26<3'd6) ? {{bias_add_26[31],bias_add_26[10:4]}} :'d6) : '0;
logic [7:0] relu_27;
assign relu_27[7:0] = (bias_add_27[31]==0) ? ((bias_add_27<3'd6) ? {{bias_add_27[31],bias_add_27[10:4]}} :'d6) : '0;
logic [7:0] relu_28;
assign relu_28[7:0] = (bias_add_28[31]==0) ? ((bias_add_28<3'd6) ? {{bias_add_28[31],bias_add_28[10:4]}} :'d6) : '0;
logic [7:0] relu_29;
assign relu_29[7:0] = (bias_add_29[31]==0) ? ((bias_add_29<3'd6) ? {{bias_add_29[31],bias_add_29[10:4]}} :'d6) : '0;
logic [7:0] relu_30;
assign relu_30[7:0] = (bias_add_30[31]==0) ? ((bias_add_30<3'd6) ? {{bias_add_30[31],bias_add_30[10:4]}} :'d6) : '0;
logic [7:0] relu_31;
assign relu_31[7:0] = (bias_add_31[31]==0) ? ((bias_add_31<3'd6) ? {{bias_add_31[31],bias_add_31[10:4]}} :'d6) : '0;
logic [7:0] relu_32;
assign relu_32[7:0] = (bias_add_32[31]==0) ? ((bias_add_32<3'd6) ? {{bias_add_32[31],bias_add_32[10:4]}} :'d6) : '0;
logic [7:0] relu_33;
assign relu_33[7:0] = (bias_add_33[31]==0) ? ((bias_add_33<3'd6) ? {{bias_add_33[31],bias_add_33[10:4]}} :'d6) : '0;
logic [7:0] relu_34;
assign relu_34[7:0] = (bias_add_34[31]==0) ? ((bias_add_34<3'd6) ? {{bias_add_34[31],bias_add_34[10:4]}} :'d6) : '0;
logic [7:0] relu_35;
assign relu_35[7:0] = (bias_add_35[31]==0) ? ((bias_add_35<3'd6) ? {{bias_add_35[31],bias_add_35[10:4]}} :'d6) : '0;
logic [7:0] relu_36;
assign relu_36[7:0] = (bias_add_36[31]==0) ? ((bias_add_36<3'd6) ? {{bias_add_36[31],bias_add_36[10:4]}} :'d6) : '0;
logic [7:0] relu_37;
assign relu_37[7:0] = (bias_add_37[31]==0) ? ((bias_add_37<3'd6) ? {{bias_add_37[31],bias_add_37[10:4]}} :'d6) : '0;
logic [7:0] relu_38;
assign relu_38[7:0] = (bias_add_38[31]==0) ? ((bias_add_38<3'd6) ? {{bias_add_38[31],bias_add_38[10:4]}} :'d6) : '0;
logic [7:0] relu_39;
assign relu_39[7:0] = (bias_add_39[31]==0) ? ((bias_add_39<3'd6) ? {{bias_add_39[31],bias_add_39[10:4]}} :'d6) : '0;
logic [7:0] relu_40;
assign relu_40[7:0] = (bias_add_40[31]==0) ? ((bias_add_40<3'd6) ? {{bias_add_40[31],bias_add_40[10:4]}} :'d6) : '0;
logic [7:0] relu_41;
assign relu_41[7:0] = (bias_add_41[31]==0) ? ((bias_add_41<3'd6) ? {{bias_add_41[31],bias_add_41[10:4]}} :'d6) : '0;
logic [7:0] relu_42;
assign relu_42[7:0] = (bias_add_42[31]==0) ? ((bias_add_42<3'd6) ? {{bias_add_42[31],bias_add_42[10:4]}} :'d6) : '0;
logic [7:0] relu_43;
assign relu_43[7:0] = (bias_add_43[31]==0) ? ((bias_add_43<3'd6) ? {{bias_add_43[31],bias_add_43[10:4]}} :'d6) : '0;
logic [7:0] relu_44;
assign relu_44[7:0] = (bias_add_44[31]==0) ? ((bias_add_44<3'd6) ? {{bias_add_44[31],bias_add_44[10:4]}} :'d6) : '0;
logic [7:0] relu_45;
assign relu_45[7:0] = (bias_add_45[31]==0) ? ((bias_add_45<3'd6) ? {{bias_add_45[31],bias_add_45[10:4]}} :'d6) : '0;
logic [7:0] relu_46;
assign relu_46[7:0] = (bias_add_46[31]==0) ? ((bias_add_46<3'd6) ? {{bias_add_46[31],bias_add_46[10:4]}} :'d6) : '0;
logic [7:0] relu_47;
assign relu_47[7:0] = (bias_add_47[31]==0) ? ((bias_add_47<3'd6) ? {{bias_add_47[31],bias_add_47[10:4]}} :'d6) : '0;
logic [7:0] relu_48;
assign relu_48[7:0] = (bias_add_48[31]==0) ? ((bias_add_48<3'd6) ? {{bias_add_48[31],bias_add_48[10:4]}} :'d6) : '0;
logic [7:0] relu_49;
assign relu_49[7:0] = (bias_add_49[31]==0) ? ((bias_add_49<3'd6) ? {{bias_add_49[31],bias_add_49[10:4]}} :'d6) : '0;
logic [7:0] relu_50;
assign relu_50[7:0] = (bias_add_50[31]==0) ? ((bias_add_50<3'd6) ? {{bias_add_50[31],bias_add_50[10:4]}} :'d6) : '0;
logic [7:0] relu_51;
assign relu_51[7:0] = (bias_add_51[31]==0) ? ((bias_add_51<3'd6) ? {{bias_add_51[31],bias_add_51[10:4]}} :'d6) : '0;
logic [7:0] relu_52;
assign relu_52[7:0] = (bias_add_52[31]==0) ? ((bias_add_52<3'd6) ? {{bias_add_52[31],bias_add_52[10:4]}} :'d6) : '0;
logic [7:0] relu_53;
assign relu_53[7:0] = (bias_add_53[31]==0) ? ((bias_add_53<3'd6) ? {{bias_add_53[31],bias_add_53[10:4]}} :'d6) : '0;
logic [7:0] relu_54;
assign relu_54[7:0] = (bias_add_54[31]==0) ? ((bias_add_54<3'd6) ? {{bias_add_54[31],bias_add_54[10:4]}} :'d6) : '0;
logic [7:0] relu_55;
assign relu_55[7:0] = (bias_add_55[31]==0) ? ((bias_add_55<3'd6) ? {{bias_add_55[31],bias_add_55[10:4]}} :'d6) : '0;
logic [7:0] relu_56;
assign relu_56[7:0] = (bias_add_56[31]==0) ? ((bias_add_56<3'd6) ? {{bias_add_56[31],bias_add_56[10:4]}} :'d6) : '0;
logic [7:0] relu_57;
assign relu_57[7:0] = (bias_add_57[31]==0) ? ((bias_add_57<3'd6) ? {{bias_add_57[31],bias_add_57[10:4]}} :'d6) : '0;
logic [7:0] relu_58;
assign relu_58[7:0] = (bias_add_58[31]==0) ? ((bias_add_58<3'd6) ? {{bias_add_58[31],bias_add_58[10:4]}} :'d6) : '0;
logic [7:0] relu_59;
assign relu_59[7:0] = (bias_add_59[31]==0) ? ((bias_add_59<3'd6) ? {{bias_add_59[31],bias_add_59[10:4]}} :'d6) : '0;
logic [7:0] relu_60;
assign relu_60[7:0] = (bias_add_60[31]==0) ? ((bias_add_60<3'd6) ? {{bias_add_60[31],bias_add_60[10:4]}} :'d6) : '0;
logic [7:0] relu_61;
assign relu_61[7:0] = (bias_add_61[31]==0) ? ((bias_add_61<3'd6) ? {{bias_add_61[31],bias_add_61[10:4]}} :'d6) : '0;
logic [7:0] relu_62;
assign relu_62[7:0] = (bias_add_62[31]==0) ? ((bias_add_62<3'd6) ? {{bias_add_62[31],bias_add_62[10:4]}} :'d6) : '0;
logic [7:0] relu_63;
assign relu_63[7:0] = (bias_add_63[31]==0) ? ((bias_add_63<3'd6) ? {{bias_add_63[31],bias_add_63[10:4]}} :'d6) : '0;

assign output_act = {
	relu_63,
	relu_62,
	relu_61,
	relu_60,
	relu_59,
	relu_58,
	relu_57,
	relu_56,
	relu_55,
	relu_54,
	relu_53,
	relu_52,
	relu_51,
	relu_50,
	relu_49,
	relu_48,
	relu_47,
	relu_46,
	relu_45,
	relu_44,
	relu_43,
	relu_42,
	relu_41,
	relu_40,
	relu_39,
	relu_38,
	relu_37,
	relu_36,
	relu_35,
	relu_34,
	relu_33,
	relu_32,
	relu_31,
	relu_30,
	relu_29,
	relu_28,
	relu_27,
	relu_26,
	relu_25,
	relu_24,
	relu_23,
	relu_22,
	relu_21,
	relu_20,
	relu_19,
	relu_18,
	relu_17,
	relu_16,
	relu_15,
	relu_14,
	relu_13,
	relu_12,
	relu_11,
	relu_10,
	relu_9,
	relu_8,
	relu_7,
	relu_6,
	relu_5,
	relu_4,
	relu_3,
	relu_2,
	relu_1,
	relu_0
};

endmodule
module conv8_dw (
    input logic clk,
    input logic rstn,
    input logic valid,
    input logic [64*72-1:0] input_act,
    output logic [512-1:0] output_act,
    output logic ready
);
logic we;
logic [8:0] zero_number; 
assign zero_number = 9'd0; 
logic [64*72-1:0] input_act_ff;
genvar i;
generate
for (i=0;i<64;i++)
    begin: genblk_13
        always_ff @(posedge clk) begin
            if (rstn == 0) begin
                input_act_ff[(i+1)*72-1:i*72] <= '0;
            end
            else begin
                input_act_ff[(i+1)*72-1:i*72] <= input_act[(i+1)*72-1:i*72];
            end
        end
    end
endgenerate
logic [71:0] input_fmap_0;
assign input_fmap_0 = input_act_ff[71:0];
logic [71:0] input_fmap_1;
assign input_fmap_1 = input_act_ff[143:72];
logic [71:0] input_fmap_2;
assign input_fmap_2 = input_act_ff[215:144];
logic [71:0] input_fmap_3;
assign input_fmap_3 = input_act_ff[287:216];
logic [71:0] input_fmap_4;
assign input_fmap_4 = input_act_ff[359:288];
logic [71:0] input_fmap_5;
assign input_fmap_5 = input_act_ff[431:360];
logic [71:0] input_fmap_6;
assign input_fmap_6 = input_act_ff[503:432];
logic [71:0] input_fmap_7;
assign input_fmap_7 = input_act_ff[575:504];
logic [71:0] input_fmap_8;
assign input_fmap_8 = input_act_ff[647:576];
logic [71:0] input_fmap_9;
assign input_fmap_9 = input_act_ff[719:648];
logic [71:0] input_fmap_10;
assign input_fmap_10 = input_act_ff[791:720];
logic [71:0] input_fmap_11;
assign input_fmap_11 = input_act_ff[863:792];
logic [71:0] input_fmap_12;
assign input_fmap_12 = input_act_ff[935:864];
logic [71:0] input_fmap_13;
assign input_fmap_13 = input_act_ff[1007:936];
logic [71:0] input_fmap_14;
assign input_fmap_14 = input_act_ff[1079:1008];
logic [71:0] input_fmap_15;
assign input_fmap_15 = input_act_ff[1151:1080];
logic [71:0] input_fmap_16;
assign input_fmap_16 = input_act_ff[1223:1152];
logic [71:0] input_fmap_17;
assign input_fmap_17 = input_act_ff[1295:1224];
logic [71:0] input_fmap_18;
assign input_fmap_18 = input_act_ff[1367:1296];
logic [71:0] input_fmap_19;
assign input_fmap_19 = input_act_ff[1439:1368];
logic [71:0] input_fmap_20;
assign input_fmap_20 = input_act_ff[1511:1440];
logic [71:0] input_fmap_21;
assign input_fmap_21 = input_act_ff[1583:1512];
logic [71:0] input_fmap_22;
assign input_fmap_22 = input_act_ff[1655:1584];
logic [71:0] input_fmap_23;
assign input_fmap_23 = input_act_ff[1727:1656];
logic [71:0] input_fmap_24;
assign input_fmap_24 = input_act_ff[1799:1728];
logic [71:0] input_fmap_25;
assign input_fmap_25 = input_act_ff[1871:1800];
logic [71:0] input_fmap_26;
assign input_fmap_26 = input_act_ff[1943:1872];
logic [71:0] input_fmap_27;
assign input_fmap_27 = input_act_ff[2015:1944];
logic [71:0] input_fmap_28;
assign input_fmap_28 = input_act_ff[2087:2016];
logic [71:0] input_fmap_29;
assign input_fmap_29 = input_act_ff[2159:2088];
logic [71:0] input_fmap_30;
assign input_fmap_30 = input_act_ff[2231:2160];
logic [71:0] input_fmap_31;
assign input_fmap_31 = input_act_ff[2303:2232];
logic [71:0] input_fmap_32;
assign input_fmap_32 = input_act_ff[2375:2304];
logic [71:0] input_fmap_33;
assign input_fmap_33 = input_act_ff[2447:2376];
logic [71:0] input_fmap_34;
assign input_fmap_34 = input_act_ff[2519:2448];
logic [71:0] input_fmap_35;
assign input_fmap_35 = input_act_ff[2591:2520];
logic [71:0] input_fmap_36;
assign input_fmap_36 = input_act_ff[2663:2592];
logic [71:0] input_fmap_37;
assign input_fmap_37 = input_act_ff[2735:2664];
logic [71:0] input_fmap_38;
assign input_fmap_38 = input_act_ff[2807:2736];
logic [71:0] input_fmap_39;
assign input_fmap_39 = input_act_ff[2879:2808];
logic [71:0] input_fmap_40;
assign input_fmap_40 = input_act_ff[2951:2880];
logic [71:0] input_fmap_41;
assign input_fmap_41 = input_act_ff[3023:2952];
logic [71:0] input_fmap_42;
assign input_fmap_42 = input_act_ff[3095:3024];
logic [71:0] input_fmap_43;
assign input_fmap_43 = input_act_ff[3167:3096];
logic [71:0] input_fmap_44;
assign input_fmap_44 = input_act_ff[3239:3168];
logic [71:0] input_fmap_45;
assign input_fmap_45 = input_act_ff[3311:3240];
logic [71:0] input_fmap_46;
assign input_fmap_46 = input_act_ff[3383:3312];
logic [71:0] input_fmap_47;
assign input_fmap_47 = input_act_ff[3455:3384];
logic [71:0] input_fmap_48;
assign input_fmap_48 = input_act_ff[3527:3456];
logic [71:0] input_fmap_49;
assign input_fmap_49 = input_act_ff[3599:3528];
logic [71:0] input_fmap_50;
assign input_fmap_50 = input_act_ff[3671:3600];
logic [71:0] input_fmap_51;
assign input_fmap_51 = input_act_ff[3743:3672];
logic [71:0] input_fmap_52;
assign input_fmap_52 = input_act_ff[3815:3744];
logic [71:0] input_fmap_53;
assign input_fmap_53 = input_act_ff[3887:3816];
logic [71:0] input_fmap_54;
assign input_fmap_54 = input_act_ff[3959:3888];
logic [71:0] input_fmap_55;
assign input_fmap_55 = input_act_ff[4031:3960];
logic [71:0] input_fmap_56;
assign input_fmap_56 = input_act_ff[4103:4032];
logic [71:0] input_fmap_57;
assign input_fmap_57 = input_act_ff[4175:4104];
logic [71:0] input_fmap_58;
assign input_fmap_58 = input_act_ff[4247:4176];
logic [71:0] input_fmap_59;
assign input_fmap_59 = input_act_ff[4319:4248];
logic [71:0] input_fmap_60;
assign input_fmap_60 = input_act_ff[4391:4320];
logic [71:0] input_fmap_61;
assign input_fmap_61 = input_act_ff[4463:4392];
logic [71:0] input_fmap_62;
assign input_fmap_62 = input_act_ff[4535:4464];
logic [71:0] input_fmap_63;
assign input_fmap_63 = input_act_ff[4607:4536];

logic signed [31:0] conv_mac_0;
logic signed [63:0] chainout_0_O0; 
logic signed [63:0] O0_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O0(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd4),.bx(input_fmap_0[15:8]),.by(-9'sd9),.cx(input_fmap_0[23:16]),.cy(-9'sd6),.dx(input_fmap_0[39:32]),.dy(-9'sd16),.chainin(63'd0),.result(O0_N0_S1),.chainout(chainout_0_O0));
logic signed [63:0] chainout_2_O0; 
logic signed [63:0] O0_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O0(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[47:40]),.ay(-9'sd7),.bx(input_fmap_0[55:48]),.by( 9'sd13),.cx(input_fmap_0[63:56]),.cy( 9'sd4),.dx(input_fmap_0[71:64]),.dy( 9'sd1),.chainin(63'd0),.result(O0_N2_S1),.chainout(chainout_2_O0));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O0_N0_S2;		always @(posedge clk) O0_N0_S2 <=     O0_N0_S1  +  O0_N2_S1 ;
 assign conv_mac_0 = O0_N0_S2;

logic signed [31:0] conv_mac_1;
logic signed [63:0] chainout_0_O1; 
logic signed [63:0] O1_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O1(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay( 9'sd4),.bx(input_fmap_1[15:8]),.by( 9'sd16),.cx(input_fmap_1[23:16]),.cy( 9'sd2),.dx(input_fmap_1[31:24]),.dy( 9'sd12),.chainin(63'd0),.result(O1_N0_S1),.chainout(chainout_0_O1));
logic signed [63:0] chainout_2_O1; 
logic signed [63:0] O1_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O1(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[39:32]),.ay( 9'sd13),.bx(input_fmap_1[47:40]),.by(-9'sd5),.cx(input_fmap_1[55:48]),.cy(-9'sd6),.dx(input_fmap_1[63:56]),.dy(-9'sd11),.chainin(63'd0),.result(O1_N2_S1),.chainout(chainout_2_O1));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O1_N0_S2;		always @(posedge clk) O1_N0_S2 <=     O1_N0_S1  +  O1_N2_S1 ;
 assign conv_mac_1 = O1_N0_S2;

logic signed [31:0] conv_mac_2;
logic signed [63:0] chainout_0_O2; 
logic signed [63:0] O2_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O2(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_2[7:0]),.ay( 9'sd3),.bx(input_fmap_2[15:8]),.by(-9'sd7),.cx(input_fmap_2[23:16]),.cy( 9'sd3),.dx(input_fmap_2[31:24]),.dy(-9'sd1),.chainin(63'd0),.result(O2_N0_S1),.chainout(chainout_0_O2));
logic signed [63:0] chainout_2_O2; 
logic signed [63:0] O2_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O2(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_2[39:32]),.ay(-9'sd29),.bx(input_fmap_2[47:40]),.by( 9'sd2),.cx(input_fmap_2[55:48]),.cy( 9'sd3),.dx(input_fmap_2[63:56]),.dy(-9'sd5),.chainin(63'd0),.result(O2_N2_S1),.chainout(chainout_2_O2));
logic signed [63:0] chainout_4_O2; 
logic signed [63:0] O2_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O2(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_2[71:64]),.ay( 9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O2_N4_S1),.chainout(chainout_4_O2));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O2_N0_S2;		always @(posedge clk) O2_N0_S2 <=     O2_N0_S1  +  O2_N2_S1 ;
 logic signed [21:0] O2_N2_S2;		always @(posedge clk) O2_N2_S2 <=     O2_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O2_N0_S3;		always @(posedge clk) O2_N0_S3 <=     O2_N0_S2  +  O2_N2_S2 ;
 assign conv_mac_2 = O2_N0_S3;

logic signed [31:0] conv_mac_3;
logic signed [63:0] chainout_0_O3; 
logic signed [63:0] O3_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O3(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_3[7:0]),.ay( 9'sd3),.bx(input_fmap_3[15:8]),.by( 9'sd10),.cx(input_fmap_3[23:16]),.cy( 9'sd7),.dx(input_fmap_3[31:24]),.dy( 9'sd2),.chainin(63'd0),.result(O3_N0_S1),.chainout(chainout_0_O3));
logic signed [63:0] chainout_2_O3; 
logic signed [63:0] O3_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O3(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_3[39:32]),.ay( 9'sd11),.bx(input_fmap_3[47:40]),.by(-9'sd1),.cx(input_fmap_3[55:48]),.cy(-9'sd5),.dx(input_fmap_3[63:56]),.dy(-9'sd21),.chainin(63'd0),.result(O3_N2_S1),.chainout(chainout_2_O3));
logic signed [63:0] chainout_4_O3; 
logic signed [63:0] O3_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O3(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_3[71:64]),.ay(-9'sd7),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O3_N4_S1),.chainout(chainout_4_O3));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O3_N0_S2;		always @(posedge clk) O3_N0_S2 <=     O3_N0_S1  +  O3_N2_S1 ;
 logic signed [21:0] O3_N2_S2;		always @(posedge clk) O3_N2_S2 <=     O3_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O3_N0_S3;		always @(posedge clk) O3_N0_S3 <=     O3_N0_S2  +  O3_N2_S2 ;
 assign conv_mac_3 = O3_N0_S3;

logic signed [31:0] conv_mac_4;
logic signed [63:0] chainout_0_O4; 
logic signed [63:0] O4_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O4(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_4[7:0]),.ay(-9'sd8),.bx(input_fmap_4[15:8]),.by(-9'sd7),.cx(input_fmap_4[23:16]),.cy(-9'sd6),.dx(input_fmap_4[31:24]),.dy(-9'sd6),.chainin(63'd0),.result(O4_N0_S1),.chainout(chainout_0_O4));
logic signed [63:0] chainout_2_O4; 
logic signed [63:0] O4_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O4(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_4[39:32]),.ay(-9'sd17),.bx(input_fmap_4[47:40]),.by(-9'sd4),.cx(input_fmap_4[55:48]),.cy( 9'sd4),.dx(input_fmap_4[63:56]),.dy( 9'sd13),.chainin(63'd0),.result(O4_N2_S1),.chainout(chainout_2_O4));
logic signed [63:0] chainout_4_O4; 
logic signed [63:0] O4_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O4(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_4[71:64]),.ay( 9'sd7),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O4_N4_S1),.chainout(chainout_4_O4));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O4_N0_S2;		always @(posedge clk) O4_N0_S2 <=     O4_N0_S1  +  O4_N2_S1 ;
 logic signed [21:0] O4_N2_S2;		always @(posedge clk) O4_N2_S2 <=     O4_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O4_N0_S3;		always @(posedge clk) O4_N0_S3 <=     O4_N0_S2  +  O4_N2_S2 ;
 assign conv_mac_4 = O4_N0_S3;

logic signed [31:0] conv_mac_5;
logic signed [63:0] chainout_0_O5; 
logic signed [63:0] O5_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O5(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_5[7:0]),.ay(-9'sd2),.bx(input_fmap_5[15:8]),.by( 9'sd2),.cx(input_fmap_5[23:16]),.cy( 9'sd3),.dx(input_fmap_5[31:24]),.dy(-9'sd7),.chainin(63'd0),.result(O5_N0_S1),.chainout(chainout_0_O5));
logic signed [63:0] chainout_2_O5; 
logic signed [63:0] O5_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O5(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_5[39:32]),.ay( 9'sd39),.bx(input_fmap_5[47:40]),.by(-9'sd2),.cx(input_fmap_5[55:48]),.cy(-9'sd4),.dx(input_fmap_5[63:56]),.dy(-9'sd17),.chainin(63'd0),.result(O5_N2_S1),.chainout(chainout_2_O5));
logic signed [63:0] chainout_4_O5; 
logic signed [63:0] O5_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O5(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_5[71:64]),.ay(-9'sd3),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O5_N4_S1),.chainout(chainout_4_O5));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O5_N0_S2;		always @(posedge clk) O5_N0_S2 <=     O5_N0_S1  +  O5_N2_S1 ;
 logic signed [21:0] O5_N2_S2;		always @(posedge clk) O5_N2_S2 <=     O5_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O5_N0_S3;		always @(posedge clk) O5_N0_S3 <=     O5_N0_S2  +  O5_N2_S2 ;
 assign conv_mac_5 = O5_N0_S3;

logic signed [31:0] conv_mac_6;
logic signed [63:0] chainout_0_O6; 
logic signed [63:0] O6_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O6(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_6[7:0]),.ay( 9'sd16),.bx(input_fmap_6[15:8]),.by( 9'sd3),.cx(input_fmap_6[23:16]),.cy(-9'sd13),.dx(input_fmap_6[31:24]),.dy(-9'sd4),.chainin(63'd0),.result(O6_N0_S1),.chainout(chainout_0_O6));
logic signed [63:0] chainout_2_O6; 
logic signed [63:0] O6_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O6(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_6[39:32]),.ay(-9'sd5),.bx(input_fmap_6[47:40]),.by( 9'sd8),.cx(input_fmap_6[55:48]),.cy(-9'sd9),.dx(input_fmap_6[63:56]),.dy( 9'sd2),.chainin(63'd0),.result(O6_N2_S1),.chainout(chainout_2_O6));
logic signed [63:0] chainout_4_O6; 
logic signed [63:0] O6_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O6(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_6[71:64]),.ay( 9'sd14),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O6_N4_S1),.chainout(chainout_4_O6));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O6_N0_S2;		always @(posedge clk) O6_N0_S2 <=     O6_N0_S1  +  O6_N2_S1 ;
 logic signed [21:0] O6_N2_S2;		always @(posedge clk) O6_N2_S2 <=     O6_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O6_N0_S3;		always @(posedge clk) O6_N0_S3 <=     O6_N0_S2  +  O6_N2_S2 ;
 assign conv_mac_6 = O6_N0_S3;

logic signed [31:0] conv_mac_7;
logic signed [63:0] chainout_0_O7; 
logic signed [63:0] O7_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O7(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_7[7:0]),.ay(-9'sd5),.bx(input_fmap_7[15:8]),.by(-9'sd7),.cx(input_fmap_7[23:16]),.cy(-9'sd5),.dx(input_fmap_7[31:24]),.dy(-9'sd4),.chainin(63'd0),.result(O7_N0_S1),.chainout(chainout_0_O7));
logic signed [63:0] chainout_2_O7; 
logic signed [63:0] O7_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O7(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_7[39:32]),.ay(-9'sd14),.bx(input_fmap_7[47:40]),.by(-9'sd4),.cx(input_fmap_7[55:48]),.cy( 9'sd3),.dx(input_fmap_7[63:56]),.dy(-9'sd1),.chainin(63'd0),.result(O7_N2_S1),.chainout(chainout_2_O7));
logic signed [63:0] chainout_4_O7; 
logic signed [63:0] O7_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O7(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_7[71:64]),.ay(-9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O7_N4_S1),.chainout(chainout_4_O7));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O7_N0_S2;		always @(posedge clk) O7_N0_S2 <=     O7_N0_S1  +  O7_N2_S1 ;
 logic signed [21:0] O7_N2_S2;		always @(posedge clk) O7_N2_S2 <=     O7_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O7_N0_S3;		always @(posedge clk) O7_N0_S3 <=     O7_N0_S2  +  O7_N2_S2 ;
 assign conv_mac_7 = O7_N0_S3;

logic signed [31:0] conv_mac_8;
logic signed [63:0] chainout_0_O8; 
logic signed [63:0] O8_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O8(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_8[7:0]),.ay(-9'sd3),.bx(input_fmap_8[15:8]),.by( 9'sd4),.cx(input_fmap_8[31:24]),.cy(-9'sd10),.dx(input_fmap_8[39:32]),.dy(-9'sd14),.chainin(63'd0),.result(O8_N0_S1),.chainout(chainout_0_O8));
logic signed [63:0] chainout_2_O8; 
logic signed [63:0] O8_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O8(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_8[47:40]),.ay(-9'sd12),.bx(input_fmap_8[55:48]),.by(-9'sd2),.cx(input_fmap_8[63:56]),.cy( 9'sd3),.dx(input_fmap_8[71:64]),.dy(-9'sd3),.chainin(63'd0),.result(O8_N2_S1),.chainout(chainout_2_O8));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O8_N0_S2;		always @(posedge clk) O8_N0_S2 <=     O8_N0_S1  +  O8_N2_S1 ;
 assign conv_mac_8 = O8_N0_S2;

logic signed [31:0] conv_mac_9;
logic signed [63:0] chainout_0_O9; 
logic signed [63:0] O9_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O9(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_9[7:0]),.ay(-9'sd6),.bx(input_fmap_9[15:8]),.by( 9'sd10),.cx(input_fmap_9[23:16]),.cy( 9'sd9),.dx(input_fmap_9[31:24]),.dy(-9'sd16),.chainin(63'd0),.result(O9_N0_S1),.chainout(chainout_0_O9));
logic signed [63:0] chainout_2_O9; 
logic signed [63:0] O9_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O9(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_9[39:32]),.ay( 9'sd27),.bx(input_fmap_9[47:40]),.by( 9'sd6),.cx(input_fmap_9[55:48]),.cy(-9'sd1),.dx(input_fmap_9[63:56]),.dy(-9'sd25),.chainin(63'd0),.result(O9_N2_S1),.chainout(chainout_2_O9));
logic signed [63:0] chainout_4_O9; 
logic signed [63:0] O9_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O9(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_9[71:64]),.ay(-9'sd10),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O9_N4_S1),.chainout(chainout_4_O9));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O9_N0_S2;		always @(posedge clk) O9_N0_S2 <=     O9_N0_S1  +  O9_N2_S1 ;
 logic signed [21:0] O9_N2_S2;		always @(posedge clk) O9_N2_S2 <=     O9_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O9_N0_S3;		always @(posedge clk) O9_N0_S3 <=     O9_N0_S2  +  O9_N2_S2 ;
 assign conv_mac_9 = O9_N0_S3;

logic signed [31:0] conv_mac_10;
logic signed [63:0] chainout_0_O10; 
logic signed [63:0] O10_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O10(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_10[7:0]),.ay( 9'sd2),.bx(input_fmap_10[15:8]),.by( 9'sd9),.cx(input_fmap_10[23:16]),.cy( 9'sd2),.dx(input_fmap_10[31:24]),.dy( 9'sd3),.chainin(63'd0),.result(O10_N0_S1),.chainout(chainout_0_O10));
logic signed [63:0] chainout_2_O10; 
logic signed [63:0] O10_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O10(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_10[39:32]),.ay( 9'sd17),.bx(input_fmap_10[47:40]),.by( 9'sd7),.cx(input_fmap_10[55:48]),.cy(-9'sd3),.dx(input_fmap_10[63:56]),.dy(-9'sd5),.chainin(63'd0),.result(O10_N2_S1),.chainout(chainout_2_O10));
logic signed [63:0] chainout_4_O10; 
logic signed [63:0] O10_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O10(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_10[71:64]),.ay(-9'sd2),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O10_N4_S1),.chainout(chainout_4_O10));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O10_N0_S2;		always @(posedge clk) O10_N0_S2 <=     O10_N0_S1  +  O10_N2_S1 ;
 logic signed [21:0] O10_N2_S2;		always @(posedge clk) O10_N2_S2 <=     O10_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O10_N0_S3;		always @(posedge clk) O10_N0_S3 <=     O10_N0_S2  +  O10_N2_S2 ;
 assign conv_mac_10 = O10_N0_S3;

logic signed [31:0] conv_mac_11;
logic signed [63:0] chainout_0_O11; 
logic signed [63:0] O11_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O11(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_11[7:0]),.ay( 9'sd1),.bx(input_fmap_11[15:8]),.by(-9'sd17),.cx(input_fmap_11[23:16]),.cy(-9'sd7),.dx(input_fmap_11[31:24]),.dy(-9'sd1),.chainin(63'd0),.result(O11_N0_S1),.chainout(chainout_0_O11));
logic signed [63:0] chainout_2_O11; 
logic signed [63:0] O11_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O11(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_11[39:32]),.ay( 9'sd26),.bx(input_fmap_11[47:40]),.by(-9'sd4),.cx(input_fmap_11[55:48]),.cy(-9'sd2),.dx(input_fmap_11[63:56]),.dy( 9'sd3),.chainin(63'd0),.result(O11_N2_S1),.chainout(chainout_2_O11));
logic signed [63:0] chainout_4_O11; 
logic signed [63:0] O11_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O11(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_11[71:64]),.ay( 9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O11_N4_S1),.chainout(chainout_4_O11));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O11_N0_S2;		always @(posedge clk) O11_N0_S2 <=     O11_N0_S1  +  O11_N2_S1 ;
 logic signed [21:0] O11_N2_S2;		always @(posedge clk) O11_N2_S2 <=     O11_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O11_N0_S3;		always @(posedge clk) O11_N0_S3 <=     O11_N0_S2  +  O11_N2_S2 ;
 assign conv_mac_11 = O11_N0_S3;

logic signed [31:0] conv_mac_12;
logic signed [63:0] chainout_0_O12; 
logic signed [63:0] O12_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O12(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_12[7:0]),.ay( 9'sd2),.bx(input_fmap_12[15:8]),.by(-9'sd3),.cx(input_fmap_12[23:16]),.cy( 9'sd4),.dx(input_fmap_12[31:24]),.dy(-9'sd4),.chainin(63'd0),.result(O12_N0_S1),.chainout(chainout_0_O12));
logic signed [63:0] chainout_2_O12; 
logic signed [63:0] O12_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O12(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_12[39:32]),.ay( 9'sd29),.bx(input_fmap_12[47:40]),.by( 9'sd1),.cx(input_fmap_12[55:48]),.cy( 9'sd1),.dx(input_fmap_12[63:56]),.dy(-9'sd4),.chainin(63'd0),.result(O12_N2_S1),.chainout(chainout_2_O12));
logic signed [63:0] chainout_4_O12; 
logic signed [63:0] O12_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O12(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_12[71:64]),.ay( 9'sd5),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O12_N4_S1),.chainout(chainout_4_O12));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O12_N0_S2;		always @(posedge clk) O12_N0_S2 <=     O12_N0_S1  +  O12_N2_S1 ;
 logic signed [21:0] O12_N2_S2;		always @(posedge clk) O12_N2_S2 <=     O12_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O12_N0_S3;		always @(posedge clk) O12_N0_S3 <=     O12_N0_S2  +  O12_N2_S2 ;
 assign conv_mac_12 = O12_N0_S3;

logic signed [31:0] conv_mac_13;
logic signed [63:0] chainout_0_O13; 
logic signed [63:0] O13_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O13(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_13[7:0]),.ay( 9'sd2),.bx(input_fmap_13[15:8]),.by(-9'sd2),.cx(input_fmap_13[23:16]),.cy( 9'sd1),.dx(input_fmap_13[31:24]),.dy( 9'sd3),.chainin(63'd0),.result(O13_N0_S1),.chainout(chainout_0_O13));
logic signed [63:0] chainout_2_O13; 
logic signed [63:0] O13_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O13(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_13[39:32]),.ay(-9'sd2),.bx(input_fmap_13[47:40]),.by(-9'sd4),.cx(input_fmap_13[55:48]),.cy(-9'sd7),.dx(input_fmap_13[63:56]),.dy(-9'sd12),.chainin(63'd0),.result(O13_N2_S1),.chainout(chainout_2_O13));
logic signed [63:0] chainout_4_O13; 
logic signed [63:0] O13_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O13(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_13[71:64]),.ay(-9'sd5),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O13_N4_S1),.chainout(chainout_4_O13));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O13_N0_S2;		always @(posedge clk) O13_N0_S2 <=     O13_N0_S1  +  O13_N2_S1 ;
 logic signed [21:0] O13_N2_S2;		always @(posedge clk) O13_N2_S2 <=     O13_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O13_N0_S3;		always @(posedge clk) O13_N0_S3 <=     O13_N0_S2  +  O13_N2_S2 ;
 assign conv_mac_13 = O13_N0_S3;

logic signed [31:0] conv_mac_14;
logic signed [63:0] chainout_0_O14; 
logic signed [63:0] O14_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O14(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_14[7:0]),.ay( 9'sd1),.bx(input_fmap_14[15:8]),.by(-9'sd5),.cx(input_fmap_14[23:16]),.cy( 9'sd5),.dx(input_fmap_14[31:24]),.dy(-9'sd5),.chainin(63'd0),.result(O14_N0_S1),.chainout(chainout_0_O14));
logic signed [63:0] chainout_2_O14; 
logic signed [63:0] O14_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O14(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_14[39:32]),.ay(-9'sd7),.bx(input_fmap_14[47:40]),.by( 9'sd23),.cx(input_fmap_14[63:56]),.cy( 9'sd5),.dx(input_fmap_14[71:64]),.dy( 9'sd6),.chainin(63'd0),.result(O14_N2_S1),.chainout(chainout_2_O14));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O14_N0_S2;		always @(posedge clk) O14_N0_S2 <=     O14_N0_S1  +  O14_N2_S1 ;
 assign conv_mac_14 = O14_N0_S2;

logic signed [31:0] conv_mac_15;
logic signed [63:0] chainout_0_O15; 
logic signed [63:0] O15_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O15(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_15[7:0]),.ay( 9'sd4),.bx(input_fmap_15[15:8]),.by(-9'sd3),.cx(input_fmap_15[23:16]),.cy( 9'sd6),.dx(input_fmap_15[31:24]),.dy( 9'sd11),.chainin(63'd0),.result(O15_N0_S1),.chainout(chainout_0_O15));
logic signed [63:0] chainout_2_O15; 
logic signed [63:0] O15_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O15(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_15[39:32]),.ay( 9'sd27),.bx(input_fmap_15[47:40]),.by(-9'sd7),.cx(input_fmap_15[55:48]),.cy(-9'sd6),.dx(input_fmap_15[63:56]),.dy(-9'sd9),.chainin(63'd0),.result(O15_N2_S1),.chainout(chainout_2_O15));
logic signed [63:0] chainout_4_O15; 
logic signed [63:0] O15_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O15(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_15[71:64]),.ay(-9'sd4),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O15_N4_S1),.chainout(chainout_4_O15));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O15_N0_S2;		always @(posedge clk) O15_N0_S2 <=     O15_N0_S1  +  O15_N2_S1 ;
 logic signed [21:0] O15_N2_S2;		always @(posedge clk) O15_N2_S2 <=     O15_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O15_N0_S3;		always @(posedge clk) O15_N0_S3 <=     O15_N0_S2  +  O15_N2_S2 ;
 assign conv_mac_15 = O15_N0_S3;

logic signed [31:0] conv_mac_16;
logic signed [63:0] chainout_0_O16; 
logic signed [63:0] O16_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O16(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_16[7:0]),.ay( 9'sd4),.bx(input_fmap_16[15:8]),.by( 9'sd17),.cx(input_fmap_16[23:16]),.cy( 9'sd4),.dx(input_fmap_16[31:24]),.dy(-9'sd5),.chainin(63'd0),.result(O16_N0_S1),.chainout(chainout_0_O16));
logic signed [63:0] chainout_2_O16; 
logic signed [63:0] O16_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O16(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_16[39:32]),.ay( 9'sd11),.bx(input_fmap_16[47:40]),.by(-9'sd6),.cx(input_fmap_16[55:48]),.cy(-9'sd3),.dx(input_fmap_16[63:56]),.dy( 9'sd5),.chainin(63'd0),.result(O16_N2_S1),.chainout(chainout_2_O16));
logic signed [63:0] chainout_4_O16; 
logic signed [63:0] O16_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O16(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_16[71:64]),.ay(-9'sd4),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O16_N4_S1),.chainout(chainout_4_O16));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O16_N0_S2;		always @(posedge clk) O16_N0_S2 <=     O16_N0_S1  +  O16_N2_S1 ;
 logic signed [21:0] O16_N2_S2;		always @(posedge clk) O16_N2_S2 <=     O16_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O16_N0_S3;		always @(posedge clk) O16_N0_S3 <=     O16_N0_S2  +  O16_N2_S2 ;
 assign conv_mac_16 = O16_N0_S3;

logic signed [31:0] conv_mac_17;
logic signed [63:0] chainout_0_O17; 
logic signed [63:0] O17_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O17(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_17[7:0]),.ay( 9'sd3),.bx(input_fmap_17[15:8]),.by(-9'sd2),.cx(input_fmap_17[23:16]),.cy(-9'sd6),.dx(input_fmap_17[31:24]),.dy(-9'sd22),.chainin(63'd0),.result(O17_N0_S1),.chainout(chainout_0_O17));
logic signed [63:0] chainout_2_O17; 
logic signed [63:0] O17_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O17(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_17[39:32]),.ay( 9'sd13),.bx(input_fmap_17[47:40]),.by( 9'sd8),.cx(input_fmap_17[55:48]),.cy(-9'sd11),.dx(input_fmap_17[63:56]),.dy( 9'sd2),.chainin(63'd0),.result(O17_N2_S1),.chainout(chainout_2_O17));
logic signed [63:0] chainout_4_O17; 
logic signed [63:0] O17_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O17(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_17[71:64]),.ay( 9'sd9),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O17_N4_S1),.chainout(chainout_4_O17));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O17_N0_S2;		always @(posedge clk) O17_N0_S2 <=     O17_N0_S1  +  O17_N2_S1 ;
 logic signed [21:0] O17_N2_S2;		always @(posedge clk) O17_N2_S2 <=     O17_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O17_N0_S3;		always @(posedge clk) O17_N0_S3 <=     O17_N0_S2  +  O17_N2_S2 ;
 assign conv_mac_17 = O17_N0_S3;

logic signed [31:0] conv_mac_18;
logic signed [63:0] chainout_0_O18; 
logic signed [63:0] O18_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O18(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_18[7:0]),.ay(-9'sd9),.bx(input_fmap_18[15:8]),.by( 9'sd4),.cx(input_fmap_18[23:16]),.cy( 9'sd1),.dx(input_fmap_18[31:24]),.dy( 9'sd4),.chainin(63'd0),.result(O18_N0_S1),.chainout(chainout_0_O18));
logic signed [63:0] chainout_2_O18; 
logic signed [63:0] O18_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O18(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_18[39:32]),.ay( 9'sd25),.bx(input_fmap_18[47:40]),.by( 9'sd8),.cx(input_fmap_18[55:48]),.cy(-9'sd9),.dx(input_fmap_18[63:56]),.dy( 9'sd1),.chainin(63'd0),.result(O18_N2_S1),.chainout(chainout_2_O18));
logic signed [63:0] chainout_4_O18; 
logic signed [63:0] O18_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O18(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_18[71:64]),.ay( 9'sd3),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O18_N4_S1),.chainout(chainout_4_O18));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O18_N0_S2;		always @(posedge clk) O18_N0_S2 <=     O18_N0_S1  +  O18_N2_S1 ;
 logic signed [21:0] O18_N2_S2;		always @(posedge clk) O18_N2_S2 <=     O18_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O18_N0_S3;		always @(posedge clk) O18_N0_S3 <=     O18_N0_S2  +  O18_N2_S2 ;
 assign conv_mac_18 = O18_N0_S3;

logic signed [31:0] conv_mac_19;
logic signed [63:0] chainout_0_O19; 
logic signed [63:0] O19_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O19(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_19[7:0]),.ay( 9'sd4),.bx(input_fmap_19[15:8]),.by(-9'sd10),.cx(input_fmap_19[23:16]),.cy( 9'sd3),.dx(input_fmap_19[31:24]),.dy(-9'sd6),.chainin(63'd0),.result(O19_N0_S1),.chainout(chainout_0_O19));
logic signed [63:0] chainout_2_O19; 
logic signed [63:0] O19_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O19(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_19[39:32]),.ay( 9'sd42),.bx(input_fmap_19[47:40]),.by(-9'sd5),.cx(input_fmap_19[55:48]),.cy( 9'sd2),.dx(input_fmap_19[63:56]),.dy(-9'sd1),.chainin(63'd0),.result(O19_N2_S1),.chainout(chainout_2_O19));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O19_N0_S2;		always @(posedge clk) O19_N0_S2 <=     O19_N0_S1  +  O19_N2_S1 ;
 assign conv_mac_19 = O19_N0_S2;

logic signed [31:0] conv_mac_20;
logic signed [63:0] chainout_0_O20; 
logic signed [63:0] O20_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O20(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_20[7:0]),.ay( 9'sd4),.bx(input_fmap_20[15:8]),.by( 9'sd8),.cx(input_fmap_20[23:16]),.cy( 9'sd1),.dx(input_fmap_20[31:24]),.dy(-9'sd2),.chainin(63'd0),.result(O20_N0_S1),.chainout(chainout_0_O20));
logic signed [63:0] chainout_2_O20; 
logic signed [63:0] O20_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O20(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_20[39:32]),.ay(-9'sd22),.bx(input_fmap_20[47:40]),.by( 9'sd3),.cx(input_fmap_20[55:48]),.cy( 9'sd1),.dx(input_fmap_20[63:56]),.dy(-9'sd8),.chainin(63'd0),.result(O20_N2_S1),.chainout(chainout_2_O20));
logic signed [63:0] chainout_4_O20; 
logic signed [63:0] O20_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O20(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_20[71:64]),.ay(-9'sd4),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O20_N4_S1),.chainout(chainout_4_O20));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O20_N0_S2;		always @(posedge clk) O20_N0_S2 <=     O20_N0_S1  +  O20_N2_S1 ;
 logic signed [21:0] O20_N2_S2;		always @(posedge clk) O20_N2_S2 <=     O20_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O20_N0_S3;		always @(posedge clk) O20_N0_S3 <=     O20_N0_S2  +  O20_N2_S2 ;
 assign conv_mac_20 = O20_N0_S3;

logic signed [31:0] conv_mac_21;
logic signed [63:0] chainout_0_O21; 
logic signed [63:0] O21_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O21(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_21[7:0]),.ay( 9'sd3),.bx(input_fmap_21[15:8]),.by(-9'sd2),.cx(input_fmap_21[23:16]),.cy( 9'sd5),.dx(input_fmap_21[31:24]),.dy(-9'sd11),.chainin(63'd0),.result(O21_N0_S1),.chainout(chainout_0_O21));
logic signed [63:0] chainout_2_O21; 
logic signed [63:0] O21_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O21(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_21[39:32]),.ay( 9'sd34),.bx(input_fmap_21[47:40]),.by(-9'sd5),.cx(input_fmap_21[55:48]),.cy(-9'sd8),.dx(input_fmap_21[63:56]),.dy( 9'sd6),.chainin(63'd0),.result(O21_N2_S1),.chainout(chainout_2_O21));
logic signed [63:0] chainout_4_O21; 
logic signed [63:0] O21_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O21(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_21[71:64]),.ay( 9'sd7),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O21_N4_S1),.chainout(chainout_4_O21));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O21_N0_S2;		always @(posedge clk) O21_N0_S2 <=     O21_N0_S1  +  O21_N2_S1 ;
 logic signed [21:0] O21_N2_S2;		always @(posedge clk) O21_N2_S2 <=     O21_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O21_N0_S3;		always @(posedge clk) O21_N0_S3 <=     O21_N0_S2  +  O21_N2_S2 ;
 assign conv_mac_21 = O21_N0_S3;

logic signed [31:0] conv_mac_22;
logic signed [63:0] chainout_0_O22; 
logic signed [63:0] O22_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O22(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_22[7:0]),.ay(-9'sd1),.bx(input_fmap_22[15:8]),.by(-9'sd3),.cx(input_fmap_22[23:16]),.cy( 9'sd5),.dx(input_fmap_22[31:24]),.dy( 9'sd4),.chainin(63'd0),.result(O22_N0_S1),.chainout(chainout_0_O22));
logic signed [63:0] chainout_2_O22; 
logic signed [63:0] O22_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O22(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_22[39:32]),.ay( 9'sd25),.bx(input_fmap_22[47:40]),.by(-9'sd2),.cx(input_fmap_22[55:48]),.cy( 9'sd6),.dx(input_fmap_22[71:64]),.dy(-9'sd3),.chainin(63'd0),.result(O22_N2_S1),.chainout(chainout_2_O22));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O22_N0_S2;		always @(posedge clk) O22_N0_S2 <=     O22_N0_S1  +  O22_N2_S1 ;
 assign conv_mac_22 = O22_N0_S2;

logic signed [31:0] conv_mac_23;
logic signed [63:0] chainout_0_O23; 
logic signed [63:0] O23_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O23(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_23[7:0]),.ay(-9'sd4),.bx(input_fmap_23[15:8]),.by(-9'sd5),.cx(input_fmap_23[23:16]),.cy(-9'sd8),.dx(input_fmap_23[31:24]),.dy( 9'sd3),.chainin(63'd0),.result(O23_N0_S1),.chainout(chainout_0_O23));
logic signed [63:0] chainout_2_O23; 
logic signed [63:0] O23_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O23(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_23[39:32]),.ay(-9'sd19),.bx(input_fmap_23[47:40]),.by(-9'sd1),.cx(input_fmap_23[55:48]),.cy( 9'sd6),.dx(input_fmap_23[63:56]),.dy( 9'sd21),.chainin(63'd0),.result(O23_N2_S1),.chainout(chainout_2_O23));
logic signed [63:0] chainout_4_O23; 
logic signed [63:0] O23_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O23(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_23[71:64]),.ay( 9'sd9),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O23_N4_S1),.chainout(chainout_4_O23));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O23_N0_S2;		always @(posedge clk) O23_N0_S2 <=     O23_N0_S1  +  O23_N2_S1 ;
 logic signed [21:0] O23_N2_S2;		always @(posedge clk) O23_N2_S2 <=     O23_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O23_N0_S3;		always @(posedge clk) O23_N0_S3 <=     O23_N0_S2  +  O23_N2_S2 ;
 assign conv_mac_23 = O23_N0_S3;

logic signed [31:0] conv_mac_24;
logic signed [63:0] chainout_0_O24; 
logic signed [63:0] O24_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O24(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_24[7:0]),.ay( 9'sd1),.bx(input_fmap_24[15:8]),.by(-9'sd1),.cx(input_fmap_24[23:16]),.cy(-9'sd6),.dx(input_fmap_24[31:24]),.dy(-9'sd1),.chainin(63'd0),.result(O24_N0_S1),.chainout(chainout_0_O24));
logic signed [63:0] chainout_2_O24; 
logic signed [63:0] O24_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O24(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_24[39:32]),.ay(-9'sd5),.bx(input_fmap_24[47:40]),.by(-9'sd5),.cx(input_fmap_24[55:48]),.cy(-9'sd6),.dx(input_fmap_24[63:56]),.dy(-9'sd4),.chainin(63'd0),.result(O24_N2_S1),.chainout(chainout_2_O24));
logic signed [63:0] chainout_4_O24; 
logic signed [63:0] O24_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O24(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_24[71:64]),.ay(-9'sd5),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O24_N4_S1),.chainout(chainout_4_O24));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O24_N0_S2;		always @(posedge clk) O24_N0_S2 <=     O24_N0_S1  +  O24_N2_S1 ;
 logic signed [21:0] O24_N2_S2;		always @(posedge clk) O24_N2_S2 <=     O24_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O24_N0_S3;		always @(posedge clk) O24_N0_S3 <=     O24_N0_S2  +  O24_N2_S2 ;
 assign conv_mac_24 = O24_N0_S3;

logic signed [31:0] conv_mac_25;
logic signed [63:0] chainout_0_O25; 
logic signed [63:0] O25_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O25(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_25[7:0]),.ay( 9'sd1),.bx(input_fmap_25[15:8]),.by(-9'sd4),.cx(input_fmap_25[23:16]),.cy( 9'sd4),.dx(input_fmap_25[31:24]),.dy(-9'sd7),.chainin(63'd0),.result(O25_N0_S1),.chainout(chainout_0_O25));
logic signed [63:0] chainout_2_O25; 
logic signed [63:0] O25_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O25(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_25[39:32]),.ay(-9'sd17),.bx(input_fmap_25[47:40]),.by(-9'sd9),.cx(input_fmap_25[55:48]),.cy( 9'sd2),.dx(input_fmap_25[63:56]),.dy(-9'sd10),.chainin(63'd0),.result(O25_N2_S1),.chainout(chainout_2_O25));
logic signed [63:0] chainout_4_O25; 
logic signed [63:0] O25_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O25(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_25[71:64]),.ay( 9'sd2),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O25_N4_S1),.chainout(chainout_4_O25));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O25_N0_S2;		always @(posedge clk) O25_N0_S2 <=     O25_N0_S1  +  O25_N2_S1 ;
 logic signed [21:0] O25_N2_S2;		always @(posedge clk) O25_N2_S2 <=     O25_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O25_N0_S3;		always @(posedge clk) O25_N0_S3 <=     O25_N0_S2  +  O25_N2_S2 ;
 assign conv_mac_25 = O25_N0_S3;

logic signed [31:0] conv_mac_26;
logic signed [63:0] chainout_0_O26; 
logic signed [63:0] O26_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O26(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_26[7:0]),.ay(-9'sd2),.bx(input_fmap_26[15:8]),.by(-9'sd6),.cx(input_fmap_26[23:16]),.cy(-9'sd2),.dx(input_fmap_26[39:32]),.dy(-9'sd10),.chainin(63'd0),.result(O26_N0_S1),.chainout(chainout_0_O26));
logic signed [63:0] chainout_2_O26; 
logic signed [63:0] O26_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O26(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_26[47:40]),.ay(-9'sd1),.bx(input_fmap_26[55:48]),.by(-9'sd3),.cx(input_fmap_26[63:56]),.cy(-9'sd6),.dx(input_fmap_26[71:64]),.dy(-9'sd6),.chainin(63'd0),.result(O26_N2_S1),.chainout(chainout_2_O26));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O26_N0_S2;		always @(posedge clk) O26_N0_S2 <=     O26_N0_S1  +  O26_N2_S1 ;
 assign conv_mac_26 = O26_N0_S2;

logic signed [31:0] conv_mac_27;
logic signed [63:0] chainout_0_O27; 
logic signed [63:0] O27_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O27(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_27[7:0]),.ay(-9'sd4),.bx(input_fmap_27[15:8]),.by(-9'sd8),.cx(input_fmap_27[23:16]),.cy(-9'sd4),.dx(input_fmap_27[31:24]),.dy(-9'sd10),.chainin(63'd0),.result(O27_N0_S1),.chainout(chainout_0_O27));
logic signed [63:0] chainout_2_O27; 
logic signed [63:0] O27_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O27(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_27[39:32]),.ay( 9'sd12),.bx(input_fmap_27[47:40]),.by( 9'sd16),.cx(input_fmap_27[55:48]),.cy(-9'sd8),.dx(input_fmap_27[63:56]),.dy( 9'sd6),.chainin(63'd0),.result(O27_N2_S1),.chainout(chainout_2_O27));
logic signed [63:0] chainout_4_O27; 
logic signed [63:0] O27_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O27(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_27[71:64]),.ay( 9'sd3),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O27_N4_S1),.chainout(chainout_4_O27));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O27_N0_S2;		always @(posedge clk) O27_N0_S2 <=     O27_N0_S1  +  O27_N2_S1 ;
 logic signed [21:0] O27_N2_S2;		always @(posedge clk) O27_N2_S2 <=     O27_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O27_N0_S3;		always @(posedge clk) O27_N0_S3 <=     O27_N0_S2  +  O27_N2_S2 ;
 assign conv_mac_27 = O27_N0_S3;

logic signed [31:0] conv_mac_28;
logic signed [63:0] chainout_0_O28; 
logic signed [63:0] O28_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O28(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_28[7:0]),.ay( 9'sd4),.bx(input_fmap_28[15:8]),.by( 9'sd9),.cx(input_fmap_28[23:16]),.cy( 9'sd2),.dx(input_fmap_28[31:24]),.dy(-9'sd1),.chainin(63'd0),.result(O28_N0_S1),.chainout(chainout_0_O28));
logic signed [63:0] chainout_2_O28; 
logic signed [63:0] O28_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O28(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_28[39:32]),.ay( 9'sd14),.bx(input_fmap_28[47:40]),.by( 9'sd3),.cx(input_fmap_28[55:48]),.cy(-9'sd8),.dx(input_fmap_28[63:56]),.dy( 9'sd1),.chainin(63'd0),.result(O28_N2_S1),.chainout(chainout_2_O28));
logic signed [63:0] chainout_4_O28; 
logic signed [63:0] O28_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O28(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_28[71:64]),.ay(-9'sd7),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O28_N4_S1),.chainout(chainout_4_O28));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O28_N0_S2;		always @(posedge clk) O28_N0_S2 <=     O28_N0_S1  +  O28_N2_S1 ;
 logic signed [21:0] O28_N2_S2;		always @(posedge clk) O28_N2_S2 <=     O28_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O28_N0_S3;		always @(posedge clk) O28_N0_S3 <=     O28_N0_S2  +  O28_N2_S2 ;
 assign conv_mac_28 = O28_N0_S3;

logic signed [31:0] conv_mac_29;
logic signed [63:0] chainout_0_O29; 
logic signed [63:0] O29_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O29(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_29[7:0]),.ay( 9'sd5),.bx(input_fmap_29[15:8]),.by( 9'sd10),.cx(input_fmap_29[23:16]),.cy( 9'sd11),.dx(input_fmap_29[31:24]),.dy( 9'sd13),.chainin(63'd0),.result(O29_N0_S1),.chainout(chainout_0_O29));
logic signed [63:0] chainout_2_O29; 
logic signed [63:0] O29_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O29(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_29[39:32]),.ay(-9'sd15),.bx(input_fmap_29[47:40]),.by(-9'sd3),.cx(input_fmap_29[55:48]),.cy( 9'sd10),.dx(input_fmap_29[63:56]),.dy(-9'sd10),.chainin(63'd0),.result(O29_N2_S1),.chainout(chainout_2_O29));
logic signed [63:0] chainout_4_O29; 
logic signed [63:0] O29_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O29(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_29[71:64]),.ay(-9'sd4),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O29_N4_S1),.chainout(chainout_4_O29));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O29_N0_S2;		always @(posedge clk) O29_N0_S2 <=     O29_N0_S1  +  O29_N2_S1 ;
 logic signed [21:0] O29_N2_S2;		always @(posedge clk) O29_N2_S2 <=     O29_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O29_N0_S3;		always @(posedge clk) O29_N0_S3 <=     O29_N0_S2  +  O29_N2_S2 ;
 assign conv_mac_29 = O29_N0_S3;

logic signed [31:0] conv_mac_30;
logic signed [63:0] chainout_0_O30; 
logic signed [63:0] O30_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O30(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_30[7:0]),.ay( 9'sd3),.bx(input_fmap_30[15:8]),.by(-9'sd3),.cx(input_fmap_30[39:32]),.cy( 9'sd23),.dx(input_fmap_30[47:40]),.dy(-9'sd3),.chainin(63'd0),.result(O30_N0_S1),.chainout(chainout_0_O30));
logic signed [63:0] chainout_2_O30; 
logic signed [63:0] O30_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O30(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_30[55:48]),.ay( 9'sd2),.bx(input_fmap_30[63:56]),.by( 9'sd1),.cx(input_fmap_30[71:64]),.cy( 9'sd3),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O30_N2_S1),.chainout(chainout_2_O30));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O30_N0_S2;		always @(posedge clk) O30_N0_S2 <=     O30_N0_S1  +  O30_N2_S1 ;
 assign conv_mac_30 = O30_N0_S2;

logic signed [31:0] conv_mac_31;
logic signed [63:0] chainout_0_O31; 
logic signed [63:0] O31_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O31(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_31[7:0]),.ay(-9'sd6),.bx(input_fmap_31[15:8]),.by(-9'sd11),.cx(input_fmap_31[23:16]),.cy( 9'sd3),.dx(input_fmap_31[39:32]),.dy( 9'sd14),.chainin(63'd0),.result(O31_N0_S1),.chainout(chainout_0_O31));
logic signed [63:0] chainout_2_O31; 
logic signed [63:0] O31_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O31(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_31[47:40]),.ay( 9'sd12),.bx(input_fmap_31[55:48]),.by( 9'sd7),.cx(input_fmap_31[63:56]),.cy( 9'sd11),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O31_N2_S1),.chainout(chainout_2_O31));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O31_N0_S2;		always @(posedge clk) O31_N0_S2 <=     O31_N0_S1  +  O31_N2_S1 ;
 assign conv_mac_31 = O31_N0_S2;

logic signed [31:0] conv_mac_32;
logic signed [63:0] chainout_0_O32; 
logic signed [63:0] O32_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O32(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_32[7:0]),.ay(-9'sd5),.bx(input_fmap_32[15:8]),.by( 9'sd1),.cx(input_fmap_32[23:16]),.cy(-9'sd3),.dx(input_fmap_32[31:24]),.dy(-9'sd5),.chainin(63'd0),.result(O32_N0_S1),.chainout(chainout_0_O32));
logic signed [63:0] chainout_2_O32; 
logic signed [63:0] O32_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O32(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_32[39:32]),.ay(-9'sd21),.bx(input_fmap_32[47:40]),.by( 9'sd1),.cx(input_fmap_32[55:48]),.cy( 9'sd9),.dx(input_fmap_32[63:56]),.dy( 9'sd31),.chainin(63'd0),.result(O32_N2_S1),.chainout(chainout_2_O32));
logic signed [63:0] chainout_4_O32; 
logic signed [63:0] O32_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O32(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_32[71:64]),.ay(-9'sd12),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O32_N4_S1),.chainout(chainout_4_O32));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O32_N0_S2;		always @(posedge clk) O32_N0_S2 <=     O32_N0_S1  +  O32_N2_S1 ;
 logic signed [21:0] O32_N2_S2;		always @(posedge clk) O32_N2_S2 <=     O32_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O32_N0_S3;		always @(posedge clk) O32_N0_S3 <=     O32_N0_S2  +  O32_N2_S2 ;
 assign conv_mac_32 = O32_N0_S3;

logic signed [31:0] conv_mac_33;
logic signed [63:0] chainout_0_O33; 
logic signed [63:0] O33_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O33(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_33[7:0]),.ay( 9'sd1),.bx(input_fmap_33[15:8]),.by(-9'sd6),.cx(input_fmap_33[23:16]),.cy(-9'sd3),.dx(input_fmap_33[31:24]),.dy(-9'sd7),.chainin(63'd0),.result(O33_N0_S1),.chainout(chainout_0_O33));
logic signed [63:0] chainout_2_O33; 
logic signed [63:0] O33_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O33(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_33[39:32]),.ay(-9'sd16),.bx(input_fmap_33[55:48]),.by(-9'sd1),.cx(input_fmap_33[63:56]),.cy( 9'sd3),.dx(input_fmap_33[71:64]),.dy( 9'sd3),.chainin(63'd0),.result(O33_N2_S1),.chainout(chainout_2_O33));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O33_N0_S2;		always @(posedge clk) O33_N0_S2 <=     O33_N0_S1  +  O33_N2_S1 ;
 assign conv_mac_33 = O33_N0_S2;

logic signed [31:0] conv_mac_34;
logic signed [63:0] chainout_0_O34; 
logic signed [63:0] O34_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O34(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_34[7:0]),.ay( 9'sd2),.bx(input_fmap_34[15:8]),.by(-9'sd9),.cx(input_fmap_34[23:16]),.cy(-9'sd8),.dx(input_fmap_34[39:32]),.dy( 9'sd22),.chainin(63'd0),.result(O34_N0_S1),.chainout(chainout_0_O34));
logic signed [63:0] chainout_2_O34; 
logic signed [63:0] O34_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O34(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_34[47:40]),.ay(-9'sd2),.bx(input_fmap_34[55:48]),.by(-9'sd2),.cx(input_fmap_34[63:56]),.cy( 9'sd11),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O34_N2_S1),.chainout(chainout_2_O34));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O34_N0_S2;		always @(posedge clk) O34_N0_S2 <=     O34_N0_S1  +  O34_N2_S1 ;
 assign conv_mac_34 = O34_N0_S2;

logic signed [31:0] conv_mac_35;
logic signed [63:0] chainout_0_O35; 
logic signed [63:0] O35_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O35(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_35[7:0]),.ay( 9'sd2),.bx(input_fmap_35[15:8]),.by(-9'sd4),.cx(input_fmap_35[23:16]),.cy( 9'sd2),.dx(input_fmap_35[31:24]),.dy( 9'sd1),.chainin(63'd0),.result(O35_N0_S1),.chainout(chainout_0_O35));
logic signed [63:0] chainout_2_O35; 
logic signed [63:0] O35_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O35(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_35[39:32]),.ay( 9'sd22),.bx(input_fmap_35[47:40]),.by( 9'sd7),.cx(input_fmap_35[63:56]),.cy( 9'sd4),.dx(input_fmap_35[71:64]),.dy( 9'sd3),.chainin(63'd0),.result(O35_N2_S1),.chainout(chainout_2_O35));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O35_N0_S2;		always @(posedge clk) O35_N0_S2 <=     O35_N0_S1  +  O35_N2_S1 ;
 assign conv_mac_35 = O35_N0_S2;

logic signed [31:0] conv_mac_36;
logic signed [63:0] chainout_0_O36; 
logic signed [63:0] O36_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O36(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_36[7:0]),.ay(-9'sd6),.bx(input_fmap_36[15:8]),.by(-9'sd9),.cx(input_fmap_36[23:16]),.cy(-9'sd2),.dx(input_fmap_36[31:24]),.dy(-9'sd2),.chainin(63'd0),.result(O36_N0_S1),.chainout(chainout_0_O36));
logic signed [63:0] chainout_2_O36; 
logic signed [63:0] O36_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O36(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_36[39:32]),.ay( 9'sd8),.bx(input_fmap_36[63:56]),.by( 9'sd26),.cx(input_fmap_36[71:64]),.cy(-9'sd2),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O36_N2_S1),.chainout(chainout_2_O36));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O36_N0_S2;		always @(posedge clk) O36_N0_S2 <=     O36_N0_S1  +  O36_N2_S1 ;
 assign conv_mac_36 = O36_N0_S2;

logic signed [31:0] conv_mac_37;
logic signed [63:0] chainout_0_O37; 
logic signed [63:0] O37_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O37(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_37[7:0]),.ay(-9'sd2),.bx(input_fmap_37[15:8]),.by(-9'sd7),.cx(input_fmap_37[23:16]),.cy( 9'sd4),.dx(input_fmap_37[39:32]),.dy(-9'sd3),.chainin(63'd0),.result(O37_N0_S1),.chainout(chainout_0_O37));
logic signed [63:0] chainout_2_O37; 
logic signed [63:0] O37_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O37(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_37[47:40]),.ay(-9'sd11),.bx(input_fmap_37[63:56]),.by(-9'sd6),.cx(input_fmap_37[71:64]),.cy(-9'sd6),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O37_N2_S1),.chainout(chainout_2_O37));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O37_N0_S2;		always @(posedge clk) O37_N0_S2 <=     O37_N0_S1  +  O37_N2_S1 ;
 assign conv_mac_37 = O37_N0_S2;

logic signed [31:0] conv_mac_38;
logic signed [63:0] chainout_0_O38; 
logic signed [63:0] O38_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O38(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_38[7:0]),.ay(-9'sd4),.bx(input_fmap_38[15:8]),.by(-9'sd12),.cx(input_fmap_38[23:16]),.cy( 9'sd1),.dx(input_fmap_38[31:24]),.dy(-9'sd16),.chainin(63'd0),.result(O38_N0_S1),.chainout(chainout_0_O38));
logic signed [63:0] chainout_2_O38; 
logic signed [63:0] O38_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O38(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_38[39:32]),.ay( 9'sd24),.bx(input_fmap_38[47:40]),.by( 9'sd13),.cx(input_fmap_38[55:48]),.cy(-9'sd4),.dx(input_fmap_38[63:56]),.dy( 9'sd6),.chainin(63'd0),.result(O38_N2_S1),.chainout(chainout_2_O38));
logic signed [63:0] chainout_4_O38; 
logic signed [63:0] O38_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O38(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_38[71:64]),.ay( 9'sd4),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O38_N4_S1),.chainout(chainout_4_O38));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O38_N0_S2;		always @(posedge clk) O38_N0_S2 <=     O38_N0_S1  +  O38_N2_S1 ;
 logic signed [21:0] O38_N2_S2;		always @(posedge clk) O38_N2_S2 <=     O38_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O38_N0_S3;		always @(posedge clk) O38_N0_S3 <=     O38_N0_S2  +  O38_N2_S2 ;
 assign conv_mac_38 = O38_N0_S3;

logic signed [31:0] conv_mac_39;
logic signed [63:0] chainout_0_O39; 
logic signed [63:0] O39_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O39(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_39[7:0]),.ay( 9'sd7),.bx(input_fmap_39[15:8]),.by(-9'sd10),.cx(input_fmap_39[23:16]),.cy(-9'sd5),.dx(input_fmap_39[31:24]),.dy( 9'sd2),.chainin(63'd0),.result(O39_N0_S1),.chainout(chainout_0_O39));
logic signed [63:0] chainout_2_O39; 
logic signed [63:0] O39_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O39(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_39[39:32]),.ay( 9'sd22),.bx(input_fmap_39[47:40]),.by(-9'sd9),.cx(input_fmap_39[55:48]),.cy(-9'sd4),.dx(input_fmap_39[63:56]),.dy( 9'sd4),.chainin(63'd0),.result(O39_N2_S1),.chainout(chainout_2_O39));
logic signed [63:0] chainout_4_O39; 
logic signed [63:0] O39_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O39(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_39[71:64]),.ay( 9'sd2),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O39_N4_S1),.chainout(chainout_4_O39));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O39_N0_S2;		always @(posedge clk) O39_N0_S2 <=     O39_N0_S1  +  O39_N2_S1 ;
 logic signed [21:0] O39_N2_S2;		always @(posedge clk) O39_N2_S2 <=     O39_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O39_N0_S3;		always @(posedge clk) O39_N0_S3 <=     O39_N0_S2  +  O39_N2_S2 ;
 assign conv_mac_39 = O39_N0_S3;

logic signed [31:0] conv_mac_40;
logic signed [63:0] chainout_0_O40; 
logic signed [63:0] O40_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O40(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_40[7:0]),.ay(-9'sd6),.bx(input_fmap_40[15:8]),.by( 9'sd12),.cx(input_fmap_40[23:16]),.cy( 9'sd1),.dx(input_fmap_40[31:24]),.dy(-9'sd7),.chainin(63'd0),.result(O40_N0_S1),.chainout(chainout_0_O40));
logic signed [63:0] chainout_2_O40; 
logic signed [63:0] O40_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O40(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_40[39:32]),.ay( 9'sd19),.bx(input_fmap_40[47:40]),.by( 9'sd6),.cx(input_fmap_40[55:48]),.cy(-9'sd2),.dx(input_fmap_40[63:56]),.dy(-9'sd8),.chainin(63'd0),.result(O40_N2_S1),.chainout(chainout_2_O40));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O40_N0_S2;		always @(posedge clk) O40_N0_S2 <=     O40_N0_S1  +  O40_N2_S1 ;
 assign conv_mac_40 = O40_N0_S2;

logic signed [31:0] conv_mac_41;
logic signed [63:0] chainout_0_O41; 
logic signed [63:0] O41_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O41(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_41[7:0]),.ay(-9'sd1),.bx(input_fmap_41[15:8]),.by(-9'sd5),.cx(input_fmap_41[23:16]),.cy( 9'sd1),.dx(input_fmap_41[31:24]),.dy(-9'sd1),.chainin(63'd0),.result(O41_N0_S1),.chainout(chainout_0_O41));
logic signed [63:0] chainout_2_O41; 
logic signed [63:0] O41_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O41(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_41[39:32]),.ay( 9'sd18),.bx(input_fmap_41[47:40]),.by( 9'sd3),.cx(input_fmap_41[55:48]),.cy( 9'sd1),.dx(input_fmap_41[63:56]),.dy( 9'sd4),.chainin(63'd0),.result(O41_N2_S1),.chainout(chainout_2_O41));
logic signed [63:0] chainout_4_O41; 
logic signed [63:0] O41_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O41(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_41[71:64]),.ay( 9'sd6),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O41_N4_S1),.chainout(chainout_4_O41));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O41_N0_S2;		always @(posedge clk) O41_N0_S2 <=     O41_N0_S1  +  O41_N2_S1 ;
 logic signed [21:0] O41_N2_S2;		always @(posedge clk) O41_N2_S2 <=     O41_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O41_N0_S3;		always @(posedge clk) O41_N0_S3 <=     O41_N0_S2  +  O41_N2_S2 ;
 assign conv_mac_41 = O41_N0_S3;

logic signed [31:0] conv_mac_42;
logic signed [63:0] chainout_0_O42; 
logic signed [63:0] O42_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O42(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_42[7:0]),.ay( 9'sd7),.bx(input_fmap_42[15:8]),.by(-9'sd5),.cx(input_fmap_42[23:16]),.cy(-9'sd1),.dx(input_fmap_42[31:24]),.dy( 9'sd15),.chainin(63'd0),.result(O42_N0_S1),.chainout(chainout_0_O42));
logic signed [63:0] chainout_2_O42; 
logic signed [63:0] O42_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O42(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_42[39:32]),.ay( 9'sd10),.bx(input_fmap_42[47:40]),.by(-9'sd11),.cx(input_fmap_42[55:48]),.cy( 9'sd1),.dx(input_fmap_42[63:56]),.dy( 9'sd14),.chainin(63'd0),.result(O42_N2_S1),.chainout(chainout_2_O42));
logic signed [63:0] chainout_4_O42; 
logic signed [63:0] O42_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O42(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_42[71:64]),.ay(-9'sd4),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O42_N4_S1),.chainout(chainout_4_O42));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O42_N0_S2;		always @(posedge clk) O42_N0_S2 <=     O42_N0_S1  +  O42_N2_S1 ;
 logic signed [21:0] O42_N2_S2;		always @(posedge clk) O42_N2_S2 <=     O42_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O42_N0_S3;		always @(posedge clk) O42_N0_S3 <=     O42_N0_S2  +  O42_N2_S2 ;
 assign conv_mac_42 = O42_N0_S3;

logic signed [31:0] conv_mac_43;
logic signed [63:0] chainout_0_O43; 
logic signed [63:0] O43_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O43(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_43[7:0]),.ay( 9'sd4),.bx(input_fmap_43[15:8]),.by(-9'sd9),.cx(input_fmap_43[31:24]),.cy(-9'sd6),.dx(input_fmap_43[39:32]),.dy( 9'sd27),.chainin(63'd0),.result(O43_N0_S1),.chainout(chainout_0_O43));
logic signed [63:0] chainout_2_O43; 
logic signed [63:0] O43_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O43(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_43[47:40]),.ay(-9'sd5),.bx(input_fmap_43[55:48]),.by( 9'sd2),.cx(input_fmap_43[63:56]),.cy(-9'sd6),.dx(input_fmap_43[71:64]),.dy( 9'sd7),.chainin(63'd0),.result(O43_N2_S1),.chainout(chainout_2_O43));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O43_N0_S2;		always @(posedge clk) O43_N0_S2 <=     O43_N0_S1  +  O43_N2_S1 ;
 assign conv_mac_43 = O43_N0_S2;

logic signed [31:0] conv_mac_44;
logic signed [63:0] chainout_0_O44; 
logic signed [63:0] O44_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O44(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_44[7:0]),.ay( 9'sd3),.bx(input_fmap_44[15:8]),.by( 9'sd10),.cx(input_fmap_44[23:16]),.cy(-9'sd6),.dx(input_fmap_44[39:32]),.dy( 9'sd11),.chainin(63'd0),.result(O44_N0_S1),.chainout(chainout_0_O44));
logic signed [63:0] chainout_2_O44; 
logic signed [63:0] O44_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O44(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_44[47:40]),.ay( 9'sd7),.bx(input_fmap_44[55:48]),.by(-9'sd1),.cx(input_fmap_44[63:56]),.cy( 9'sd2),.dx(input_fmap_44[71:64]),.dy( 9'sd5),.chainin(63'd0),.result(O44_N2_S1),.chainout(chainout_2_O44));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O44_N0_S2;		always @(posedge clk) O44_N0_S2 <=     O44_N0_S1  +  O44_N2_S1 ;
 assign conv_mac_44 = O44_N0_S2;

logic signed [31:0] conv_mac_45;
logic signed [63:0] chainout_0_O45; 
logic signed [63:0] O45_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O45(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_45[15:8]),.ay(-9'sd9),.bx(input_fmap_45[31:24]),.by( 9'sd3),.cx(input_fmap_45[39:32]),.cy(-9'sd13),.dx(input_fmap_45[47:40]),.dy( 9'sd4),.chainin(63'd0),.result(O45_N0_S1),.chainout(chainout_0_O45));
logic signed [63:0] chainout_2_O45; 
logic signed [63:0] O45_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O45(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_45[55:48]),.ay(-9'sd5),.bx(input_fmap_45[63:56]),.by(-9'sd7),.cx(input_fmap_45[71:64]),.cy(-9'sd3),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O45_N2_S1),.chainout(chainout_2_O45));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O45_N0_S2;		always @(posedge clk) O45_N0_S2 <=     O45_N0_S1  +  O45_N2_S1 ;
 assign conv_mac_45 = O45_N0_S2;

logic signed [31:0] conv_mac_46;
logic signed [63:0] chainout_0_O46; 
logic signed [63:0] O46_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O46(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_46[7:0]),.ay(-9'sd7),.bx(input_fmap_46[15:8]),.by( 9'sd13),.cx(input_fmap_46[23:16]),.cy( 9'sd4),.dx(input_fmap_46[31:24]),.dy(-9'sd4),.chainin(63'd0),.result(O46_N0_S1),.chainout(chainout_0_O46));
logic signed [63:0] chainout_2_O46; 
logic signed [63:0] O46_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O46(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_46[39:32]),.ay( 9'sd23),.bx(input_fmap_46[47:40]),.by( 9'sd4),.cx(input_fmap_46[55:48]),.cy(-9'sd2),.dx(input_fmap_46[63:56]),.dy(-9'sd17),.chainin(63'd0),.result(O46_N2_S1),.chainout(chainout_2_O46));
logic signed [63:0] chainout_4_O46; 
logic signed [63:0] O46_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O46(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_46[71:64]),.ay(-9'sd2),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O46_N4_S1),.chainout(chainout_4_O46));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O46_N0_S2;		always @(posedge clk) O46_N0_S2 <=     O46_N0_S1  +  O46_N2_S1 ;
 logic signed [21:0] O46_N2_S2;		always @(posedge clk) O46_N2_S2 <=     O46_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O46_N0_S3;		always @(posedge clk) O46_N0_S3 <=     O46_N0_S2  +  O46_N2_S2 ;
 assign conv_mac_46 = O46_N0_S3;

logic signed [31:0] conv_mac_47;
logic signed [63:0] chainout_0_O47; 
logic signed [63:0] O47_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O47(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_47[7:0]),.ay(-9'sd3),.bx(input_fmap_47[15:8]),.by(-9'sd6),.cx(input_fmap_47[31:24]),.cy(-9'sd8),.dx(input_fmap_47[39:32]),.dy( 9'sd29),.chainin(63'd0),.result(O47_N0_S1),.chainout(chainout_0_O47));
logic signed [63:0] chainout_2_O47; 
logic signed [63:0] O47_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O47(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_47[47:40]),.ay( 9'sd11),.bx(input_fmap_47[55:48]),.by(-9'sd4),.cx(input_fmap_47[63:56]),.cy(-9'sd2),.dx(input_fmap_47[71:64]),.dy( 9'sd3),.chainin(63'd0),.result(O47_N2_S1),.chainout(chainout_2_O47));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O47_N0_S2;		always @(posedge clk) O47_N0_S2 <=     O47_N0_S1  +  O47_N2_S1 ;
 assign conv_mac_47 = O47_N0_S2;

logic signed [31:0] conv_mac_48;
logic signed [63:0] chainout_0_O48; 
logic signed [63:0] O48_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O48(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_48[7:0]),.ay( 9'sd2),.bx(input_fmap_48[15:8]),.by( 9'sd1),.cx(input_fmap_48[23:16]),.cy( 9'sd4),.dx(input_fmap_48[31:24]),.dy(-9'sd14),.chainin(63'd0),.result(O48_N0_S1),.chainout(chainout_0_O48));
logic signed [63:0] chainout_2_O48; 
logic signed [63:0] O48_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O48(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_48[39:32]),.ay(-9'sd11),.bx(input_fmap_48[47:40]),.by( 9'sd18),.cx(input_fmap_48[55:48]),.cy(-9'sd4),.dx(input_fmap_48[63:56]),.dy(-9'sd1),.chainin(63'd0),.result(O48_N2_S1),.chainout(chainout_2_O48));
logic signed [63:0] chainout_4_O48; 
logic signed [63:0] O48_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O48(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_48[71:64]),.ay( 9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O48_N4_S1),.chainout(chainout_4_O48));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O48_N0_S2;		always @(posedge clk) O48_N0_S2 <=     O48_N0_S1  +  O48_N2_S1 ;
 logic signed [21:0] O48_N2_S2;		always @(posedge clk) O48_N2_S2 <=     O48_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O48_N0_S3;		always @(posedge clk) O48_N0_S3 <=     O48_N0_S2  +  O48_N2_S2 ;
 assign conv_mac_48 = O48_N0_S3;

logic signed [31:0] conv_mac_49;
logic signed [63:0] chainout_0_O49; 
logic signed [63:0] O49_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O49(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_49[7:0]),.ay( 9'sd3),.bx(input_fmap_49[15:8]),.by( 9'sd12),.cx(input_fmap_49[23:16]),.cy( 9'sd4),.dx(input_fmap_49[31:24]),.dy(-9'sd7),.chainin(63'd0),.result(O49_N0_S1),.chainout(chainout_0_O49));
logic signed [63:0] chainout_2_O49; 
logic signed [63:0] O49_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O49(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_49[39:32]),.ay( 9'sd7),.bx(input_fmap_49[47:40]),.by( 9'sd7),.cx(input_fmap_49[55:48]),.cy(-9'sd9),.dx(input_fmap_49[63:56]),.dy(-9'sd18),.chainin(63'd0),.result(O49_N2_S1),.chainout(chainout_2_O49));
logic signed [63:0] chainout_4_O49; 
logic signed [63:0] O49_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O49(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_49[71:64]),.ay(-9'sd10),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O49_N4_S1),.chainout(chainout_4_O49));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O49_N0_S2;		always @(posedge clk) O49_N0_S2 <=     O49_N0_S1  +  O49_N2_S1 ;
 logic signed [21:0] O49_N2_S2;		always @(posedge clk) O49_N2_S2 <=     O49_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O49_N0_S3;		always @(posedge clk) O49_N0_S3 <=     O49_N0_S2  +  O49_N2_S2 ;
 assign conv_mac_49 = O49_N0_S3;

logic signed [31:0] conv_mac_50;
logic signed [63:0] chainout_0_O50; 
logic signed [63:0] O50_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O50(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_50[15:8]),.ay(-9'sd6),.bx(input_fmap_50[23:16]),.by(-9'sd2),.cx(input_fmap_50[31:24]),.cy( 9'sd2),.dx(input_fmap_50[39:32]),.dy(-9'sd11),.chainin(63'd0),.result(O50_N0_S1),.chainout(chainout_0_O50));
logic signed [63:0] chainout_2_O50; 
logic signed [63:0] O50_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O50(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_50[55:48]),.ay(-9'sd9),.bx(input_fmap_50[63:56]),.by(-9'sd6),.cx(input_fmap_50[71:64]),.cy(-9'sd5),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O50_N2_S1),.chainout(chainout_2_O50));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O50_N0_S2;		always @(posedge clk) O50_N0_S2 <=     O50_N0_S1  +  O50_N2_S1 ;
 assign conv_mac_50 = O50_N0_S2;

logic signed [31:0] conv_mac_51;
logic signed [63:0] chainout_0_O51; 
logic signed [63:0] O51_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O51(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_51[7:0]),.ay( 9'sd2),.bx(input_fmap_51[15:8]),.by( 9'sd17),.cx(input_fmap_51[23:16]),.cy(-9'sd1),.dx(input_fmap_51[31:24]),.dy( 9'sd13),.chainin(63'd0),.result(O51_N0_S1),.chainout(chainout_0_O51));
logic signed [63:0] chainout_2_O51; 
logic signed [63:0] O51_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O51(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_51[39:32]),.ay( 9'sd13),.bx(input_fmap_51[47:40]),.by(-9'sd1),.cx(input_fmap_51[55:48]),.cy(-9'sd1),.dx(input_fmap_51[63:56]),.dy(-9'sd7),.chainin(63'd0),.result(O51_N2_S1),.chainout(chainout_2_O51));
logic signed [63:0] chainout_4_O51; 
logic signed [63:0] O51_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O51(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_51[71:64]),.ay( 9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O51_N4_S1),.chainout(chainout_4_O51));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O51_N0_S2;		always @(posedge clk) O51_N0_S2 <=     O51_N0_S1  +  O51_N2_S1 ;
 logic signed [21:0] O51_N2_S2;		always @(posedge clk) O51_N2_S2 <=     O51_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O51_N0_S3;		always @(posedge clk) O51_N0_S3 <=     O51_N0_S2  +  O51_N2_S2 ;
 assign conv_mac_51 = O51_N0_S3;

logic signed [31:0] conv_mac_52;
logic signed [63:0] chainout_0_O52; 
logic signed [63:0] O52_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O52(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_52[7:0]),.ay( 9'sd1),.bx(input_fmap_52[15:8]),.by( 9'sd21),.cx(input_fmap_52[23:16]),.cy( 9'sd2),.dx(input_fmap_52[31:24]),.dy( 9'sd1),.chainin(63'd0),.result(O52_N0_S1),.chainout(chainout_0_O52));
logic signed [63:0] chainout_2_O52; 
logic signed [63:0] O52_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O52(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_52[39:32]),.ay(-9'sd2),.bx(input_fmap_52[47:40]),.by( 9'sd4),.cx(input_fmap_52[55:48]),.cy(-9'sd2),.dx(input_fmap_52[63:56]),.dy(-9'sd8),.chainin(63'd0),.result(O52_N2_S1),.chainout(chainout_2_O52));
logic signed [63:0] chainout_4_O52; 
logic signed [63:0] O52_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O52(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_52[71:64]),.ay(-9'sd3),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O52_N4_S1),.chainout(chainout_4_O52));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O52_N0_S2;		always @(posedge clk) O52_N0_S2 <=     O52_N0_S1  +  O52_N2_S1 ;
 logic signed [21:0] O52_N2_S2;		always @(posedge clk) O52_N2_S2 <=     O52_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O52_N0_S3;		always @(posedge clk) O52_N0_S3 <=     O52_N0_S2  +  O52_N2_S2 ;
 assign conv_mac_52 = O52_N0_S3;

logic signed [31:0] conv_mac_53;
logic signed [63:0] chainout_0_O53; 
logic signed [63:0] O53_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O53(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_53[7:0]),.ay( 9'sd9),.bx(input_fmap_53[15:8]),.by( 9'sd6),.cx(input_fmap_53[23:16]),.cy(-9'sd9),.dx(input_fmap_53[31:24]),.dy( 9'sd6),.chainin(63'd0),.result(O53_N0_S1),.chainout(chainout_0_O53));
logic signed [63:0] chainout_2_O53; 
logic signed [63:0] O53_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O53(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_53[39:32]),.ay(-9'sd10),.bx(input_fmap_53[47:40]),.by(-9'sd12),.cx(input_fmap_53[55:48]),.cy(-9'sd1),.dx(input_fmap_53[71:64]),.dy(-9'sd4),.chainin(63'd0),.result(O53_N2_S1),.chainout(chainout_2_O53));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O53_N0_S2;		always @(posedge clk) O53_N0_S2 <=     O53_N0_S1  +  O53_N2_S1 ;
 assign conv_mac_53 = O53_N0_S2;

logic signed [31:0] conv_mac_54;
logic signed [63:0] chainout_0_O54; 
logic signed [63:0] O54_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O54(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_54[23:16]),.ay( 9'sd3),.bx(input_fmap_54[31:24]),.by(-9'sd2),.cx(input_fmap_54[39:32]),.cy( 9'sd25),.dx(input_fmap_54[47:40]),.dy(-9'sd3),.chainin(63'd0),.result(O54_N0_S1),.chainout(chainout_0_O54));
logic signed [63:0] chainout_2_O54; 
logic signed [63:0] O54_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O54(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_54[63:56]),.ay(-9'sd3),.bx(input_fmap_54[71:64]),.by(-9'sd2),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O54_N2_S1),.chainout(chainout_2_O54));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O54_N0_S2;		always @(posedge clk) O54_N0_S2 <=     O54_N0_S1  +  O54_N2_S1 ;
 assign conv_mac_54 = O54_N0_S2;

logic signed [31:0] conv_mac_55;
logic signed [63:0] chainout_0_O55; 
logic signed [63:0] O55_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O55(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_55[7:0]),.ay( 9'sd2),.bx(input_fmap_55[15:8]),.by( 9'sd1),.cx(input_fmap_55[23:16]),.cy( 9'sd3),.dx(input_fmap_55[31:24]),.dy(-9'sd10),.chainin(63'd0),.result(O55_N0_S1),.chainout(chainout_0_O55));
logic signed [63:0] chainout_2_O55; 
logic signed [63:0] O55_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O55(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_55[39:32]),.ay( 9'sd23),.bx(input_fmap_55[47:40]),.by( 9'sd6),.cx(input_fmap_55[55:48]),.cy( 9'sd1),.dx(input_fmap_55[63:56]),.dy(-9'sd19),.chainin(63'd0),.result(O55_N2_S1),.chainout(chainout_2_O55));
logic signed [63:0] chainout_4_O55; 
logic signed [63:0] O55_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O55(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_55[71:64]),.ay(-9'sd6),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O55_N4_S1),.chainout(chainout_4_O55));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O55_N0_S2;		always @(posedge clk) O55_N0_S2 <=     O55_N0_S1  +  O55_N2_S1 ;
 logic signed [21:0] O55_N2_S2;		always @(posedge clk) O55_N2_S2 <=     O55_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O55_N0_S3;		always @(posedge clk) O55_N0_S3 <=     O55_N0_S2  +  O55_N2_S2 ;
 assign conv_mac_55 = O55_N0_S3;

logic signed [31:0] conv_mac_56;
logic signed [63:0] chainout_0_O56; 
logic signed [63:0] O56_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O56(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_56[7:0]),.ay(-9'sd1),.bx(input_fmap_56[15:8]),.by(-9'sd10),.cx(input_fmap_56[23:16]),.cy(-9'sd1),.dx(input_fmap_56[31:24]),.dy( 9'sd3),.chainin(63'd0),.result(O56_N0_S1),.chainout(chainout_0_O56));
logic signed [63:0] chainout_2_O56; 
logic signed [63:0] O56_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O56(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_56[39:32]),.ay( 9'sd21),.bx(input_fmap_56[47:40]),.by(-9'sd4),.cx(input_fmap_56[55:48]),.cy( 9'sd3),.dx(input_fmap_56[63:56]),.dy( 9'sd17),.chainin(63'd0),.result(O56_N2_S1),.chainout(chainout_2_O56));
logic signed [63:0] chainout_4_O56; 
logic signed [63:0] O56_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O56(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_56[71:64]),.ay(-9'sd3),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O56_N4_S1),.chainout(chainout_4_O56));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O56_N0_S2;		always @(posedge clk) O56_N0_S2 <=     O56_N0_S1  +  O56_N2_S1 ;
 logic signed [21:0] O56_N2_S2;		always @(posedge clk) O56_N2_S2 <=     O56_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O56_N0_S3;		always @(posedge clk) O56_N0_S3 <=     O56_N0_S2  +  O56_N2_S2 ;
 assign conv_mac_56 = O56_N0_S3;

logic signed [31:0] conv_mac_57;
logic signed [63:0] chainout_0_O57; 
logic signed [63:0] O57_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O57(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_57[7:0]),.ay(-9'sd4),.bx(input_fmap_57[15:8]),.by( 9'sd4),.cx(input_fmap_57[23:16]),.cy( 9'sd6),.dx(input_fmap_57[31:24]),.dy(-9'sd9),.chainin(63'd0),.result(O57_N0_S1),.chainout(chainout_0_O57));
logic signed [63:0] chainout_2_O57; 
logic signed [63:0] O57_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O57(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_57[39:32]),.ay( 9'sd39),.bx(input_fmap_57[47:40]),.by(-9'sd2),.cx(input_fmap_57[55:48]),.cy(-9'sd3),.dx(input_fmap_57[63:56]),.dy(-9'sd13),.chainin(63'd0),.result(O57_N2_S1),.chainout(chainout_2_O57));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O57_N0_S2;		always @(posedge clk) O57_N0_S2 <=     O57_N0_S1  +  O57_N2_S1 ;
 assign conv_mac_57 = O57_N0_S2;

logic signed [31:0] conv_mac_58;
logic signed [63:0] chainout_0_O58; 
logic signed [63:0] O58_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O58(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_58[7:0]),.ay(-9'sd1),.bx(input_fmap_58[15:8]),.by( 9'sd7),.cx(input_fmap_58[23:16]),.cy( 9'sd4),.dx(input_fmap_58[31:24]),.dy(-9'sd3),.chainin(63'd0),.result(O58_N0_S1),.chainout(chainout_0_O58));
logic signed [63:0] chainout_2_O58; 
logic signed [63:0] O58_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O58(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_58[39:32]),.ay( 9'sd27),.bx(input_fmap_58[55:48]),.by(-9'sd1),.cx(input_fmap_58[63:56]),.cy(-9'sd6),.dx(input_fmap_58[71:64]),.dy( 9'sd2),.chainin(63'd0),.result(O58_N2_S1),.chainout(chainout_2_O58));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O58_N0_S2;		always @(posedge clk) O58_N0_S2 <=     O58_N0_S1  +  O58_N2_S1 ;
 assign conv_mac_58 = O58_N0_S2;

logic signed [31:0] conv_mac_59;
logic signed [63:0] chainout_0_O59; 
logic signed [63:0] O59_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O59(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_59[7:0]),.ay(-9'sd3),.bx(input_fmap_59[15:8]),.by( 9'sd3),.cx(input_fmap_59[23:16]),.cy( 9'sd2),.dx(input_fmap_59[39:32]),.dy( 9'sd30),.chainin(63'd0),.result(O59_N0_S1),.chainout(chainout_0_O59));
logic signed [63:0] chainout_2_O59; 
logic signed [63:0] O59_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O59(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_59[47:40]),.ay(-9'sd3),.bx(input_fmap_59[55:48]),.by( 9'sd6),.cx(input_fmap_59[63:56]),.cy(-9'sd5),.dx(input_fmap_59[71:64]),.dy( 9'sd2),.chainin(63'd0),.result(O59_N2_S1),.chainout(chainout_2_O59));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O59_N0_S2;		always @(posedge clk) O59_N0_S2 <=     O59_N0_S1  +  O59_N2_S1 ;
 assign conv_mac_59 = O59_N0_S2;

logic signed [31:0] conv_mac_60;
logic signed [63:0] chainout_0_O60; 
logic signed [63:0] O60_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O60(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_60[7:0]),.ay( 9'sd5),.bx(input_fmap_60[15:8]),.by( 9'sd7),.cx(input_fmap_60[23:16]),.cy(-9'sd3),.dx(input_fmap_60[31:24]),.dy( 9'sd11),.chainin(63'd0),.result(O60_N0_S1),.chainout(chainout_0_O60));
logic signed [63:0] chainout_2_O60; 
logic signed [63:0] O60_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O60(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_60[39:32]),.ay(-9'sd27),.bx(input_fmap_60[47:40]),.by(-9'sd5),.cx(input_fmap_60[55:48]),.cy( 9'sd4),.dx(input_fmap_60[63:56]),.dy(-9'sd2),.chainin(63'd0),.result(O60_N2_S1),.chainout(chainout_2_O60));
logic signed [63:0] chainout_4_O60; 
logic signed [63:0] O60_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O60(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_60[71:64]),.ay(-9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O60_N4_S1),.chainout(chainout_4_O60));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O60_N0_S2;		always @(posedge clk) O60_N0_S2 <=     O60_N0_S1  +  O60_N2_S1 ;
 logic signed [21:0] O60_N2_S2;		always @(posedge clk) O60_N2_S2 <=     O60_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O60_N0_S3;		always @(posedge clk) O60_N0_S3 <=     O60_N0_S2  +  O60_N2_S2 ;
 assign conv_mac_60 = O60_N0_S3;

logic signed [31:0] conv_mac_61;
logic signed [63:0] chainout_0_O61; 
logic signed [63:0] O61_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O61(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_61[7:0]),.ay( 9'sd8),.bx(input_fmap_61[15:8]),.by( 9'sd1),.cx(input_fmap_61[23:16]),.cy( 9'sd3),.dx(input_fmap_61[31:24]),.dy( 9'sd11),.chainin(63'd0),.result(O61_N0_S1),.chainout(chainout_0_O61));
logic signed [63:0] chainout_2_O61; 
logic signed [63:0] O61_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O61(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_61[39:32]),.ay(-9'sd23),.bx(input_fmap_61[47:40]),.by(-9'sd9),.cx(input_fmap_61[55:48]),.cy( 9'sd4),.dx(input_fmap_61[63:56]),.dy(-9'sd11),.chainin(63'd0),.result(O61_N2_S1),.chainout(chainout_2_O61));
logic signed [63:0] chainout_4_O61; 
logic signed [63:0] O61_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O61(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_61[71:64]),.ay(-9'sd6),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O61_N4_S1),.chainout(chainout_4_O61));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O61_N0_S2;		always @(posedge clk) O61_N0_S2 <=     O61_N0_S1  +  O61_N2_S1 ;
 logic signed [21:0] O61_N2_S2;		always @(posedge clk) O61_N2_S2 <=     O61_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O61_N0_S3;		always @(posedge clk) O61_N0_S3 <=     O61_N0_S2  +  O61_N2_S2 ;
 assign conv_mac_61 = O61_N0_S3;

logic signed [31:0] conv_mac_62;
logic signed [63:0] chainout_0_O62; 
logic signed [63:0] O62_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O62(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_62[7:0]),.ay(-9'sd3),.bx(input_fmap_62[15:8]),.by( 9'sd9),.cx(input_fmap_62[23:16]),.cy( 9'sd8),.dx(input_fmap_62[31:24]),.dy(-9'sd5),.chainin(63'd0),.result(O62_N0_S1),.chainout(chainout_0_O62));
logic signed [63:0] chainout_2_O62; 
logic signed [63:0] O62_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O62(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_62[39:32]),.ay(-9'sd11),.bx(input_fmap_62[47:40]),.by( 9'sd14),.cx(input_fmap_62[55:48]),.cy(-9'sd6),.dx(input_fmap_62[63:56]),.dy(-9'sd2),.chainin(63'd0),.result(O62_N2_S1),.chainout(chainout_2_O62));
logic signed [63:0] chainout_4_O62; 
logic signed [63:0] O62_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O62(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_62[71:64]),.ay( 9'sd4),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O62_N4_S1),.chainout(chainout_4_O62));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O62_N0_S2;		always @(posedge clk) O62_N0_S2 <=     O62_N0_S1  +  O62_N2_S1 ;
 logic signed [21:0] O62_N2_S2;		always @(posedge clk) O62_N2_S2 <=     O62_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O62_N0_S3;		always @(posedge clk) O62_N0_S3 <=     O62_N0_S2  +  O62_N2_S2 ;
 assign conv_mac_62 = O62_N0_S3;

logic signed [31:0] conv_mac_63;
logic signed [63:0] chainout_0_O63; 
logic signed [63:0] O63_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O63(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_63[7:0]),.ay(-9'sd2),.bx(input_fmap_63[15:8]),.by(-9'sd7),.cx(input_fmap_63[23:16]),.cy(-9'sd6),.dx(input_fmap_63[31:24]),.dy(-9'sd3),.chainin(63'd0),.result(O63_N0_S1),.chainout(chainout_0_O63));
logic signed [63:0] chainout_2_O63; 
logic signed [63:0] O63_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O63(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_63[39:32]),.ay(-9'sd6),.bx(input_fmap_63[47:40]),.by(-9'sd3),.cx(input_fmap_63[55:48]),.cy( 9'sd1),.dx(input_fmap_63[63:56]),.dy(-9'sd8),.chainin(63'd0),.result(O63_N2_S1),.chainout(chainout_2_O63));
logic signed [63:0] chainout_4_O63; 
logic signed [63:0] O63_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O63(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_63[71:64]),.ay(-9'sd3),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O63_N4_S1),.chainout(chainout_4_O63));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O63_N0_S2;		always @(posedge clk) O63_N0_S2 <=     O63_N0_S1  +  O63_N2_S1 ;
 logic signed [21:0] O63_N2_S2;		always @(posedge clk) O63_N2_S2 <=     O63_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O63_N0_S3;		always @(posedge clk) O63_N0_S3 <=     O63_N0_S2  +  O63_N2_S2 ;
 assign conv_mac_63 = O63_N0_S3;

logic valid_D1;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D1<= 0 ;
	else valid_D1<=valid;
end
logic valid_D2;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D2<= 0 ;
	else valid_D2<=valid_D1;
end
logic valid_D3;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D3<= 0 ;
	else valid_D3<=valid_D2;
end
logic valid_D4;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D4<= 0 ;
	else valid_D4<=valid_D3;
end
always_ff @(posedge clk) begin
	if (rstn == 0) ready <= 0 ;
	else ready <=valid_D4;
end
logic [31:0] bias_add_0;
assign bias_add_0 = conv_mac_0 + 6'd22;
logic [31:0] bias_add_1;
assign bias_add_1 = conv_mac_1 - 3'd2;
logic [31:0] bias_add_2;
assign bias_add_2 = conv_mac_2 + 7'd63;
logic [31:0] bias_add_3;
assign bias_add_3 = conv_mac_3;
logic [31:0] bias_add_4;
assign bias_add_4 = conv_mac_4 + 7'd39;
logic [31:0] bias_add_5;
assign bias_add_5 = conv_mac_5 + 6'd26;
logic [31:0] bias_add_6;
assign bias_add_6 = conv_mac_6 + 6'd18;
logic [31:0] bias_add_7;
assign bias_add_7 = conv_mac_7 + 7'd42;
logic [31:0] bias_add_8;
assign bias_add_8 = conv_mac_8 + 7'd59;
logic [31:0] bias_add_9;
assign bias_add_9 = conv_mac_9 + 5'd8;
logic [31:0] bias_add_10;
assign bias_add_10 = conv_mac_10 + 2'd1;
logic [31:0] bias_add_11;
assign bias_add_11 = conv_mac_11 + 4'd6;
logic [31:0] bias_add_12;
assign bias_add_12 = conv_mac_12 - 5'd11;
logic [31:0] bias_add_13;
assign bias_add_13 = conv_mac_13 + 6'd20;
logic [31:0] bias_add_14;
assign bias_add_14 = conv_mac_14 - 5'd10;
logic [31:0] bias_add_15;
assign bias_add_15 = conv_mac_15 + 5'd11;
logic [31:0] bias_add_16;
assign bias_add_16 = conv_mac_16 + 3'd3;
logic [31:0] bias_add_17;
assign bias_add_17 = conv_mac_17 + 5'd8;
logic [31:0] bias_add_18;
assign bias_add_18 = conv_mac_18 - 4'd6;
logic [31:0] bias_add_19;
assign bias_add_19 = conv_mac_19 + 5'd12;
logic [31:0] bias_add_20;
assign bias_add_20 = conv_mac_20 + 6'd26;
logic [31:0] bias_add_21;
assign bias_add_21 = conv_mac_21 - 5'd13;
logic [31:0] bias_add_22;
assign bias_add_22 = conv_mac_22 - 5'd8;
logic [31:0] bias_add_23;
assign bias_add_23 = conv_mac_23 + 5'd9;
logic [31:0] bias_add_24;
assign bias_add_24 = conv_mac_24 + 6'd25;
logic [31:0] bias_add_25;
assign bias_add_25 = conv_mac_25 + 6'd18;
logic [31:0] bias_add_26;
assign bias_add_26 = conv_mac_26 + 5'd15;
logic [31:0] bias_add_27;
assign bias_add_27 = conv_mac_27 + 5'd12;
logic [31:0] bias_add_28;
assign bias_add_28 = conv_mac_28 - 5'd11;
logic [31:0] bias_add_29;
assign bias_add_29 = conv_mac_29 + 4'd4;
logic [31:0] bias_add_30;
assign bias_add_30 = conv_mac_30 - 3'd3;
logic [31:0] bias_add_31;
assign bias_add_31 = conv_mac_31 - 3'd2;
logic [31:0] bias_add_32;
assign bias_add_32 = conv_mac_32 + 4'd6;
logic [31:0] bias_add_33;
assign bias_add_33 = conv_mac_33 + 7'd35;
logic [31:0] bias_add_34;
assign bias_add_34 = conv_mac_34 + 4'd6;
logic [31:0] bias_add_35;
assign bias_add_35 = conv_mac_35 - 5'd9;
logic [31:0] bias_add_36;
assign bias_add_36 = conv_mac_36 + 5'd13;
logic [31:0] bias_add_37;
assign bias_add_37 = conv_mac_37 + 7'd42;
logic [31:0] bias_add_38;
assign bias_add_38 = conv_mac_38 + 4'd6;
logic [31:0] bias_add_39;
assign bias_add_39 = conv_mac_39 - 2'd1;
logic [31:0] bias_add_40;
assign bias_add_40 = conv_mac_40 - 2'd1;
logic [31:0] bias_add_41;
assign bias_add_41 = conv_mac_41 - 6'd18;
logic [31:0] bias_add_42;
assign bias_add_42 = conv_mac_42 - 5'd13;
logic [31:0] bias_add_43;
assign bias_add_43 = conv_mac_43 - 6'd17;
logic [31:0] bias_add_44;
assign bias_add_44 = conv_mac_44 - 5'd12;
logic [31:0] bias_add_45;
assign bias_add_45 = conv_mac_45 + 6'd29;
logic [31:0] bias_add_46;
assign bias_add_46 = conv_mac_46 + 4'd6;
logic [31:0] bias_add_47;
assign bias_add_47 = conv_mac_47 + 5'd10;
logic [31:0] bias_add_48;
assign bias_add_48 = conv_mac_48 + 6'd22;
logic [31:0] bias_add_49;
assign bias_add_49 = conv_mac_49 + 5'd8;
logic [31:0] bias_add_50;
assign bias_add_50 = conv_mac_50 + 6'd30;
logic [31:0] bias_add_51;
assign bias_add_51 = conv_mac_51 - 4'd4;
logic [31:0] bias_add_52;
assign bias_add_52 = conv_mac_52 - 3'd2;
logic [31:0] bias_add_53;
assign bias_add_53 = conv_mac_53 + 6'd26;
logic [31:0] bias_add_54;
assign bias_add_54 = conv_mac_54 - 3'd3;
logic [31:0] bias_add_55;
assign bias_add_55 = conv_mac_55 + 3'd2;
logic [31:0] bias_add_56;
assign bias_add_56 = conv_mac_56 - 2'd1;
logic [31:0] bias_add_57;
assign bias_add_57 = conv_mac_57 + 5'd12;
logic [31:0] bias_add_58;
assign bias_add_58 = conv_mac_58 - 2'd1;
logic [31:0] bias_add_59;
assign bias_add_59 = conv_mac_59 + 3'd2;
logic [31:0] bias_add_60;
assign bias_add_60 = conv_mac_60 + 6'd24;
logic [31:0] bias_add_61;
assign bias_add_61 = conv_mac_61 + 7'd40;
logic [31:0] bias_add_62;
assign bias_add_62 = conv_mac_62 + 3'd3;
logic [31:0] bias_add_63;
assign bias_add_63 = conv_mac_63 + 6'd19;

logic [7:0] relu_0;
assign relu_0[7:0] = (bias_add_0[31]==0) ? ((bias_add_0<3'd6) ? {{bias_add_0[31],bias_add_0[10:4]}} :'d6) : '0;
logic [7:0] relu_1;
assign relu_1[7:0] = (bias_add_1[31]==0) ? ((bias_add_1<3'd6) ? {{bias_add_1[31],bias_add_1[10:4]}} :'d6) : '0;
logic [7:0] relu_2;
assign relu_2[7:0] = (bias_add_2[31]==0) ? ((bias_add_2<3'd6) ? {{bias_add_2[31],bias_add_2[10:4]}} :'d6) : '0;
logic [7:0] relu_3;
assign relu_3[7:0] = (bias_add_3[31]==0) ? ((bias_add_3<3'd6) ? {{bias_add_3[31],bias_add_3[10:4]}} :'d6) : '0;
logic [7:0] relu_4;
assign relu_4[7:0] = (bias_add_4[31]==0) ? ((bias_add_4<3'd6) ? {{bias_add_4[31],bias_add_4[10:4]}} :'d6) : '0;
logic [7:0] relu_5;
assign relu_5[7:0] = (bias_add_5[31]==0) ? ((bias_add_5<3'd6) ? {{bias_add_5[31],bias_add_5[10:4]}} :'d6) : '0;
logic [7:0] relu_6;
assign relu_6[7:0] = (bias_add_6[31]==0) ? ((bias_add_6<3'd6) ? {{bias_add_6[31],bias_add_6[10:4]}} :'d6) : '0;
logic [7:0] relu_7;
assign relu_7[7:0] = (bias_add_7[31]==0) ? ((bias_add_7<3'd6) ? {{bias_add_7[31],bias_add_7[10:4]}} :'d6) : '0;
logic [7:0] relu_8;
assign relu_8[7:0] = (bias_add_8[31]==0) ? ((bias_add_8<3'd6) ? {{bias_add_8[31],bias_add_8[10:4]}} :'d6) : '0;
logic [7:0] relu_9;
assign relu_9[7:0] = (bias_add_9[31]==0) ? ((bias_add_9<3'd6) ? {{bias_add_9[31],bias_add_9[10:4]}} :'d6) : '0;
logic [7:0] relu_10;
assign relu_10[7:0] = (bias_add_10[31]==0) ? ((bias_add_10<3'd6) ? {{bias_add_10[31],bias_add_10[10:4]}} :'d6) : '0;
logic [7:0] relu_11;
assign relu_11[7:0] = (bias_add_11[31]==0) ? ((bias_add_11<3'd6) ? {{bias_add_11[31],bias_add_11[10:4]}} :'d6) : '0;
logic [7:0] relu_12;
assign relu_12[7:0] = (bias_add_12[31]==0) ? ((bias_add_12<3'd6) ? {{bias_add_12[31],bias_add_12[10:4]}} :'d6) : '0;
logic [7:0] relu_13;
assign relu_13[7:0] = (bias_add_13[31]==0) ? ((bias_add_13<3'd6) ? {{bias_add_13[31],bias_add_13[10:4]}} :'d6) : '0;
logic [7:0] relu_14;
assign relu_14[7:0] = (bias_add_14[31]==0) ? ((bias_add_14<3'd6) ? {{bias_add_14[31],bias_add_14[10:4]}} :'d6) : '0;
logic [7:0] relu_15;
assign relu_15[7:0] = (bias_add_15[31]==0) ? ((bias_add_15<3'd6) ? {{bias_add_15[31],bias_add_15[10:4]}} :'d6) : '0;
logic [7:0] relu_16;
assign relu_16[7:0] = (bias_add_16[31]==0) ? ((bias_add_16<3'd6) ? {{bias_add_16[31],bias_add_16[10:4]}} :'d6) : '0;
logic [7:0] relu_17;
assign relu_17[7:0] = (bias_add_17[31]==0) ? ((bias_add_17<3'd6) ? {{bias_add_17[31],bias_add_17[10:4]}} :'d6) : '0;
logic [7:0] relu_18;
assign relu_18[7:0] = (bias_add_18[31]==0) ? ((bias_add_18<3'd6) ? {{bias_add_18[31],bias_add_18[10:4]}} :'d6) : '0;
logic [7:0] relu_19;
assign relu_19[7:0] = (bias_add_19[31]==0) ? ((bias_add_19<3'd6) ? {{bias_add_19[31],bias_add_19[10:4]}} :'d6) : '0;
logic [7:0] relu_20;
assign relu_20[7:0] = (bias_add_20[31]==0) ? ((bias_add_20<3'd6) ? {{bias_add_20[31],bias_add_20[10:4]}} :'d6) : '0;
logic [7:0] relu_21;
assign relu_21[7:0] = (bias_add_21[31]==0) ? ((bias_add_21<3'd6) ? {{bias_add_21[31],bias_add_21[10:4]}} :'d6) : '0;
logic [7:0] relu_22;
assign relu_22[7:0] = (bias_add_22[31]==0) ? ((bias_add_22<3'd6) ? {{bias_add_22[31],bias_add_22[10:4]}} :'d6) : '0;
logic [7:0] relu_23;
assign relu_23[7:0] = (bias_add_23[31]==0) ? ((bias_add_23<3'd6) ? {{bias_add_23[31],bias_add_23[10:4]}} :'d6) : '0;
logic [7:0] relu_24;
assign relu_24[7:0] = (bias_add_24[31]==0) ? ((bias_add_24<3'd6) ? {{bias_add_24[31],bias_add_24[10:4]}} :'d6) : '0;
logic [7:0] relu_25;
assign relu_25[7:0] = (bias_add_25[31]==0) ? ((bias_add_25<3'd6) ? {{bias_add_25[31],bias_add_25[10:4]}} :'d6) : '0;
logic [7:0] relu_26;
assign relu_26[7:0] = (bias_add_26[31]==0) ? ((bias_add_26<3'd6) ? {{bias_add_26[31],bias_add_26[10:4]}} :'d6) : '0;
logic [7:0] relu_27;
assign relu_27[7:0] = (bias_add_27[31]==0) ? ((bias_add_27<3'd6) ? {{bias_add_27[31],bias_add_27[10:4]}} :'d6) : '0;
logic [7:0] relu_28;
assign relu_28[7:0] = (bias_add_28[31]==0) ? ((bias_add_28<3'd6) ? {{bias_add_28[31],bias_add_28[10:4]}} :'d6) : '0;
logic [7:0] relu_29;
assign relu_29[7:0] = (bias_add_29[31]==0) ? ((bias_add_29<3'd6) ? {{bias_add_29[31],bias_add_29[10:4]}} :'d6) : '0;
logic [7:0] relu_30;
assign relu_30[7:0] = (bias_add_30[31]==0) ? ((bias_add_30<3'd6) ? {{bias_add_30[31],bias_add_30[10:4]}} :'d6) : '0;
logic [7:0] relu_31;
assign relu_31[7:0] = (bias_add_31[31]==0) ? ((bias_add_31<3'd6) ? {{bias_add_31[31],bias_add_31[10:4]}} :'d6) : '0;
logic [7:0] relu_32;
assign relu_32[7:0] = (bias_add_32[31]==0) ? ((bias_add_32<3'd6) ? {{bias_add_32[31],bias_add_32[10:4]}} :'d6) : '0;
logic [7:0] relu_33;
assign relu_33[7:0] = (bias_add_33[31]==0) ? ((bias_add_33<3'd6) ? {{bias_add_33[31],bias_add_33[10:4]}} :'d6) : '0;
logic [7:0] relu_34;
assign relu_34[7:0] = (bias_add_34[31]==0) ? ((bias_add_34<3'd6) ? {{bias_add_34[31],bias_add_34[10:4]}} :'d6) : '0;
logic [7:0] relu_35;
assign relu_35[7:0] = (bias_add_35[31]==0) ? ((bias_add_35<3'd6) ? {{bias_add_35[31],bias_add_35[10:4]}} :'d6) : '0;
logic [7:0] relu_36;
assign relu_36[7:0] = (bias_add_36[31]==0) ? ((bias_add_36<3'd6) ? {{bias_add_36[31],bias_add_36[10:4]}} :'d6) : '0;
logic [7:0] relu_37;
assign relu_37[7:0] = (bias_add_37[31]==0) ? ((bias_add_37<3'd6) ? {{bias_add_37[31],bias_add_37[10:4]}} :'d6) : '0;
logic [7:0] relu_38;
assign relu_38[7:0] = (bias_add_38[31]==0) ? ((bias_add_38<3'd6) ? {{bias_add_38[31],bias_add_38[10:4]}} :'d6) : '0;
logic [7:0] relu_39;
assign relu_39[7:0] = (bias_add_39[31]==0) ? ((bias_add_39<3'd6) ? {{bias_add_39[31],bias_add_39[10:4]}} :'d6) : '0;
logic [7:0] relu_40;
assign relu_40[7:0] = (bias_add_40[31]==0) ? ((bias_add_40<3'd6) ? {{bias_add_40[31],bias_add_40[10:4]}} :'d6) : '0;
logic [7:0] relu_41;
assign relu_41[7:0] = (bias_add_41[31]==0) ? ((bias_add_41<3'd6) ? {{bias_add_41[31],bias_add_41[10:4]}} :'d6) : '0;
logic [7:0] relu_42;
assign relu_42[7:0] = (bias_add_42[31]==0) ? ((bias_add_42<3'd6) ? {{bias_add_42[31],bias_add_42[10:4]}} :'d6) : '0;
logic [7:0] relu_43;
assign relu_43[7:0] = (bias_add_43[31]==0) ? ((bias_add_43<3'd6) ? {{bias_add_43[31],bias_add_43[10:4]}} :'d6) : '0;
logic [7:0] relu_44;
assign relu_44[7:0] = (bias_add_44[31]==0) ? ((bias_add_44<3'd6) ? {{bias_add_44[31],bias_add_44[10:4]}} :'d6) : '0;
logic [7:0] relu_45;
assign relu_45[7:0] = (bias_add_45[31]==0) ? ((bias_add_45<3'd6) ? {{bias_add_45[31],bias_add_45[10:4]}} :'d6) : '0;
logic [7:0] relu_46;
assign relu_46[7:0] = (bias_add_46[31]==0) ? ((bias_add_46<3'd6) ? {{bias_add_46[31],bias_add_46[10:4]}} :'d6) : '0;
logic [7:0] relu_47;
assign relu_47[7:0] = (bias_add_47[31]==0) ? ((bias_add_47<3'd6) ? {{bias_add_47[31],bias_add_47[10:4]}} :'d6) : '0;
logic [7:0] relu_48;
assign relu_48[7:0] = (bias_add_48[31]==0) ? ((bias_add_48<3'd6) ? {{bias_add_48[31],bias_add_48[10:4]}} :'d6) : '0;
logic [7:0] relu_49;
assign relu_49[7:0] = (bias_add_49[31]==0) ? ((bias_add_49<3'd6) ? {{bias_add_49[31],bias_add_49[10:4]}} :'d6) : '0;
logic [7:0] relu_50;
assign relu_50[7:0] = (bias_add_50[31]==0) ? ((bias_add_50<3'd6) ? {{bias_add_50[31],bias_add_50[10:4]}} :'d6) : '0;
logic [7:0] relu_51;
assign relu_51[7:0] = (bias_add_51[31]==0) ? ((bias_add_51<3'd6) ? {{bias_add_51[31],bias_add_51[10:4]}} :'d6) : '0;
logic [7:0] relu_52;
assign relu_52[7:0] = (bias_add_52[31]==0) ? ((bias_add_52<3'd6) ? {{bias_add_52[31],bias_add_52[10:4]}} :'d6) : '0;
logic [7:0] relu_53;
assign relu_53[7:0] = (bias_add_53[31]==0) ? ((bias_add_53<3'd6) ? {{bias_add_53[31],bias_add_53[10:4]}} :'d6) : '0;
logic [7:0] relu_54;
assign relu_54[7:0] = (bias_add_54[31]==0) ? ((bias_add_54<3'd6) ? {{bias_add_54[31],bias_add_54[10:4]}} :'d6) : '0;
logic [7:0] relu_55;
assign relu_55[7:0] = (bias_add_55[31]==0) ? ((bias_add_55<3'd6) ? {{bias_add_55[31],bias_add_55[10:4]}} :'d6) : '0;
logic [7:0] relu_56;
assign relu_56[7:0] = (bias_add_56[31]==0) ? ((bias_add_56<3'd6) ? {{bias_add_56[31],bias_add_56[10:4]}} :'d6) : '0;
logic [7:0] relu_57;
assign relu_57[7:0] = (bias_add_57[31]==0) ? ((bias_add_57<3'd6) ? {{bias_add_57[31],bias_add_57[10:4]}} :'d6) : '0;
logic [7:0] relu_58;
assign relu_58[7:0] = (bias_add_58[31]==0) ? ((bias_add_58<3'd6) ? {{bias_add_58[31],bias_add_58[10:4]}} :'d6) : '0;
logic [7:0] relu_59;
assign relu_59[7:0] = (bias_add_59[31]==0) ? ((bias_add_59<3'd6) ? {{bias_add_59[31],bias_add_59[10:4]}} :'d6) : '0;
logic [7:0] relu_60;
assign relu_60[7:0] = (bias_add_60[31]==0) ? ((bias_add_60<3'd6) ? {{bias_add_60[31],bias_add_60[10:4]}} :'d6) : '0;
logic [7:0] relu_61;
assign relu_61[7:0] = (bias_add_61[31]==0) ? ((bias_add_61<3'd6) ? {{bias_add_61[31],bias_add_61[10:4]}} :'d6) : '0;
logic [7:0] relu_62;
assign relu_62[7:0] = (bias_add_62[31]==0) ? ((bias_add_62<3'd6) ? {{bias_add_62[31],bias_add_62[10:4]}} :'d6) : '0;
logic [7:0] relu_63;
assign relu_63[7:0] = (bias_add_63[31]==0) ? ((bias_add_63<3'd6) ? {{bias_add_63[31],bias_add_63[10:4]}} :'d6) : '0;

assign output_act = {
	relu_63,
	relu_62,
	relu_61,
	relu_60,
	relu_59,
	relu_58,
	relu_57,
	relu_56,
	relu_55,
	relu_54,
	relu_53,
	relu_52,
	relu_51,
	relu_50,
	relu_49,
	relu_48,
	relu_47,
	relu_46,
	relu_45,
	relu_44,
	relu_43,
	relu_42,
	relu_41,
	relu_40,
	relu_39,
	relu_38,
	relu_37,
	relu_36,
	relu_35,
	relu_34,
	relu_33,
	relu_32,
	relu_31,
	relu_30,
	relu_29,
	relu_28,
	relu_27,
	relu_26,
	relu_25,
	relu_24,
	relu_23,
	relu_22,
	relu_21,
	relu_20,
	relu_19,
	relu_18,
	relu_17,
	relu_16,
	relu_15,
	relu_14,
	relu_13,
	relu_12,
	relu_11,
	relu_10,
	relu_9,
	relu_8,
	relu_7,
	relu_6,
	relu_5,
	relu_4,
	relu_3,
	relu_2,
	relu_1,
	relu_0
};

endmodule
module conv1_pw (
    input logic clk,
    input logic rstn,
    input logic valid,
    input logic [64-1:0] input_act,
    output logic [64-1:0] output_act,
    output logic ready
);
logic we;
logic [8:0] zero_number; 
assign zero_number = 9'd0; 
//1
logic [64-1:0] input_act_ff ;
always_ff @(posedge clk) begin
    if (rstn == 0) begin
        input_act_ff <= '0;
      //  ready <= '0;
    end
    else begin
        input_act_ff <= input_act;
     //   ready <= valid;
    end
end
logic [7:0] input_fmap_0;
assign input_fmap_0 = input_act_ff[7:0];
logic [7:0] input_fmap_1;
assign input_fmap_1 = input_act_ff[15:8];
logic [7:0] input_fmap_2;
assign input_fmap_2 = input_act_ff[23:16];
logic [7:0] input_fmap_3;
assign input_fmap_3 = input_act_ff[31:24];
logic [7:0] input_fmap_4;
assign input_fmap_4 = input_act_ff[39:32];
logic [7:0] input_fmap_5;
assign input_fmap_5 = input_act_ff[47:40];
logic [7:0] input_fmap_6;
assign input_fmap_6 = input_act_ff[55:48];
logic [7:0] input_fmap_7;
assign input_fmap_7 = input_act_ff[63:56];

logic [11-1:0] O0_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv1_pw_O0_I0_R0_C03_rom_inst (.q(O0_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O0_I0_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_pw_O0_I0_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv1_pw_O0_I0_R0_C03_rom_inst (.q(O0_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [10-1:0] O0_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv1_pw_O0_I6_R0_C01_rom_inst (.q(O0_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I6_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O0_I6_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_pw_O0_I6_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv1_pw_O0_I6_R0_C01_rom_inst (.q(O0_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [12-1:0] O0_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv1_pw_O0_I7_R0_C04_rom_inst (.q(O0_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I7_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O0_I7_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_pw_O0_I7_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv1_pw_O0_I7_R0_C04_rom_inst (.q(O0_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [10-1:0] O1_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv1_pw_O1_I2_R0_C01_rom_inst (.q(O1_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O1_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_pw_O1_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv1_pw_O1_I2_R0_C01_rom_inst (.q(O1_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [10-1:0] O1_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv1_pw_O1_I4_R0_C01_rom_inst (.q(O1_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I4_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O1_I4_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_pw_O1_I4_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv1_pw_O1_I4_R0_C01_rom_inst (.q(O1_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [12-1:0] O1_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv1_pw_O1_I5_R0_C04_rom_inst (.q(O1_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I5_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O1_I5_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_pw_O1_I5_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv1_pw_O1_I5_R0_C04_rom_inst (.q(O1_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [10-1:0] O1_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv1_pw_O1_I6_R0_C01_rom_inst (.q(O1_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I6_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O1_I6_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_pw_O1_I6_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv1_pw_O1_I6_R0_C01_rom_inst (.q(O1_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [10-1:0] O1_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv1_pw_O1_I7_R0_C01_rom_inst (.q(O1_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I7_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O1_I7_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_pw_O1_I7_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv1_pw_O1_I7_R0_C01_rom_inst (.q(O1_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [13-1:0] O2_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv1_pw_O2_I1_R0_C012_rom_inst (.q(O2_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O2_I1_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O2_I1_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_pw_O2_I1_R0_C012_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv1_pw_O2_I1_R0_C012_rom_inst (.q(O2_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [10-1:0] O3_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv1_pw_O3_I3_R0_C01_rom_inst (.q(O3_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O3_I3_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_pw_O3_I3_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv1_pw_O3_I3_R0_C01_rom_inst (.q(O3_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [11-1:0] O3_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv1_pw_O3_I5_R0_C03_rom_inst (.q(O3_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I5_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O3_I5_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_pw_O3_I5_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv1_pw_O3_I5_R0_C03_rom_inst (.q(O3_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [10-1:0] O4_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv1_pw_O4_I0_R0_C01_rom_inst (.q(O4_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I0_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I0_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_pw_O4_I0_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv1_pw_O4_I0_R0_C01_rom_inst (.q(O4_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [12-1:0] O4_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv1_pw_O4_I1_R0_C06_rom_inst (.q(O4_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I1_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O4_I1_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_pw_O4_I1_R0_C06_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv1_pw_O4_I1_R0_C06_rom_inst (.q(O4_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [10-1:0] O4_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv1_pw_O4_I2_R0_C01_rom_inst (.q(O4_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_pw_O4_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv1_pw_O4_I2_R0_C01_rom_inst (.q(O4_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [10-1:0] O4_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv1_pw_O4_I3_R0_C01_rom_inst (.q(O4_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I3_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I3_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_pw_O4_I3_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv1_pw_O4_I3_R0_C01_rom_inst (.q(O4_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [11-1:0] O4_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv1_pw_O4_I4_R0_C02_rom_inst (.q(O4_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O4_I4_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_pw_O4_I4_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv1_pw_O4_I4_R0_C02_rom_inst (.q(O4_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [10-1:0] O4_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv1_pw_O4_I5_R0_C01_rom_inst (.q(O4_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I5_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I5_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_pw_O4_I5_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv1_pw_O4_I5_R0_C01_rom_inst (.q(O4_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [10-1:0] O4_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv1_pw_O4_I6_R0_C01_rom_inst (.q(O4_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I6_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I6_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_pw_O4_I6_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv1_pw_O4_I6_R0_C01_rom_inst (.q(O4_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [10-1:0] O4_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv1_pw_O4_I7_R0_C01_rom_inst (.q(O4_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I7_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I7_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_pw_O4_I7_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv1_pw_O4_I7_R0_C01_rom_inst (.q(O4_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [13-1:0] O5_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv1_pw_O5_I0_R0_C011_rom_inst (.q(O5_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I0_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O5_I0_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_pw_O5_I0_R0_C011_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv1_pw_O5_I0_R0_C011_rom_inst (.q(O5_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [10-1:0] O5_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv1_pw_O5_I2_R0_C01_rom_inst (.q(O5_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_pw_O5_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv1_pw_O5_I2_R0_C01_rom_inst (.q(O5_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [10-1:0] O5_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv1_pw_O5_I3_R0_C01_rom_inst (.q(O5_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I3_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I3_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_pw_O5_I3_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv1_pw_O5_I3_R0_C01_rom_inst (.q(O5_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [10-1:0] O5_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv1_pw_O5_I4_R0_C01_rom_inst (.q(O5_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I4_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I4_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_pw_O5_I4_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv1_pw_O5_I4_R0_C01_rom_inst (.q(O5_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [11-1:0] O5_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv1_pw_O5_I5_R0_C02_rom_inst (.q(O5_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O5_I5_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_pw_O5_I5_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv1_pw_O5_I5_R0_C02_rom_inst (.q(O5_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [10-1:0] O5_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv1_pw_O5_I6_R0_C01_rom_inst (.q(O5_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I6_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I6_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_pw_O5_I6_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv1_pw_O5_I6_R0_C01_rom_inst (.q(O5_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [11-1:0] O5_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv1_pw_O5_I7_R0_C02_rom_inst (.q(O5_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I7_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O5_I7_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_pw_O5_I7_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv1_pw_O5_I7_R0_C02_rom_inst (.q(O5_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [11-1:0] O6_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv1_pw_O6_I0_R0_C02_rom_inst (.q(O6_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I0_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O6_I0_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_pw_O6_I0_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv1_pw_O6_I0_R0_C02_rom_inst (.q(O6_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [10-1:0] O6_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv1_pw_O6_I2_R0_C01_rom_inst (.q(O6_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O6_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_pw_O6_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv1_pw_O6_I2_R0_C01_rom_inst (.q(O6_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [12-1:0] O6_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv1_pw_O6_I6_R0_C05_rom_inst (.q(O6_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O6_I6_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_pw_O6_I6_R0_C05_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv1_pw_O6_I6_R0_C05_rom_inst (.q(O6_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [10-1:0] O6_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv1_pw_O6_I7_R0_C01_rom_inst (.q(O6_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I7_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O6_I7_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_pw_O6_I7_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv1_pw_O6_I7_R0_C01_rom_inst (.q(O6_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [10-1:0] O7_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv1_pw_O7_I0_R0_C01_rom_inst (.q(O7_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I0_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O7_I0_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_pw_O7_I0_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv1_pw_O7_I0_R0_C01_rom_inst (.q(O7_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [13-1:0] O7_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv1_pw_O7_I1_R0_C010_rom_inst (.q(O7_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I1_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O7_I1_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_pw_O7_I1_R0_C010_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv1_pw_O7_I1_R0_C010_rom_inst (.q(O7_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [11-1:0] O7_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv1_pw_O7_I2_R0_C02_rom_inst (.q(O7_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I2_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O7_I2_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv1_pw_O7_I2_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv1_pw_O7_I2_R0_C02_rom_inst (.q(O7_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic signed [31:0] conv_mac_0;
logic signed [31:0] O0_N0_S0;		always @(posedge clk) O0_N0_S0 <=     O0_I0_R0_C0_SM1   +  O0_I6_R0_C0_SM1  ;
 logic signed [31:0] O0_N2_S0;		always @(posedge clk) O0_N2_S0 <=     O0_I7_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O0_N0_S1;		always @(posedge clk) O0_N0_S1 <=     O0_N0_S0  +  O0_N2_S0 ;
 assign conv_mac_0 = O0_N0_S1;

logic signed [31:0] conv_mac_1;
logic signed [31:0] O1_N0_S0;		always @(posedge clk) O1_N0_S0 <=     O1_I2_R0_C0_SM1   +  O1_I4_R0_C0_SM1  ;
 logic signed [31:0] O1_N2_S0;		always @(posedge clk) O1_N2_S0 <=     O1_I5_R0_C0_SM1   +  O1_I6_R0_C0_SM1  ;
 logic signed [31:0] O1_N4_S0;		always @(posedge clk) O1_N4_S0 <=     O1_I7_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O1_N0_S1;		always @(posedge clk) O1_N0_S1 <=     O1_N0_S0  +  O1_N2_S0 ;
 logic signed [31:0] O1_N2_S1;		always @(posedge clk) O1_N2_S1 <=     O1_N4_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O1_N0_S2;		always @(posedge clk) O1_N0_S2 <=     O1_N0_S1  +  O1_N2_S1 ;
 assign conv_mac_1 = O1_N0_S2;

logic signed [31:0] conv_mac_2;
logic signed [31:0] O2_N0_S0;		always @(posedge clk) O2_N0_S0 <=     O2_I1_R0_C0_SM1      ;
 assign conv_mac_2 = O2_N0_S0;

logic signed [31:0] conv_mac_3;
logic signed [31:0] O3_N0_S0;		always @(posedge clk) O3_N0_S0 <=     O3_I3_R0_C0_SM1   +  O3_I5_R0_C0_SM1  ;
 assign conv_mac_3 = O3_N0_S0;

logic signed [31:0] conv_mac_4;
logic signed [31:0] O4_N0_S0;		always @(posedge clk) O4_N0_S0 <=     O4_I0_R0_C0_SM1   +  O4_I1_R0_C0_SM1  ;
 logic signed [31:0] O4_N2_S0;		always @(posedge clk) O4_N2_S0 <=     O4_I2_R0_C0_SM1   +  O4_I3_R0_C0_SM1  ;
 logic signed [31:0] O4_N4_S0;		always @(posedge clk) O4_N4_S0 <=     O4_I4_R0_C0_SM1   +  O4_I5_R0_C0_SM1  ;
 logic signed [31:0] O4_N6_S0;		always @(posedge clk) O4_N6_S0 <=     O4_I6_R0_C0_SM1   +  O4_I7_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O4_N0_S1;		always @(posedge clk) O4_N0_S1 <=     O4_N0_S0  +  O4_N2_S0 ;
 logic signed [31:0] O4_N2_S1;		always @(posedge clk) O4_N2_S1 <=     O4_N4_S0  +  O4_N6_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O4_N0_S2;		always @(posedge clk) O4_N0_S2 <=     O4_N0_S1  +  O4_N2_S1 ;
 assign conv_mac_4 = O4_N0_S2;

logic signed [31:0] conv_mac_5;
logic signed [31:0] O5_N0_S0;		always @(posedge clk) O5_N0_S0 <=     O5_I0_R0_C0_SM1   +  O5_I2_R0_C0_SM1  ;
 logic signed [31:0] O5_N2_S0;		always @(posedge clk) O5_N2_S0 <=     O5_I3_R0_C0_SM1   +  O5_I4_R0_C0_SM1  ;
 logic signed [31:0] O5_N4_S0;		always @(posedge clk) O5_N4_S0 <=     O5_I5_R0_C0_SM1   +  O5_I6_R0_C0_SM1  ;
 logic signed [31:0] O5_N6_S0;		always @(posedge clk) O5_N6_S0 <=     O5_I7_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O5_N0_S1;		always @(posedge clk) O5_N0_S1 <=     O5_N0_S0  +  O5_N2_S0 ;
 logic signed [31:0] O5_N2_S1;		always @(posedge clk) O5_N2_S1 <=     O5_N4_S0  +  O5_N6_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O5_N0_S2;		always @(posedge clk) O5_N0_S2 <=     O5_N0_S1  +  O5_N2_S1 ;
 assign conv_mac_5 = O5_N0_S2;

logic signed [31:0] conv_mac_6;
logic signed [31:0] O6_N0_S0;		always @(posedge clk) O6_N0_S0 <=     O6_I0_R0_C0_SM1   +  O6_I2_R0_C0_SM1  ;
 logic signed [31:0] O6_N2_S0;		always @(posedge clk) O6_N2_S0 <=     O6_I6_R0_C0_SM1   +  O6_I7_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O6_N0_S1;		always @(posedge clk) O6_N0_S1 <=     O6_N0_S0  +  O6_N2_S0 ;
 assign conv_mac_6 = O6_N0_S1;

logic signed [31:0] conv_mac_7;
logic signed [31:0] O7_N0_S0;		always @(posedge clk) O7_N0_S0 <=     O7_I0_R0_C0_SM1   +  O7_I1_R0_C0_SM1  ;
 logic signed [31:0] O7_N2_S0;		always @(posedge clk) O7_N2_S0 <=     O7_I2_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O7_N0_S1;		always @(posedge clk) O7_N0_S1 <=     O7_N0_S0  +  O7_N2_S0 ;
 assign conv_mac_7 = O7_N0_S1;

logic valid_D1;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D1<= 0 ;
	else valid_D1<=valid;
end
logic valid_D2;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D2<= 0 ;
	else valid_D2<=valid_D1;
end
logic valid_D3;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D3<= 0 ;
	else valid_D3<=valid_D2;
end
logic valid_D4;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D4<= 0 ;
	else valid_D4<=valid_D3;
end
always_ff @(posedge clk) begin
	if (rstn == 0) ready <= 0 ;
	else ready <=valid_D4;
end
logic [31:0] bias_add_0;
assign bias_add_0 = conv_mac_0 + 6'd22;
logic [31:0] bias_add_1;
assign bias_add_1 = conv_mac_1 + 7'd42;
logic [31:0] bias_add_2;
assign bias_add_2 = conv_mac_2 - 4'd7;
logic [31:0] bias_add_3;
assign bias_add_3 = conv_mac_3 + 6'd24;
logic [31:0] bias_add_4;
assign bias_add_4 = conv_mac_4 - 4'd7;
logic [31:0] bias_add_5;
assign bias_add_5 = conv_mac_5 + 7'd48;
logic [31:0] bias_add_6;
assign bias_add_6 = conv_mac_6 + 6'd25;
logic [31:0] bias_add_7;
assign bias_add_7 = conv_mac_7 + 5'd9;

logic [7:0] relu_0;
assign relu_0[7:0] = (bias_add_0[31]==0) ? ((bias_add_0<3'd6) ? {{bias_add_0[31],bias_add_0[10:4]}} :'d6) : '0;
logic [7:0] relu_1;
assign relu_1[7:0] = (bias_add_1[31]==0) ? ((bias_add_1<3'd6) ? {{bias_add_1[31],bias_add_1[10:4]}} :'d6) : '0;
logic [7:0] relu_2;
assign relu_2[7:0] = (bias_add_2[31]==0) ? ((bias_add_2<3'd6) ? {{bias_add_2[31],bias_add_2[10:4]}} :'d6) : '0;
logic [7:0] relu_3;
assign relu_3[7:0] = (bias_add_3[31]==0) ? ((bias_add_3<3'd6) ? {{bias_add_3[31],bias_add_3[10:4]}} :'d6) : '0;
logic [7:0] relu_4;
assign relu_4[7:0] = (bias_add_4[31]==0) ? ((bias_add_4<3'd6) ? {{bias_add_4[31],bias_add_4[10:4]}} :'d6) : '0;
logic [7:0] relu_5;
assign relu_5[7:0] = (bias_add_5[31]==0) ? ((bias_add_5<3'd6) ? {{bias_add_5[31],bias_add_5[10:4]}} :'d6) : '0;
logic [7:0] relu_6;
assign relu_6[7:0] = (bias_add_6[31]==0) ? ((bias_add_6<3'd6) ? {{bias_add_6[31],bias_add_6[10:4]}} :'d6) : '0;
logic [7:0] relu_7;
assign relu_7[7:0] = (bias_add_7[31]==0) ? ((bias_add_7<3'd6) ? {{bias_add_7[31],bias_add_7[10:4]}} :'d6) : '0;

assign output_act = {
	relu_7,
	relu_6,
	relu_5,
	relu_4,
	relu_3,
	relu_2,
	relu_1,
	relu_0
};

endmodule
module conv2_pw (
    input logic clk,
    input logic rstn,
    input logic valid,
    input logic [64-1:0] input_act,
    output logic [128-1:0] output_act,
    output logic ready
);
logic we;
logic [8:0] zero_number; 
assign zero_number = 9'd0; 
//1
logic [64-1:0] input_act_ff ;
always_ff @(posedge clk) begin
    if (rstn == 0) begin
        input_act_ff <= '0;
      //  ready <= '0;
    end
    else begin
        input_act_ff <= input_act;
     //   ready <= valid;
    end
end
logic [7:0] input_fmap_0;
assign input_fmap_0 = input_act_ff[7:0];
logic [7:0] input_fmap_1;
assign input_fmap_1 = input_act_ff[15:8];
logic [7:0] input_fmap_2;
assign input_fmap_2 = input_act_ff[23:16];
logic [7:0] input_fmap_3;
assign input_fmap_3 = input_act_ff[31:24];
logic [7:0] input_fmap_4;
assign input_fmap_4 = input_act_ff[39:32];
logic [7:0] input_fmap_5;
assign input_fmap_5 = input_act_ff[47:40];
logic [7:0] input_fmap_6;
assign input_fmap_6 = input_act_ff[55:48];
logic [7:0] input_fmap_7;
assign input_fmap_7 = input_act_ff[63:56];

logic [12-1:0] O0_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv2_pw_O0_I0_R0_C06_rom_inst (.q(O0_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O0_I0_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O0_I0_R0_C06_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv2_pw_O0_I0_R0_C06_rom_inst (.q(O0_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [11-1:0] O0_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_pw_O0_I1_R0_C02_rom_inst (.q(O0_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I1_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O0_I1_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O0_I1_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_pw_O0_I1_R0_C02_rom_inst (.q(O0_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [13-1:0] O0_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_pw_O0_I2_R0_C08_rom_inst (.q(O0_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I2_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O0_I2_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O0_I2_R0_C08_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_pw_O0_I2_R0_C08_rom_inst (.q(O0_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [12-1:0] O0_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv2_pw_O0_I3_R0_C06_rom_inst (.q(O0_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I3_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O0_I3_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O0_I3_R0_C06_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv2_pw_O0_I3_R0_C06_rom_inst (.q(O0_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [13-1:0] O0_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_pw_O0_I4_R0_C010_rom_inst (.q(O0_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I4_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O0_I4_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O0_I4_R0_C010_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_pw_O0_I4_R0_C010_rom_inst (.q(O0_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [11-1:0] O0_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_pw_O0_I5_R0_C02_rom_inst (.q(O0_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I5_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O0_I5_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O0_I5_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_pw_O0_I5_R0_C02_rom_inst (.q(O0_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [13-1:0] O0_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_pw_O0_I6_R0_C014_rom_inst (.q(O0_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I6_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O0_I6_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O0_I6_R0_C014_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_pw_O0_I6_R0_C014_rom_inst (.q(O0_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [10-1:0] O1_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv2_pw_O1_I0_R0_C01_rom_inst (.q(O1_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I0_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O1_I0_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O1_I0_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv2_pw_O1_I0_R0_C01_rom_inst (.q(O1_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [11-1:0] O1_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_pw_O1_I1_R0_C02_rom_inst (.q(O1_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O1_I1_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O1_I1_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_pw_O1_I1_R0_C02_rom_inst (.q(O1_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [11-1:0] O1_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_pw_O1_I2_R0_C03_rom_inst (.q(O1_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I2_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O1_I2_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O1_I2_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_pw_O1_I2_R0_C03_rom_inst (.q(O1_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [12-1:0] O1_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv2_pw_O1_I3_R0_C04_rom_inst (.q(O1_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I3_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O1_I3_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O1_I3_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv2_pw_O1_I3_R0_C04_rom_inst (.q(O1_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [10-1:0] O1_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv2_pw_O1_I5_R0_C01_rom_inst (.q(O1_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I5_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O1_I5_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O1_I5_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv2_pw_O1_I5_R0_C01_rom_inst (.q(O1_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [11-1:0] O1_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_pw_O1_I7_R0_C03_rom_inst (.q(O1_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I7_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O1_I7_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O1_I7_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_pw_O1_I7_R0_C03_rom_inst (.q(O1_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [10-1:0] O2_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv2_pw_O2_I0_R0_C01_rom_inst (.q(O2_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O2_I0_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O2_I0_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O2_I0_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv2_pw_O2_I0_R0_C01_rom_inst (.q(O2_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [13-1:0] O2_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_pw_O2_I1_R0_C013_rom_inst (.q(O2_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O2_I1_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O2_I1_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O2_I1_R0_C013_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_pw_O2_I1_R0_C013_rom_inst (.q(O2_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [11-1:0] O2_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_pw_O2_I3_R0_C03_rom_inst (.q(O2_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O2_I3_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O2_I3_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O2_I3_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_pw_O2_I3_R0_C03_rom_inst (.q(O2_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [11-1:0] O2_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_pw_O2_I5_R0_C02_rom_inst (.q(O2_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O2_I5_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O2_I5_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O2_I5_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_pw_O2_I5_R0_C02_rom_inst (.q(O2_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [10-1:0] O2_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv2_pw_O2_I7_R0_C01_rom_inst (.q(O2_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O2_I7_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O2_I7_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O2_I7_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv2_pw_O2_I7_R0_C01_rom_inst (.q(O2_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [10-1:0] O3_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv2_pw_O3_I1_R0_C01_rom_inst (.q(O3_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I1_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O3_I1_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O3_I1_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv2_pw_O3_I1_R0_C01_rom_inst (.q(O3_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [11-1:0] O3_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_pw_O3_I3_R0_C03_rom_inst (.q(O3_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O3_I3_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O3_I3_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_pw_O3_I3_R0_C03_rom_inst (.q(O3_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [10-1:0] O3_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv2_pw_O3_I5_R0_C01_rom_inst (.q(O3_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I5_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O3_I5_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O3_I5_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv2_pw_O3_I5_R0_C01_rom_inst (.q(O3_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [11-1:0] O3_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_pw_O3_I6_R0_C02_rom_inst (.q(O3_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I6_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O3_I6_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O3_I6_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_pw_O3_I6_R0_C02_rom_inst (.q(O3_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [11-1:0] O4_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_pw_O4_I0_R0_C02_rom_inst (.q(O4_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I0_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O4_I0_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O4_I0_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_pw_O4_I0_R0_C02_rom_inst (.q(O4_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [10-1:0] O4_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv2_pw_O4_I1_R0_C01_rom_inst (.q(O4_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I1_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I1_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O4_I1_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv2_pw_O4_I1_R0_C01_rom_inst (.q(O4_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [12-1:0] O4_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv2_pw_O4_I2_R0_C04_rom_inst (.q(O4_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I2_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O4_I2_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O4_I2_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv2_pw_O4_I2_R0_C04_rom_inst (.q(O4_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [11-1:0] O4_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_pw_O4_I3_R0_C02_rom_inst (.q(O4_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I3_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O4_I3_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O4_I3_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_pw_O4_I3_R0_C02_rom_inst (.q(O4_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [11-1:0] O4_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_pw_O4_I4_R0_C02_rom_inst (.q(O4_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O4_I4_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O4_I4_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_pw_O4_I4_R0_C02_rom_inst (.q(O4_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [10-1:0] O4_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv2_pw_O4_I5_R0_C01_rom_inst (.q(O4_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I5_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I5_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O4_I5_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv2_pw_O4_I5_R0_C01_rom_inst (.q(O4_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [12-1:0] O4_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv2_pw_O4_I6_R0_C04_rom_inst (.q(O4_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I6_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O4_I6_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O4_I6_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv2_pw_O4_I6_R0_C04_rom_inst (.q(O4_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [11-1:0] O4_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_pw_O4_I7_R0_C02_rom_inst (.q(O4_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I7_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O4_I7_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O4_I7_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_pw_O4_I7_R0_C02_rom_inst (.q(O4_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [13-1:0] O5_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_pw_O5_I0_R0_C09_rom_inst (.q(O5_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I0_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O5_I0_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O5_I0_R0_C09_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_pw_O5_I0_R0_C09_rom_inst (.q(O5_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [11-1:0] O5_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_pw_O5_I2_R0_C02_rom_inst (.q(O5_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I2_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O5_I2_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O5_I2_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_pw_O5_I2_R0_C02_rom_inst (.q(O5_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [10-1:0] O5_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv2_pw_O5_I3_R0_C01_rom_inst (.q(O5_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I3_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I3_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O5_I3_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv2_pw_O5_I3_R0_C01_rom_inst (.q(O5_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [10-1:0] O5_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv2_pw_O5_I4_R0_C01_rom_inst (.q(O5_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I4_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I4_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O5_I4_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv2_pw_O5_I4_R0_C01_rom_inst (.q(O5_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [12-1:0] O5_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv2_pw_O5_I5_R0_C04_rom_inst (.q(O5_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O5_I5_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O5_I5_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv2_pw_O5_I5_R0_C04_rom_inst (.q(O5_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [13-1:0] O5_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_pw_O5_I6_R0_C013_rom_inst (.q(O5_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I6_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O5_I6_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O5_I6_R0_C013_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_pw_O5_I6_R0_C013_rom_inst (.q(O5_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [10-1:0] O6_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv2_pw_O6_I2_R0_C01_rom_inst (.q(O6_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O6_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O6_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv2_pw_O6_I2_R0_C01_rom_inst (.q(O6_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [10-1:0] O6_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv2_pw_O6_I3_R0_C01_rom_inst (.q(O6_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I3_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O6_I3_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O6_I3_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv2_pw_O6_I3_R0_C01_rom_inst (.q(O6_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [11-1:0] O6_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_pw_O6_I4_R0_C03_rom_inst (.q(O6_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I4_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O6_I4_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O6_I4_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_pw_O6_I4_R0_C03_rom_inst (.q(O6_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [10-1:0] O6_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv2_pw_O6_I5_R0_C01_rom_inst (.q(O6_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I5_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O6_I5_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O6_I5_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv2_pw_O6_I5_R0_C01_rom_inst (.q(O6_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [10-1:0] O6_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv2_pw_O6_I6_R0_C01_rom_inst (.q(O6_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O6_I6_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O6_I6_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv2_pw_O6_I6_R0_C01_rom_inst (.q(O6_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [11-1:0] O6_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_pw_O6_I7_R0_C03_rom_inst (.q(O6_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I7_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O6_I7_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O6_I7_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_pw_O6_I7_R0_C03_rom_inst (.q(O6_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [11-1:0] O7_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_pw_O7_I0_R0_C02_rom_inst (.q(O7_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I0_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O7_I0_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O7_I0_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_pw_O7_I0_R0_C02_rom_inst (.q(O7_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [11-1:0] O7_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_pw_O7_I1_R0_C02_rom_inst (.q(O7_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I1_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O7_I1_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O7_I1_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_pw_O7_I1_R0_C02_rom_inst (.q(O7_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [13-1:0] O7_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_pw_O7_I3_R0_C013_rom_inst (.q(O7_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I3_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O7_I3_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O7_I3_R0_C013_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_pw_O7_I3_R0_C013_rom_inst (.q(O7_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [11-1:0] O7_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_pw_O7_I4_R0_C03_rom_inst (.q(O7_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I4_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O7_I4_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O7_I4_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_pw_O7_I4_R0_C03_rom_inst (.q(O7_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [12-1:0] O7_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv2_pw_O7_I5_R0_C06_rom_inst (.q(O7_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I5_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O7_I5_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O7_I5_R0_C06_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv2_pw_O7_I5_R0_C06_rom_inst (.q(O7_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [11-1:0] O7_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_pw_O7_I6_R0_C03_rom_inst (.q(O7_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I6_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O7_I6_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O7_I6_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_pw_O7_I6_R0_C03_rom_inst (.q(O7_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [13-1:0] O8_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_pw_O8_I1_R0_C09_rom_inst (.q(O8_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O8_I1_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O8_I1_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O8_I1_R0_C09_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_pw_O8_I1_R0_C09_rom_inst (.q(O8_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [10-1:0] O9_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv2_pw_O9_I0_R0_C01_rom_inst (.q(O9_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O9_I0_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O9_I0_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O9_I0_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv2_pw_O9_I0_R0_C01_rom_inst (.q(O9_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [11-1:0] O9_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_pw_O9_I2_R0_C02_rom_inst (.q(O9_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O9_I2_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O9_I2_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O9_I2_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_pw_O9_I2_R0_C02_rom_inst (.q(O9_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [11-1:0] O9_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_pw_O9_I3_R0_C02_rom_inst (.q(O9_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O9_I3_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O9_I3_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O9_I3_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_pw_O9_I3_R0_C02_rom_inst (.q(O9_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [11-1:0] O9_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_pw_O9_I4_R0_C03_rom_inst (.q(O9_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O9_I4_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O9_I4_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O9_I4_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_pw_O9_I4_R0_C03_rom_inst (.q(O9_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [10-1:0] O9_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv2_pw_O9_I5_R0_C01_rom_inst (.q(O9_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O9_I5_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O9_I5_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O9_I5_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv2_pw_O9_I5_R0_C01_rom_inst (.q(O9_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [10-1:0] O9_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv2_pw_O9_I6_R0_C01_rom_inst (.q(O9_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O9_I6_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O9_I6_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O9_I6_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv2_pw_O9_I6_R0_C01_rom_inst (.q(O9_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [13-1:0] O9_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_pw_O9_I7_R0_C010_rom_inst (.q(O9_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O9_I7_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O9_I7_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O9_I7_R0_C010_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_pw_O9_I7_R0_C010_rom_inst (.q(O9_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [13-1:0] O10_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_pw_O10_I0_R0_C08_rom_inst (.q(O10_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O10_I0_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O10_I0_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O10_I0_R0_C08_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_pw_O10_I0_R0_C08_rom_inst (.q(O10_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [11-1:0] O10_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_pw_O10_I5_R0_C02_rom_inst (.q(O10_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O10_I5_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O10_I5_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O10_I5_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_pw_O10_I5_R0_C02_rom_inst (.q(O10_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [11-1:0] O10_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_pw_O10_I6_R0_C03_rom_inst (.q(O10_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O10_I6_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O10_I6_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O10_I6_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_pw_O10_I6_R0_C03_rom_inst (.q(O10_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [10-1:0] O11_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv2_pw_O11_I0_R0_C01_rom_inst (.q(O11_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I0_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O11_I0_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O11_I0_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv2_pw_O11_I0_R0_C01_rom_inst (.q(O11_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [13-1:0] O11_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_pw_O11_I1_R0_C011_rom_inst (.q(O11_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I1_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O11_I1_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O11_I1_R0_C011_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_pw_O11_I1_R0_C011_rom_inst (.q(O11_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [12-1:0] O11_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv2_pw_O11_I3_R0_C07_rom_inst (.q(O11_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I3_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O11_I3_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O11_I3_R0_C07_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv2_pw_O11_I3_R0_C07_rom_inst (.q(O11_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [11-1:0] O11_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_pw_O11_I4_R0_C02_rom_inst (.q(O11_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I4_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O11_I4_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O11_I4_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_pw_O11_I4_R0_C02_rom_inst (.q(O11_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [10-1:0] O11_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv2_pw_O11_I7_R0_C01_rom_inst (.q(O11_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I7_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O11_I7_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O11_I7_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv2_pw_O11_I7_R0_C01_rom_inst (.q(O11_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [11-1:0] O12_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_pw_O12_I0_R0_C02_rom_inst (.q(O12_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I0_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O12_I0_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O12_I0_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_pw_O12_I0_R0_C02_rom_inst (.q(O12_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [12-1:0] O12_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv2_pw_O12_I1_R0_C04_rom_inst (.q(O12_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I1_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O12_I1_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O12_I1_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv2_pw_O12_I1_R0_C04_rom_inst (.q(O12_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [13-1:0] O12_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_pw_O12_I3_R0_C09_rom_inst (.q(O12_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I3_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O12_I3_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O12_I3_R0_C09_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_pw_O12_I3_R0_C09_rom_inst (.q(O12_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [11-1:0] O12_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_pw_O12_I4_R0_C03_rom_inst (.q(O12_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I4_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O12_I4_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O12_I4_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_pw_O12_I4_R0_C03_rom_inst (.q(O12_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [11-1:0] O12_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_pw_O12_I5_R0_C02_rom_inst (.q(O12_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I5_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O12_I5_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O12_I5_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_pw_O12_I5_R0_C02_rom_inst (.q(O12_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [10-1:0] O12_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv2_pw_O12_I6_R0_C01_rom_inst (.q(O12_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I6_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O12_I6_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O12_I6_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv2_pw_O12_I6_R0_C01_rom_inst (.q(O12_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [10-1:0] O12_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv2_pw_O12_I7_R0_C01_rom_inst (.q(O12_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I7_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O12_I7_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O12_I7_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv2_pw_O12_I7_R0_C01_rom_inst (.q(O12_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [10-1:0] O13_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv2_pw_O13_I0_R0_C01_rom_inst (.q(O13_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O13_I0_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O13_I0_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O13_I0_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv2_pw_O13_I0_R0_C01_rom_inst (.q(O13_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [11-1:0] O13_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_pw_O13_I1_R0_C03_rom_inst (.q(O13_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O13_I1_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O13_I1_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O13_I1_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_pw_O13_I1_R0_C03_rom_inst (.q(O13_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [10-1:0] O13_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv2_pw_O13_I2_R0_C01_rom_inst (.q(O13_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O13_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O13_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O13_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv2_pw_O13_I2_R0_C01_rom_inst (.q(O13_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [13-1:0] O13_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_pw_O13_I3_R0_C010_rom_inst (.q(O13_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O13_I3_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O13_I3_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O13_I3_R0_C010_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_pw_O13_I3_R0_C010_rom_inst (.q(O13_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [10-1:0] O13_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv2_pw_O13_I4_R0_C01_rom_inst (.q(O13_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O13_I4_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O13_I4_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O13_I4_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv2_pw_O13_I4_R0_C01_rom_inst (.q(O13_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [12-1:0] O13_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv2_pw_O13_I5_R0_C04_rom_inst (.q(O13_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O13_I5_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O13_I5_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O13_I5_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv2_pw_O13_I5_R0_C04_rom_inst (.q(O13_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [12-1:0] O13_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv2_pw_O13_I6_R0_C06_rom_inst (.q(O13_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O13_I6_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O13_I6_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O13_I6_R0_C06_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv2_pw_O13_I6_R0_C06_rom_inst (.q(O13_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [10-1:0] O14_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv2_pw_O14_I0_R0_C01_rom_inst (.q(O14_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I0_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O14_I0_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O14_I0_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv2_pw_O14_I0_R0_C01_rom_inst (.q(O14_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [10-1:0] O14_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv2_pw_O14_I1_R0_C01_rom_inst (.q(O14_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I1_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O14_I1_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O14_I1_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv2_pw_O14_I1_R0_C01_rom_inst (.q(O14_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [13-1:0] O14_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv2_pw_O14_I2_R0_C09_rom_inst (.q(O14_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I2_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O14_I2_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O14_I2_R0_C09_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv2_pw_O14_I2_R0_C09_rom_inst (.q(O14_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [11-1:0] O14_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_pw_O14_I3_R0_C03_rom_inst (.q(O14_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I3_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O14_I3_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O14_I3_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_pw_O14_I3_R0_C03_rom_inst (.q(O14_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [12-1:0] O14_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv2_pw_O14_I4_R0_C05_rom_inst (.q(O14_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I4_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O14_I4_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O14_I4_R0_C05_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv2_pw_O14_I4_R0_C05_rom_inst (.q(O14_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [11-1:0] O14_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_pw_O14_I5_R0_C02_rom_inst (.q(O14_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I5_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O14_I5_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O14_I5_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_pw_O14_I5_R0_C02_rom_inst (.q(O14_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [11-1:0] O14_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_pw_O14_I6_R0_C02_rom_inst (.q(O14_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I6_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O14_I6_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O14_I6_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_pw_O14_I6_R0_C02_rom_inst (.q(O14_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [10-1:0] O15_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv2_pw_O15_I0_R0_C01_rom_inst (.q(O15_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I0_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O15_I0_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O15_I0_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv2_pw_O15_I0_R0_C01_rom_inst (.q(O15_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [10-1:0] O15_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv2_pw_O15_I1_R0_C01_rom_inst (.q(O15_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I1_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O15_I1_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O15_I1_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv2_pw_O15_I1_R0_C01_rom_inst (.q(O15_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [12-1:0] O15_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv2_pw_O15_I2_R0_C05_rom_inst (.q(O15_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I2_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O15_I2_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O15_I2_R0_C05_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv2_pw_O15_I2_R0_C05_rom_inst (.q(O15_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [11-1:0] O15_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv2_pw_O15_I3_R0_C02_rom_inst (.q(O15_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I3_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O15_I3_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O15_I3_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv2_pw_O15_I3_R0_C02_rom_inst (.q(O15_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [12-1:0] O15_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv2_pw_O15_I4_R0_C05_rom_inst (.q(O15_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I4_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O15_I4_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O15_I4_R0_C05_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv2_pw_O15_I4_R0_C05_rom_inst (.q(O15_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [10-1:0] O15_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv2_pw_O15_I6_R0_C01_rom_inst (.q(O15_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I6_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O15_I6_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O15_I6_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv2_pw_O15_I6_R0_C01_rom_inst (.q(O15_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [12-1:0] O15_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv2_pw_O15_I7_R0_C04_rom_inst (.q(O15_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I7_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O15_I7_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv2_pw_O15_I7_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv2_pw_O15_I7_R0_C04_rom_inst (.q(O15_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic signed [31:0] conv_mac_0;
logic signed [31:0] O0_N0_S0;		always @(posedge clk) O0_N0_S0 <=     O0_I0_R0_C0_SM1   +  O0_I1_R0_C0_SM1  ;
 logic signed [31:0] O0_N2_S0;		always @(posedge clk) O0_N2_S0 <=     O0_I2_R0_C0_SM1   +  O0_I3_R0_C0_SM1  ;
 logic signed [31:0] O0_N4_S0;		always @(posedge clk) O0_N4_S0 <=     O0_I4_R0_C0_SM1   +  O0_I5_R0_C0_SM1  ;
 logic signed [31:0] O0_N6_S0;		always @(posedge clk) O0_N6_S0 <=     O0_I6_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O0_N0_S1;		always @(posedge clk) O0_N0_S1 <=     O0_N0_S0  +  O0_N2_S0 ;
 logic signed [31:0] O0_N2_S1;		always @(posedge clk) O0_N2_S1 <=     O0_N4_S0  +  O0_N6_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O0_N0_S2;		always @(posedge clk) O0_N0_S2 <=     O0_N0_S1  +  O0_N2_S1 ;
 assign conv_mac_0 = O0_N0_S2;

logic signed [31:0] conv_mac_1;
logic signed [31:0] O1_N0_S0;		always @(posedge clk) O1_N0_S0 <=     O1_I0_R0_C0_SM1   +  O1_I1_R0_C0_SM1  ;
 logic signed [31:0] O1_N2_S0;		always @(posedge clk) O1_N2_S0 <=     O1_I2_R0_C0_SM1   +  O1_I3_R0_C0_SM1  ;
 logic signed [31:0] O1_N4_S0;		always @(posedge clk) O1_N4_S0 <=     O1_I5_R0_C0_SM1   +  O1_I7_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O1_N0_S1;		always @(posedge clk) O1_N0_S1 <=     O1_N0_S0  +  O1_N2_S0 ;
 logic signed [31:0] O1_N2_S1;		always @(posedge clk) O1_N2_S1 <=     O1_N4_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O1_N0_S2;		always @(posedge clk) O1_N0_S2 <=     O1_N0_S1  +  O1_N2_S1 ;
 assign conv_mac_1 = O1_N0_S2;

logic signed [31:0] conv_mac_2;
logic signed [31:0] O2_N0_S0;		always @(posedge clk) O2_N0_S0 <=     O2_I0_R0_C0_SM1   +  O2_I1_R0_C0_SM1  ;
 logic signed [31:0] O2_N2_S0;		always @(posedge clk) O2_N2_S0 <=     O2_I3_R0_C0_SM1   +  O2_I5_R0_C0_SM1  ;
 logic signed [31:0] O2_N4_S0;		always @(posedge clk) O2_N4_S0 <=     O2_I7_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O2_N0_S1;		always @(posedge clk) O2_N0_S1 <=     O2_N0_S0  +  O2_N2_S0 ;
 logic signed [31:0] O2_N2_S1;		always @(posedge clk) O2_N2_S1 <=     O2_N4_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O2_N0_S2;		always @(posedge clk) O2_N0_S2 <=     O2_N0_S1  +  O2_N2_S1 ;
 assign conv_mac_2 = O2_N0_S2;

logic signed [31:0] conv_mac_3;
logic signed [31:0] O3_N0_S0;		always @(posedge clk) O3_N0_S0 <=     O3_I1_R0_C0_SM1   +  O3_I3_R0_C0_SM1  ;
 logic signed [31:0] O3_N2_S0;		always @(posedge clk) O3_N2_S0 <=     O3_I5_R0_C0_SM1   +  O3_I6_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O3_N0_S1;		always @(posedge clk) O3_N0_S1 <=     O3_N0_S0  +  O3_N2_S0 ;
 assign conv_mac_3 = O3_N0_S1;

logic signed [31:0] conv_mac_4;
logic signed [31:0] O4_N0_S0;		always @(posedge clk) O4_N0_S0 <=     O4_I0_R0_C0_SM1   +  O4_I1_R0_C0_SM1  ;
 logic signed [31:0] O4_N2_S0;		always @(posedge clk) O4_N2_S0 <=     O4_I2_R0_C0_SM1   +  O4_I3_R0_C0_SM1  ;
 logic signed [31:0] O4_N4_S0;		always @(posedge clk) O4_N4_S0 <=     O4_I4_R0_C0_SM1   +  O4_I5_R0_C0_SM1  ;
 logic signed [31:0] O4_N6_S0;		always @(posedge clk) O4_N6_S0 <=     O4_I6_R0_C0_SM1   +  O4_I7_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O4_N0_S1;		always @(posedge clk) O4_N0_S1 <=     O4_N0_S0  +  O4_N2_S0 ;
 logic signed [31:0] O4_N2_S1;		always @(posedge clk) O4_N2_S1 <=     O4_N4_S0  +  O4_N6_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O4_N0_S2;		always @(posedge clk) O4_N0_S2 <=     O4_N0_S1  +  O4_N2_S1 ;
 assign conv_mac_4 = O4_N0_S2;

logic signed [31:0] conv_mac_5;
logic signed [31:0] O5_N0_S0;		always @(posedge clk) O5_N0_S0 <=     O5_I0_R0_C0_SM1   +  O5_I2_R0_C0_SM1  ;
 logic signed [31:0] O5_N2_S0;		always @(posedge clk) O5_N2_S0 <=     O5_I3_R0_C0_SM1   +  O5_I4_R0_C0_SM1  ;
 logic signed [31:0] O5_N4_S0;		always @(posedge clk) O5_N4_S0 <=     O5_I5_R0_C0_SM1   +  O5_I6_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O5_N0_S1;		always @(posedge clk) O5_N0_S1 <=     O5_N0_S0  +  O5_N2_S0 ;
 logic signed [31:0] O5_N2_S1;		always @(posedge clk) O5_N2_S1 <=     O5_N4_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O5_N0_S2;		always @(posedge clk) O5_N0_S2 <=     O5_N0_S1  +  O5_N2_S1 ;
 assign conv_mac_5 = O5_N0_S2;

logic signed [31:0] conv_mac_6;
logic signed [31:0] O6_N0_S0;		always @(posedge clk) O6_N0_S0 <=     O6_I2_R0_C0_SM1   +  O6_I3_R0_C0_SM1  ;
 logic signed [31:0] O6_N2_S0;		always @(posedge clk) O6_N2_S0 <=     O6_I4_R0_C0_SM1   +  O6_I5_R0_C0_SM1  ;
 logic signed [31:0] O6_N4_S0;		always @(posedge clk) O6_N4_S0 <=     O6_I6_R0_C0_SM1   +  O6_I7_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O6_N0_S1;		always @(posedge clk) O6_N0_S1 <=     O6_N0_S0  +  O6_N2_S0 ;
 logic signed [31:0] O6_N2_S1;		always @(posedge clk) O6_N2_S1 <=     O6_N4_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O6_N0_S2;		always @(posedge clk) O6_N0_S2 <=     O6_N0_S1  +  O6_N2_S1 ;
 assign conv_mac_6 = O6_N0_S2;

logic signed [31:0] conv_mac_7;
logic signed [31:0] O7_N0_S0;		always @(posedge clk) O7_N0_S0 <=     O7_I0_R0_C0_SM1   +  O7_I1_R0_C0_SM1  ;
 logic signed [31:0] O7_N2_S0;		always @(posedge clk) O7_N2_S0 <=     O7_I3_R0_C0_SM1   +  O7_I4_R0_C0_SM1  ;
 logic signed [31:0] O7_N4_S0;		always @(posedge clk) O7_N4_S0 <=     O7_I5_R0_C0_SM1   +  O7_I6_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O7_N0_S1;		always @(posedge clk) O7_N0_S1 <=     O7_N0_S0  +  O7_N2_S0 ;
 logic signed [31:0] O7_N2_S1;		always @(posedge clk) O7_N2_S1 <=     O7_N4_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O7_N0_S2;		always @(posedge clk) O7_N0_S2 <=     O7_N0_S1  +  O7_N2_S1 ;
 assign conv_mac_7 = O7_N0_S2;

logic signed [31:0] conv_mac_8;
logic signed [31:0] O8_N0_S0;		always @(posedge clk) O8_N0_S0 <=     O8_I1_R0_C0_SM1      ;
 assign conv_mac_8 = O8_N0_S0;

logic signed [31:0] conv_mac_9;
logic signed [31:0] O9_N0_S0;		always @(posedge clk) O9_N0_S0 <=     O9_I0_R0_C0_SM1   +  O9_I2_R0_C0_SM1  ;
 logic signed [31:0] O9_N2_S0;		always @(posedge clk) O9_N2_S0 <=     O9_I3_R0_C0_SM1   +  O9_I4_R0_C0_SM1  ;
 logic signed [31:0] O9_N4_S0;		always @(posedge clk) O9_N4_S0 <=     O9_I5_R0_C0_SM1   +  O9_I6_R0_C0_SM1  ;
 logic signed [31:0] O9_N6_S0;		always @(posedge clk) O9_N6_S0 <=     O9_I7_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O9_N0_S1;		always @(posedge clk) O9_N0_S1 <=     O9_N0_S0  +  O9_N2_S0 ;
 logic signed [31:0] O9_N2_S1;		always @(posedge clk) O9_N2_S1 <=     O9_N4_S0  +  O9_N6_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O9_N0_S2;		always @(posedge clk) O9_N0_S2 <=     O9_N0_S1  +  O9_N2_S1 ;
 assign conv_mac_9 = O9_N0_S2;

logic signed [31:0] conv_mac_10;
logic signed [31:0] O10_N0_S0;		always @(posedge clk) O10_N0_S0 <=     O10_I0_R0_C0_SM1   +  O10_I5_R0_C0_SM1  ;
 logic signed [31:0] O10_N2_S0;		always @(posedge clk) O10_N2_S0 <=     O10_I6_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O10_N0_S1;		always @(posedge clk) O10_N0_S1 <=     O10_N0_S0  +  O10_N2_S0 ;
 assign conv_mac_10 = O10_N0_S1;

logic signed [31:0] conv_mac_11;
logic signed [31:0] O11_N0_S0;		always @(posedge clk) O11_N0_S0 <=     O11_I0_R0_C0_SM1   +  O11_I1_R0_C0_SM1  ;
 logic signed [31:0] O11_N2_S0;		always @(posedge clk) O11_N2_S0 <=     O11_I3_R0_C0_SM1   +  O11_I4_R0_C0_SM1  ;
 logic signed [31:0] O11_N4_S0;		always @(posedge clk) O11_N4_S0 <=     O11_I7_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O11_N0_S1;		always @(posedge clk) O11_N0_S1 <=     O11_N0_S0  +  O11_N2_S0 ;
 logic signed [31:0] O11_N2_S1;		always @(posedge clk) O11_N2_S1 <=     O11_N4_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O11_N0_S2;		always @(posedge clk) O11_N0_S2 <=     O11_N0_S1  +  O11_N2_S1 ;
 assign conv_mac_11 = O11_N0_S2;

logic signed [31:0] conv_mac_12;
logic signed [31:0] O12_N0_S0;		always @(posedge clk) O12_N0_S0 <=     O12_I0_R0_C0_SM1   +  O12_I1_R0_C0_SM1  ;
 logic signed [31:0] O12_N2_S0;		always @(posedge clk) O12_N2_S0 <=     O12_I3_R0_C0_SM1   +  O12_I4_R0_C0_SM1  ;
 logic signed [31:0] O12_N4_S0;		always @(posedge clk) O12_N4_S0 <=     O12_I5_R0_C0_SM1   +  O12_I6_R0_C0_SM1  ;
 logic signed [31:0] O12_N6_S0;		always @(posedge clk) O12_N6_S0 <=     O12_I7_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O12_N0_S1;		always @(posedge clk) O12_N0_S1 <=     O12_N0_S0  +  O12_N2_S0 ;
 logic signed [31:0] O12_N2_S1;		always @(posedge clk) O12_N2_S1 <=     O12_N4_S0  +  O12_N6_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O12_N0_S2;		always @(posedge clk) O12_N0_S2 <=     O12_N0_S1  +  O12_N2_S1 ;
 assign conv_mac_12 = O12_N0_S2;

logic signed [31:0] conv_mac_13;
logic signed [31:0] O13_N0_S0;		always @(posedge clk) O13_N0_S0 <=     O13_I0_R0_C0_SM1   +  O13_I1_R0_C0_SM1  ;
 logic signed [31:0] O13_N2_S0;		always @(posedge clk) O13_N2_S0 <=     O13_I2_R0_C0_SM1   +  O13_I3_R0_C0_SM1  ;
 logic signed [31:0] O13_N4_S0;		always @(posedge clk) O13_N4_S0 <=     O13_I4_R0_C0_SM1   +  O13_I5_R0_C0_SM1  ;
 logic signed [31:0] O13_N6_S0;		always @(posedge clk) O13_N6_S0 <=     O13_I6_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O13_N0_S1;		always @(posedge clk) O13_N0_S1 <=     O13_N0_S0  +  O13_N2_S0 ;
 logic signed [31:0] O13_N2_S1;		always @(posedge clk) O13_N2_S1 <=     O13_N4_S0  +  O13_N6_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O13_N0_S2;		always @(posedge clk) O13_N0_S2 <=     O13_N0_S1  +  O13_N2_S1 ;
 assign conv_mac_13 = O13_N0_S2;

logic signed [31:0] conv_mac_14;
logic signed [31:0] O14_N0_S0;		always @(posedge clk) O14_N0_S0 <=     O14_I0_R0_C0_SM1   +  O14_I1_R0_C0_SM1  ;
 logic signed [31:0] O14_N2_S0;		always @(posedge clk) O14_N2_S0 <=     O14_I2_R0_C0_SM1   +  O14_I3_R0_C0_SM1  ;
 logic signed [31:0] O14_N4_S0;		always @(posedge clk) O14_N4_S0 <=     O14_I4_R0_C0_SM1   +  O14_I5_R0_C0_SM1  ;
 logic signed [31:0] O14_N6_S0;		always @(posedge clk) O14_N6_S0 <=     O14_I6_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O14_N0_S1;		always @(posedge clk) O14_N0_S1 <=     O14_N0_S0  +  O14_N2_S0 ;
 logic signed [31:0] O14_N2_S1;		always @(posedge clk) O14_N2_S1 <=     O14_N4_S0  +  O14_N6_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O14_N0_S2;		always @(posedge clk) O14_N0_S2 <=     O14_N0_S1  +  O14_N2_S1 ;
 assign conv_mac_14 = O14_N0_S2;

logic signed [31:0] conv_mac_15;
logic signed [31:0] O15_N0_S0;		always @(posedge clk) O15_N0_S0 <=     O15_I0_R0_C0_SM1   +  O15_I1_R0_C0_SM1  ;
 logic signed [31:0] O15_N2_S0;		always @(posedge clk) O15_N2_S0 <=     O15_I2_R0_C0_SM1   +  O15_I3_R0_C0_SM1  ;
 logic signed [31:0] O15_N4_S0;		always @(posedge clk) O15_N4_S0 <=     O15_I4_R0_C0_SM1   +  O15_I6_R0_C0_SM1  ;
 logic signed [31:0] O15_N6_S0;		always @(posedge clk) O15_N6_S0 <=     O15_I7_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O15_N0_S1;		always @(posedge clk) O15_N0_S1 <=     O15_N0_S0  +  O15_N2_S0 ;
 logic signed [31:0] O15_N2_S1;		always @(posedge clk) O15_N2_S1 <=     O15_N4_S0  +  O15_N6_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O15_N0_S2;		always @(posedge clk) O15_N0_S2 <=     O15_N0_S1  +  O15_N2_S1 ;
 assign conv_mac_15 = O15_N0_S2;

logic valid_D1;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D1<= 0 ;
	else valid_D1<=valid;
end
logic valid_D2;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D2<= 0 ;
	else valid_D2<=valid_D1;
end
logic valid_D3;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D3<= 0 ;
	else valid_D3<=valid_D2;
end
logic valid_D4;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D4<= 0 ;
	else valid_D4<=valid_D3;
end
always_ff @(posedge clk) begin
	if (rstn == 0) ready <= 0 ;
	else ready <=valid_D4;
end
logic [31:0] bias_add_0;
assign bias_add_0 = conv_mac_0 - 6'd25;
logic [31:0] bias_add_1;
assign bias_add_1 = conv_mac_1 + 5'd13;
logic [31:0] bias_add_2;
assign bias_add_2 = conv_mac_2 - 3'd3;
logic [31:0] bias_add_3;
assign bias_add_3 = conv_mac_3 + 5'd10;
logic [31:0] bias_add_4;
assign bias_add_4 = conv_mac_4 + 7'd37;
logic [31:0] bias_add_5;
assign bias_add_5 = conv_mac_5 + 8'd75;
logic [31:0] bias_add_6;
assign bias_add_6 = conv_mac_6 + 6'd22;
logic [31:0] bias_add_7;
assign bias_add_7 = conv_mac_7 - 6'd18;
logic [31:0] bias_add_8;
assign bias_add_8 = conv_mac_8 + 4'd6;
logic [31:0] bias_add_9;
assign bias_add_9 = conv_mac_9 + 6'd17;
logic [31:0] bias_add_10;
assign bias_add_10 = conv_mac_10 + 4'd5;
logic [31:0] bias_add_11;
assign bias_add_11 = conv_mac_11 + 5'd10;
logic [31:0] bias_add_12;
assign bias_add_12 = conv_mac_12 - 5'd12;
logic [31:0] bias_add_13;
assign bias_add_13 = conv_mac_13 + 6'd26;
logic [31:0] bias_add_14;
assign bias_add_14 = conv_mac_14 - 3'd2;
logic [31:0] bias_add_15;
assign bias_add_15 = conv_mac_15 + 7'd33;

logic [7:0] relu_0;
assign relu_0[7:0] = (bias_add_0[31]==0) ? ((bias_add_0<3'd6) ? {{bias_add_0[31],bias_add_0[10:4]}} :'d6) : '0;
logic [7:0] relu_1;
assign relu_1[7:0] = (bias_add_1[31]==0) ? ((bias_add_1<3'd6) ? {{bias_add_1[31],bias_add_1[10:4]}} :'d6) : '0;
logic [7:0] relu_2;
assign relu_2[7:0] = (bias_add_2[31]==0) ? ((bias_add_2<3'd6) ? {{bias_add_2[31],bias_add_2[10:4]}} :'d6) : '0;
logic [7:0] relu_3;
assign relu_3[7:0] = (bias_add_3[31]==0) ? ((bias_add_3<3'd6) ? {{bias_add_3[31],bias_add_3[10:4]}} :'d6) : '0;
logic [7:0] relu_4;
assign relu_4[7:0] = (bias_add_4[31]==0) ? ((bias_add_4<3'd6) ? {{bias_add_4[31],bias_add_4[10:4]}} :'d6) : '0;
logic [7:0] relu_5;
assign relu_5[7:0] = (bias_add_5[31]==0) ? ((bias_add_5<3'd6) ? {{bias_add_5[31],bias_add_5[10:4]}} :'d6) : '0;
logic [7:0] relu_6;
assign relu_6[7:0] = (bias_add_6[31]==0) ? ((bias_add_6<3'd6) ? {{bias_add_6[31],bias_add_6[10:4]}} :'d6) : '0;
logic [7:0] relu_7;
assign relu_7[7:0] = (bias_add_7[31]==0) ? ((bias_add_7<3'd6) ? {{bias_add_7[31],bias_add_7[10:4]}} :'d6) : '0;
logic [7:0] relu_8;
assign relu_8[7:0] = (bias_add_8[31]==0) ? ((bias_add_8<3'd6) ? {{bias_add_8[31],bias_add_8[10:4]}} :'d6) : '0;
logic [7:0] relu_9;
assign relu_9[7:0] = (bias_add_9[31]==0) ? ((bias_add_9<3'd6) ? {{bias_add_9[31],bias_add_9[10:4]}} :'d6) : '0;
logic [7:0] relu_10;
assign relu_10[7:0] = (bias_add_10[31]==0) ? ((bias_add_10<3'd6) ? {{bias_add_10[31],bias_add_10[10:4]}} :'d6) : '0;
logic [7:0] relu_11;
assign relu_11[7:0] = (bias_add_11[31]==0) ? ((bias_add_11<3'd6) ? {{bias_add_11[31],bias_add_11[10:4]}} :'d6) : '0;
logic [7:0] relu_12;
assign relu_12[7:0] = (bias_add_12[31]==0) ? ((bias_add_12<3'd6) ? {{bias_add_12[31],bias_add_12[10:4]}} :'d6) : '0;
logic [7:0] relu_13;
assign relu_13[7:0] = (bias_add_13[31]==0) ? ((bias_add_13<3'd6) ? {{bias_add_13[31],bias_add_13[10:4]}} :'d6) : '0;
logic [7:0] relu_14;
assign relu_14[7:0] = (bias_add_14[31]==0) ? ((bias_add_14<3'd6) ? {{bias_add_14[31],bias_add_14[10:4]}} :'d6) : '0;
logic [7:0] relu_15;
assign relu_15[7:0] = (bias_add_15[31]==0) ? ((bias_add_15<3'd6) ? {{bias_add_15[31],bias_add_15[10:4]}} :'d6) : '0;

assign output_act = {
	relu_15,
	relu_14,
	relu_13,
	relu_12,
	relu_11,
	relu_10,
	relu_9,
	relu_8,
	relu_7,
	relu_6,
	relu_5,
	relu_4,
	relu_3,
	relu_2,
	relu_1,
	relu_0
};

endmodule
module conv3_pw (
    input logic clk,
    input logic rstn,
    input logic valid,
    input logic [128-1:0] input_act,
    output logic [128-1:0] output_act,
    output logic ready
);
logic we;
logic [8:0] zero_number; 
assign zero_number = 9'd0; 
//1
logic [128-1:0] input_act_ff ;
always_ff @(posedge clk) begin
    if (rstn == 0) begin
        input_act_ff <= '0;
      //  ready <= '0;
    end
    else begin
        input_act_ff <= input_act;
     //   ready <= valid;
    end
end
logic [7:0] input_fmap_0;
assign input_fmap_0 = input_act_ff[7:0];
logic [7:0] input_fmap_1;
assign input_fmap_1 = input_act_ff[15:8];
logic [7:0] input_fmap_2;
assign input_fmap_2 = input_act_ff[23:16];
logic [7:0] input_fmap_3;
assign input_fmap_3 = input_act_ff[31:24];
logic [7:0] input_fmap_4;
assign input_fmap_4 = input_act_ff[39:32];
logic [7:0] input_fmap_5;
assign input_fmap_5 = input_act_ff[47:40];
logic [7:0] input_fmap_6;
assign input_fmap_6 = input_act_ff[55:48];
logic [7:0] input_fmap_7;
assign input_fmap_7 = input_act_ff[63:56];
logic [7:0] input_fmap_8;
assign input_fmap_8 = input_act_ff[71:64];
logic [7:0] input_fmap_9;
assign input_fmap_9 = input_act_ff[79:72];
logic [7:0] input_fmap_10;
assign input_fmap_10 = input_act_ff[87:80];
logic [7:0] input_fmap_11;
assign input_fmap_11 = input_act_ff[95:88];
logic [7:0] input_fmap_12;
assign input_fmap_12 = input_act_ff[103:96];
logic [7:0] input_fmap_13;
assign input_fmap_13 = input_act_ff[111:104];
logic [7:0] input_fmap_14;
assign input_fmap_14 = input_act_ff[119:112];
logic [7:0] input_fmap_15;
assign input_fmap_15 = input_act_ff[127:120];

logic [10-1:0] O0_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O0_I2_R0_C01_rom_inst (.q(O0_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O0_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O0_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O0_I2_R0_C01_rom_inst (.q(O0_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [11-1:0] O0_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_pw_O0_I3_R0_C03_rom_inst (.q(O0_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I3_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O0_I3_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O0_I3_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_pw_O0_I3_R0_C03_rom_inst (.q(O0_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [10-1:0] O0_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O0_I4_R0_C01_rom_inst (.q(O0_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I4_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O0_I4_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O0_I4_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O0_I4_R0_C01_rom_inst (.q(O0_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [10-1:0] O0_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O0_I5_R0_C01_rom_inst (.q(O0_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I5_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O0_I5_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O0_I5_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O0_I5_R0_C01_rom_inst (.q(O0_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [10-1:0] O0_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O0_I8_R0_C01_rom_inst (.q(O0_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I8_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O0_I8_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O0_I8_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O0_I8_R0_C01_rom_inst (.q(O0_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [10-1:0] O0_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O0_I11_R0_C01_rom_inst (.q(O0_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I11_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O0_I11_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O0_I11_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O0_I11_R0_C01_rom_inst (.q(O0_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [10-1:0] O0_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O0_I12_R0_C01_rom_inst (.q(O0_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I12_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O0_I12_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O0_I12_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O0_I12_R0_C01_rom_inst (.q(O0_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [10-1:0] O0_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O0_I13_R0_C01_rom_inst (.q(O0_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I13_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O0_I13_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O0_I13_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O0_I13_R0_C01_rom_inst (.q(O0_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [10-1:0] O0_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O0_I15_R0_C01_rom_inst (.q(O0_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I15_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O0_I15_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O0_I15_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O0_I15_R0_C01_rom_inst (.q(O0_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [11-1:0] O1_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_pw_O1_I1_R0_C02_rom_inst (.q(O1_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O1_I1_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O1_I1_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_pw_O1_I1_R0_C02_rom_inst (.q(O1_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [11-1:0] O1_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_pw_O1_I2_R0_C02_rom_inst (.q(O1_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I2_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O1_I2_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O1_I2_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_pw_O1_I2_R0_C02_rom_inst (.q(O1_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [11-1:0] O1_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_pw_O1_I4_R0_C02_rom_inst (.q(O1_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I4_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O1_I4_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O1_I4_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_pw_O1_I4_R0_C02_rom_inst (.q(O1_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [10-1:0] O1_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O1_I5_R0_C01_rom_inst (.q(O1_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I5_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O1_I5_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O1_I5_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O1_I5_R0_C01_rom_inst (.q(O1_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [10-1:0] O1_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O1_I6_R0_C01_rom_inst (.q(O1_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I6_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O1_I6_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O1_I6_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O1_I6_R0_C01_rom_inst (.q(O1_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [10-1:0] O1_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O1_I7_R0_C01_rom_inst (.q(O1_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I7_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O1_I7_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O1_I7_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O1_I7_R0_C01_rom_inst (.q(O1_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [11-1:0] O1_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_pw_O1_I9_R0_C03_rom_inst (.q(O1_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I9_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O1_I9_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O1_I9_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_pw_O1_I9_R0_C03_rom_inst (.q(O1_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [10-1:0] O1_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O1_I11_R0_C01_rom_inst (.q(O1_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I11_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O1_I11_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O1_I11_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O1_I11_R0_C01_rom_inst (.q(O1_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [10-1:0] O1_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O1_I12_R0_C01_rom_inst (.q(O1_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I12_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O1_I12_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O1_I12_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O1_I12_R0_C01_rom_inst (.q(O1_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [10-1:0] O1_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O1_I13_R0_C01_rom_inst (.q(O1_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I13_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O1_I13_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O1_I13_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O1_I13_R0_C01_rom_inst (.q(O1_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [10-1:0] O1_I14_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O1_I14_R0_C01_rom_inst (.q(O1_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I14_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O1_I14_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O1_I14_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O1_I14_R0_C01_rom_inst (.q(O1_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clock  (clk));
logic [11-1:0] O1_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_pw_O1_I15_R0_C02_rom_inst (.q(O1_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I15_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O1_I15_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O1_I15_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_pw_O1_I15_R0_C02_rom_inst (.q(O1_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [10-1:0] O2_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O2_I0_R0_C01_rom_inst (.q(O2_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O2_I0_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O2_I0_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O2_I0_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O2_I0_R0_C01_rom_inst (.q(O2_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [10-1:0] O2_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O2_I1_R0_C01_rom_inst (.q(O2_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O2_I1_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O2_I1_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O2_I1_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O2_I1_R0_C01_rom_inst (.q(O2_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [11-1:0] O2_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_pw_O2_I2_R0_C02_rom_inst (.q(O2_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O2_I2_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O2_I2_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_pw_O2_I2_R0_C02_rom_inst (.q(O2_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [11-1:0] O2_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_pw_O2_I3_R0_C02_rom_inst (.q(O2_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O2_I3_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O2_I3_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O2_I3_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_pw_O2_I3_R0_C02_rom_inst (.q(O2_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [10-1:0] O2_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O2_I4_R0_C01_rom_inst (.q(O2_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O2_I4_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O2_I4_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O2_I4_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O2_I4_R0_C01_rom_inst (.q(O2_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [10-1:0] O2_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O2_I5_R0_C01_rom_inst (.q(O2_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O2_I5_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O2_I5_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O2_I5_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O2_I5_R0_C01_rom_inst (.q(O2_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [10-1:0] O2_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O2_I6_R0_C01_rom_inst (.q(O2_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O2_I6_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O2_I6_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O2_I6_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O2_I6_R0_C01_rom_inst (.q(O2_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [11-1:0] O2_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_pw_O2_I7_R0_C02_rom_inst (.q(O2_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O2_I7_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O2_I7_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O2_I7_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_pw_O2_I7_R0_C02_rom_inst (.q(O2_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [11-1:0] O2_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_pw_O2_I8_R0_C02_rom_inst (.q(O2_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O2_I8_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O2_I8_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O2_I8_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_pw_O2_I8_R0_C02_rom_inst (.q(O2_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [10-1:0] O2_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O2_I9_R0_C01_rom_inst (.q(O2_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O2_I9_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O2_I9_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O2_I9_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O2_I9_R0_C01_rom_inst (.q(O2_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [10-1:0] O2_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O2_I11_R0_C01_rom_inst (.q(O2_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O2_I11_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O2_I11_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O2_I11_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O2_I11_R0_C01_rom_inst (.q(O2_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [11-1:0] O2_I14_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_pw_O2_I14_R0_C03_rom_inst (.q(O2_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clk(clk),.d(0),.we(0));
//assign O2_I14_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O2_I14_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O2_I14_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_pw_O2_I14_R0_C03_rom_inst (.q(O2_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clock  (clk));
logic [12-1:0] O2_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_pw_O2_I15_R0_C04_rom_inst (.q(O2_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O2_I15_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O2_I15_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O2_I15_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_pw_O2_I15_R0_C04_rom_inst (.q(O2_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [10-1:0] O3_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O3_I1_R0_C01_rom_inst (.q(O3_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I1_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O3_I1_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O3_I1_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O3_I1_R0_C01_rom_inst (.q(O3_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [11-1:0] O3_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_pw_O3_I4_R0_C02_rom_inst (.q(O3_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I4_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O3_I4_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O3_I4_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_pw_O3_I4_R0_C02_rom_inst (.q(O3_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [10-1:0] O3_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O3_I5_R0_C01_rom_inst (.q(O3_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I5_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O3_I5_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O3_I5_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O3_I5_R0_C01_rom_inst (.q(O3_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [13-1:0] O3_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv3_pw_O3_I6_R0_C08_rom_inst (.q(O3_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I6_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O3_I6_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O3_I6_R0_C08_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv3_pw_O3_I6_R0_C08_rom_inst (.q(O3_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [10-1:0] O3_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O3_I9_R0_C01_rom_inst (.q(O3_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I9_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O3_I9_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O3_I9_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O3_I9_R0_C01_rom_inst (.q(O3_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [10-1:0] O3_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O3_I13_R0_C01_rom_inst (.q(O3_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I13_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O3_I13_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O3_I13_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O3_I13_R0_C01_rom_inst (.q(O3_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [10-1:0] O3_I14_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O3_I14_R0_C01_rom_inst (.q(O3_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I14_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O3_I14_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O3_I14_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O3_I14_R0_C01_rom_inst (.q(O3_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clock  (clk));
logic [11-1:0] O3_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_pw_O3_I15_R0_C02_rom_inst (.q(O3_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I15_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O3_I15_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O3_I15_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_pw_O3_I15_R0_C02_rom_inst (.q(O3_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [10-1:0] O4_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O4_I1_R0_C01_rom_inst (.q(O4_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I1_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I1_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O4_I1_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O4_I1_R0_C01_rom_inst (.q(O4_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [10-1:0] O4_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O4_I2_R0_C01_rom_inst (.q(O4_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O4_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O4_I2_R0_C01_rom_inst (.q(O4_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [10-1:0] O4_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O4_I3_R0_C01_rom_inst (.q(O4_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I3_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I3_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O4_I3_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O4_I3_R0_C01_rom_inst (.q(O4_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [10-1:0] O4_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O4_I5_R0_C01_rom_inst (.q(O4_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I5_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I5_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O4_I5_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O4_I5_R0_C01_rom_inst (.q(O4_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [10-1:0] O4_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O4_I6_R0_C01_rom_inst (.q(O4_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I6_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I6_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O4_I6_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O4_I6_R0_C01_rom_inst (.q(O4_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [12-1:0] O4_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_pw_O4_I9_R0_C04_rom_inst (.q(O4_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I9_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O4_I9_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O4_I9_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_pw_O4_I9_R0_C04_rom_inst (.q(O4_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [10-1:0] O4_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O4_I13_R0_C01_rom_inst (.q(O4_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I13_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I13_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O4_I13_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O4_I13_R0_C01_rom_inst (.q(O4_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [11-1:0] O4_I14_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_pw_O4_I14_R0_C02_rom_inst (.q(O4_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I14_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O4_I14_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O4_I14_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_pw_O4_I14_R0_C02_rom_inst (.q(O4_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clock  (clk));
logic [11-1:0] O4_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_pw_O4_I15_R0_C03_rom_inst (.q(O4_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I15_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O4_I15_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O4_I15_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_pw_O4_I15_R0_C03_rom_inst (.q(O4_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [10-1:0] O5_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O5_I0_R0_C01_rom_inst (.q(O5_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I0_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I0_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O5_I0_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O5_I0_R0_C01_rom_inst (.q(O5_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [10-1:0] O5_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O5_I3_R0_C01_rom_inst (.q(O5_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I3_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I3_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O5_I3_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O5_I3_R0_C01_rom_inst (.q(O5_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [10-1:0] O5_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O5_I4_R0_C01_rom_inst (.q(O5_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I4_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I4_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O5_I4_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O5_I4_R0_C01_rom_inst (.q(O5_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [10-1:0] O5_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O5_I5_R0_C01_rom_inst (.q(O5_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I5_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O5_I5_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O5_I5_R0_C01_rom_inst (.q(O5_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [11-1:0] O5_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_pw_O5_I7_R0_C02_rom_inst (.q(O5_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I7_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O5_I7_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O5_I7_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_pw_O5_I7_R0_C02_rom_inst (.q(O5_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [10-1:0] O5_I10_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O5_I10_R0_C01_rom_inst (.q(O5_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I10_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I10_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O5_I10_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O5_I10_R0_C01_rom_inst (.q(O5_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clock  (clk));
logic [12-1:0] O5_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_pw_O5_I13_R0_C04_rom_inst (.q(O5_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I13_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O5_I13_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O5_I13_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_pw_O5_I13_R0_C04_rom_inst (.q(O5_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [10-1:0] O5_I14_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O5_I14_R0_C01_rom_inst (.q(O5_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I14_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I14_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O5_I14_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O5_I14_R0_C01_rom_inst (.q(O5_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clock  (clk));
logic [10-1:0] O6_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O6_I0_R0_C01_rom_inst (.q(O6_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I0_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O6_I0_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O6_I0_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O6_I0_R0_C01_rom_inst (.q(O6_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [12-1:0] O6_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_pw_O6_I1_R0_C05_rom_inst (.q(O6_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I1_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O6_I1_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O6_I1_R0_C05_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_pw_O6_I1_R0_C05_rom_inst (.q(O6_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [12-1:0] O6_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_pw_O6_I2_R0_C05_rom_inst (.q(O6_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I2_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O6_I2_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O6_I2_R0_C05_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_pw_O6_I2_R0_C05_rom_inst (.q(O6_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [10-1:0] O6_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O6_I6_R0_C01_rom_inst (.q(O6_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O6_I6_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O6_I6_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O6_I6_R0_C01_rom_inst (.q(O6_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [10-1:0] O6_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O6_I8_R0_C01_rom_inst (.q(O6_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I8_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O6_I8_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O6_I8_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O6_I8_R0_C01_rom_inst (.q(O6_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [10-1:0] O6_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O6_I9_R0_C01_rom_inst (.q(O6_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I9_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O6_I9_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O6_I9_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O6_I9_R0_C01_rom_inst (.q(O6_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [11-1:0] O7_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_pw_O7_I0_R0_C03_rom_inst (.q(O7_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I0_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O7_I0_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O7_I0_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_pw_O7_I0_R0_C03_rom_inst (.q(O7_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [10-1:0] O7_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O7_I2_R0_C01_rom_inst (.q(O7_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O7_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O7_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O7_I2_R0_C01_rom_inst (.q(O7_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [12-1:0] O7_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_pw_O7_I3_R0_C04_rom_inst (.q(O7_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I3_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O7_I3_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O7_I3_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_pw_O7_I3_R0_C04_rom_inst (.q(O7_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [11-1:0] O7_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_pw_O7_I4_R0_C02_rom_inst (.q(O7_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I4_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O7_I4_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O7_I4_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_pw_O7_I4_R0_C02_rom_inst (.q(O7_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [13-1:0] O7_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv3_pw_O7_I5_R0_C010_rom_inst (.q(O7_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I5_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O7_I5_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O7_I5_R0_C010_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv3_pw_O7_I5_R0_C010_rom_inst (.q(O7_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [11-1:0] O7_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_pw_O7_I7_R0_C02_rom_inst (.q(O7_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O7_I7_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O7_I7_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_pw_O7_I7_R0_C02_rom_inst (.q(O7_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [13-1:0] O7_I10_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv3_pw_O7_I10_R0_C011_rom_inst (.q(O7_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I10_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O7_I10_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O7_I10_R0_C011_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv3_pw_O7_I10_R0_C011_rom_inst (.q(O7_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clock  (clk));
logic [11-1:0] O7_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_pw_O7_I13_R0_C02_rom_inst (.q(O7_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I13_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O7_I13_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O7_I13_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_pw_O7_I13_R0_C02_rom_inst (.q(O7_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [10-1:0] O7_I14_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O7_I14_R0_C01_rom_inst (.q(O7_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I14_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O7_I14_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O7_I14_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O7_I14_R0_C01_rom_inst (.q(O7_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clock  (clk));
logic [10-1:0] O8_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O8_I1_R0_C01_rom_inst (.q(O8_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O8_I1_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O8_I1_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O8_I1_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O8_I1_R0_C01_rom_inst (.q(O8_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [10-1:0] O8_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O8_I5_R0_C01_rom_inst (.q(O8_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O8_I5_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O8_I5_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O8_I5_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O8_I5_R0_C01_rom_inst (.q(O8_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [12-1:0] O8_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_pw_O8_I6_R0_C06_rom_inst (.q(O8_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O8_I6_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O8_I6_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O8_I6_R0_C06_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_pw_O8_I6_R0_C06_rom_inst (.q(O8_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [10-1:0] O8_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O8_I9_R0_C01_rom_inst (.q(O8_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O8_I9_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O8_I9_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O8_I9_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O8_I9_R0_C01_rom_inst (.q(O8_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [10-1:0] O8_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O8_I12_R0_C01_rom_inst (.q(O8_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O8_I12_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O8_I12_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O8_I12_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O8_I12_R0_C01_rom_inst (.q(O8_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [10-1:0] O8_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O8_I13_R0_C01_rom_inst (.q(O8_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O8_I13_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O8_I13_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O8_I13_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O8_I13_R0_C01_rom_inst (.q(O8_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [10-1:0] O8_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O8_I15_R0_C01_rom_inst (.q(O8_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O8_I15_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O8_I15_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O8_I15_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O8_I15_R0_C01_rom_inst (.q(O8_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [10-1:0] O9_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O9_I3_R0_C01_rom_inst (.q(O9_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O9_I3_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O9_I3_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O9_I3_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O9_I3_R0_C01_rom_inst (.q(O9_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [10-1:0] O9_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O9_I4_R0_C01_rom_inst (.q(O9_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O9_I4_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O9_I4_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O9_I4_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O9_I4_R0_C01_rom_inst (.q(O9_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [10-1:0] O9_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O9_I5_R0_C01_rom_inst (.q(O9_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O9_I5_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O9_I5_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O9_I5_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O9_I5_R0_C01_rom_inst (.q(O9_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [13-1:0] O9_I10_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv3_pw_O9_I10_R0_C08_rom_inst (.q(O9_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clk(clk),.d(0),.we(0));
//assign O9_I10_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O9_I10_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O9_I10_R0_C08_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv3_pw_O9_I10_R0_C08_rom_inst (.q(O9_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clock  (clk));
logic [10-1:0] O9_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O9_I13_R0_C01_rom_inst (.q(O9_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O9_I13_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O9_I13_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O9_I13_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O9_I13_R0_C01_rom_inst (.q(O9_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [11-1:0] O10_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_pw_O10_I3_R0_C02_rom_inst (.q(O10_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O10_I3_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O10_I3_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O10_I3_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_pw_O10_I3_R0_C02_rom_inst (.q(O10_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [12-1:0] O10_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_pw_O10_I5_R0_C07_rom_inst (.q(O10_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O10_I5_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O10_I5_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O10_I5_R0_C07_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_pw_O10_I5_R0_C07_rom_inst (.q(O10_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [11-1:0] O10_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_pw_O10_I6_R0_C02_rom_inst (.q(O10_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O10_I6_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O10_I6_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O10_I6_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_pw_O10_I6_R0_C02_rom_inst (.q(O10_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [10-1:0] O10_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O10_I7_R0_C01_rom_inst (.q(O10_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O10_I7_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O10_I7_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O10_I7_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O10_I7_R0_C01_rom_inst (.q(O10_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [13-1:0] O10_I10_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv3_pw_O10_I10_R0_C011_rom_inst (.q(O10_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clk(clk),.d(0),.we(0));
//assign O10_I10_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O10_I10_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O10_I10_R0_C011_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv3_pw_O10_I10_R0_C011_rom_inst (.q(O10_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clock  (clk));
logic [10-1:0] O10_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O10_I11_R0_C01_rom_inst (.q(O10_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O10_I11_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O10_I11_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O10_I11_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O10_I11_R0_C01_rom_inst (.q(O10_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [10-1:0] O10_I14_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O10_I14_R0_C01_rom_inst (.q(O10_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clk(clk),.d(0),.we(0));
//assign O10_I14_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O10_I14_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O10_I14_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O10_I14_R0_C01_rom_inst (.q(O10_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clock  (clk));
logic [11-1:0] O11_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_pw_O11_I1_R0_C02_rom_inst (.q(O11_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I1_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O11_I1_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O11_I1_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_pw_O11_I1_R0_C02_rom_inst (.q(O11_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [10-1:0] O11_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O11_I3_R0_C01_rom_inst (.q(O11_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I3_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O11_I3_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O11_I3_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O11_I3_R0_C01_rom_inst (.q(O11_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [10-1:0] O11_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O11_I4_R0_C01_rom_inst (.q(O11_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I4_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O11_I4_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O11_I4_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O11_I4_R0_C01_rom_inst (.q(O11_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [11-1:0] O11_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_pw_O11_I8_R0_C03_rom_inst (.q(O11_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I8_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O11_I8_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O11_I8_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_pw_O11_I8_R0_C03_rom_inst (.q(O11_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [10-1:0] O11_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O11_I9_R0_C01_rom_inst (.q(O11_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I9_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O11_I9_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O11_I9_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O11_I9_R0_C01_rom_inst (.q(O11_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [11-1:0] O11_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_pw_O11_I11_R0_C03_rom_inst (.q(O11_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I11_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O11_I11_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O11_I11_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_pw_O11_I11_R0_C03_rom_inst (.q(O11_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [11-1:0] O11_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_pw_O11_I12_R0_C02_rom_inst (.q(O11_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I12_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O11_I12_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O11_I12_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_pw_O11_I12_R0_C02_rom_inst (.q(O11_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [10-1:0] O11_I14_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O11_I14_R0_C01_rom_inst (.q(O11_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I14_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O11_I14_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O11_I14_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O11_I14_R0_C01_rom_inst (.q(O11_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clock  (clk));
logic [10-1:0] O12_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O12_I2_R0_C01_rom_inst (.q(O12_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O12_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O12_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O12_I2_R0_C01_rom_inst (.q(O12_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [13-1:0] O12_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv3_pw_O12_I3_R0_C011_rom_inst (.q(O12_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I3_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O12_I3_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O12_I3_R0_C011_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv3_pw_O12_I3_R0_C011_rom_inst (.q(O12_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [10-1:0] O12_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O12_I4_R0_C01_rom_inst (.q(O12_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I4_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O12_I4_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O12_I4_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O12_I4_R0_C01_rom_inst (.q(O12_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [12-1:0] O12_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_pw_O12_I5_R0_C07_rom_inst (.q(O12_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I5_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O12_I5_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O12_I5_R0_C07_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_pw_O12_I5_R0_C07_rom_inst (.q(O12_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [11-1:0] O12_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_pw_O12_I6_R0_C02_rom_inst (.q(O12_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I6_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O12_I6_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O12_I6_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_pw_O12_I6_R0_C02_rom_inst (.q(O12_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [10-1:0] O12_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O12_I7_R0_C01_rom_inst (.q(O12_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I7_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O12_I7_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O12_I7_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O12_I7_R0_C01_rom_inst (.q(O12_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [12-1:0] O12_I10_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_pw_O12_I10_R0_C04_rom_inst (.q(O12_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I10_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O12_I10_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O12_I10_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_pw_O12_I10_R0_C04_rom_inst (.q(O12_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clock  (clk));
logic [10-1:0] O12_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O12_I11_R0_C01_rom_inst (.q(O12_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I11_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O12_I11_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O12_I11_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O12_I11_R0_C01_rom_inst (.q(O12_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [10-1:0] O12_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O12_I12_R0_C01_rom_inst (.q(O12_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I12_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O12_I12_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O12_I12_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O12_I12_R0_C01_rom_inst (.q(O12_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [10-1:0] O12_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O12_I13_R0_C01_rom_inst (.q(O12_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I13_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O12_I13_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O12_I13_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O12_I13_R0_C01_rom_inst (.q(O12_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [10-1:0] O13_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O13_I1_R0_C01_rom_inst (.q(O13_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O13_I1_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O13_I1_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O13_I1_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O13_I1_R0_C01_rom_inst (.q(O13_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [10-1:0] O13_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O13_I2_R0_C01_rom_inst (.q(O13_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O13_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O13_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O13_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O13_I2_R0_C01_rom_inst (.q(O13_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [10-1:0] O13_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O13_I4_R0_C01_rom_inst (.q(O13_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O13_I4_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O13_I4_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O13_I4_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O13_I4_R0_C01_rom_inst (.q(O13_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [10-1:0] O13_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O13_I6_R0_C01_rom_inst (.q(O13_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O13_I6_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O13_I6_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O13_I6_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O13_I6_R0_C01_rom_inst (.q(O13_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [12-1:0] O13_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_pw_O13_I8_R0_C05_rom_inst (.q(O13_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O13_I8_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O13_I8_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O13_I8_R0_C05_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_pw_O13_I8_R0_C05_rom_inst (.q(O13_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [12-1:0] O13_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_pw_O13_I11_R0_C05_rom_inst (.q(O13_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O13_I11_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O13_I11_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O13_I11_R0_C05_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_pw_O13_I11_R0_C05_rom_inst (.q(O13_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [12-1:0] O13_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_pw_O13_I12_R0_C05_rom_inst (.q(O13_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O13_I12_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O13_I12_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O13_I12_R0_C05_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_pw_O13_I12_R0_C05_rom_inst (.q(O13_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [10-1:0] O14_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O14_I0_R0_C01_rom_inst (.q(O14_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I0_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O14_I0_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O14_I0_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O14_I0_R0_C01_rom_inst (.q(O14_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [10-1:0] O14_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O14_I1_R0_C01_rom_inst (.q(O14_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I1_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O14_I1_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O14_I1_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O14_I1_R0_C01_rom_inst (.q(O14_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [10-1:0] O14_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O14_I2_R0_C01_rom_inst (.q(O14_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O14_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O14_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O14_I2_R0_C01_rom_inst (.q(O14_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [10-1:0] O14_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O14_I3_R0_C01_rom_inst (.q(O14_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I3_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O14_I3_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O14_I3_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O14_I3_R0_C01_rom_inst (.q(O14_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [11-1:0] O14_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_pw_O14_I6_R0_C02_rom_inst (.q(O14_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I6_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O14_I6_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O14_I6_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_pw_O14_I6_R0_C02_rom_inst (.q(O14_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [10-1:0] O14_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O14_I7_R0_C01_rom_inst (.q(O14_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I7_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O14_I7_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O14_I7_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O14_I7_R0_C01_rom_inst (.q(O14_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [10-1:0] O14_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O14_I9_R0_C01_rom_inst (.q(O14_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I9_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O14_I9_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O14_I9_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O14_I9_R0_C01_rom_inst (.q(O14_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [10-1:0] O14_I14_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O14_I14_R0_C01_rom_inst (.q(O14_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I14_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O14_I14_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O14_I14_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O14_I14_R0_C01_rom_inst (.q(O14_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clock  (clk));
logic [10-1:0] O15_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O15_I0_R0_C01_rom_inst (.q(O15_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I0_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O15_I0_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O15_I0_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O15_I0_R0_C01_rom_inst (.q(O15_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [11-1:0] O15_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_pw_O15_I1_R0_C02_rom_inst (.q(O15_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I1_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O15_I1_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O15_I1_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_pw_O15_I1_R0_C02_rom_inst (.q(O15_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [10-1:0] O15_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O15_I2_R0_C01_rom_inst (.q(O15_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O15_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O15_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O15_I2_R0_C01_rom_inst (.q(O15_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [11-1:0] O15_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_pw_O15_I3_R0_C03_rom_inst (.q(O15_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I3_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O15_I3_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O15_I3_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_pw_O15_I3_R0_C03_rom_inst (.q(O15_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [10-1:0] O15_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O15_I4_R0_C01_rom_inst (.q(O15_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I4_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O15_I4_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O15_I4_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O15_I4_R0_C01_rom_inst (.q(O15_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [10-1:0] O15_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O15_I5_R0_C01_rom_inst (.q(O15_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I5_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O15_I5_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O15_I5_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O15_I5_R0_C01_rom_inst (.q(O15_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [10-1:0] O15_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O15_I6_R0_C01_rom_inst (.q(O15_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I6_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O15_I6_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O15_I6_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O15_I6_R0_C01_rom_inst (.q(O15_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [11-1:0] O15_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_pw_O15_I7_R0_C03_rom_inst (.q(O15_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I7_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O15_I7_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O15_I7_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_pw_O15_I7_R0_C03_rom_inst (.q(O15_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [10-1:0] O15_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O15_I8_R0_C01_rom_inst (.q(O15_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I8_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O15_I8_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O15_I8_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O15_I8_R0_C01_rom_inst (.q(O15_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [11-1:0] O15_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv3_pw_O15_I9_R0_C03_rom_inst (.q(O15_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I9_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O15_I9_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O15_I9_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv3_pw_O15_I9_R0_C03_rom_inst (.q(O15_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [10-1:0] O15_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O15_I11_R0_C01_rom_inst (.q(O15_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I11_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O15_I11_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O15_I11_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O15_I11_R0_C01_rom_inst (.q(O15_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [10-1:0] O15_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O15_I12_R0_C01_rom_inst (.q(O15_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I12_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O15_I12_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O15_I12_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O15_I12_R0_C01_rom_inst (.q(O15_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [10-1:0] O15_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv3_pw_O15_I13_R0_C01_rom_inst (.q(O15_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I13_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O15_I13_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O15_I13_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv3_pw_O15_I13_R0_C01_rom_inst (.q(O15_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [12-1:0] O15_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv3_pw_O15_I15_R0_C04_rom_inst (.q(O15_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I15_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O15_I15_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv3_pw_O15_I15_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv3_pw_O15_I15_R0_C04_rom_inst (.q(O15_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic signed [31:0] conv_mac_0;
logic signed [31:0] O0_N0_S0;		always @(posedge clk) O0_N0_S0 <=     O0_I2_R0_C0_SM1   +  O0_I3_R0_C0_SM1  ;
 logic signed [31:0] O0_N2_S0;		always @(posedge clk) O0_N2_S0 <=     O0_I4_R0_C0_SM1   +  O0_I5_R0_C0_SM1  ;
 logic signed [31:0] O0_N4_S0;		always @(posedge clk) O0_N4_S0 <=     O0_I8_R0_C0_SM1   +  O0_I11_R0_C0_SM1  ;
 logic signed [31:0] O0_N6_S0;		always @(posedge clk) O0_N6_S0 <=     O0_I12_R0_C0_SM1   +  O0_I13_R0_C0_SM1  ;
 logic signed [31:0] O0_N8_S0;		always @(posedge clk) O0_N8_S0 <=     O0_I15_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O0_N0_S1;		always @(posedge clk) O0_N0_S1 <=     O0_N0_S0  +  O0_N2_S0 ;
 logic signed [31:0] O0_N2_S1;		always @(posedge clk) O0_N2_S1 <=     O0_N4_S0  +  O0_N6_S0 ;
 logic signed [31:0] O0_N4_S1;		always @(posedge clk) O0_N4_S1 <=     O0_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O0_N0_S2;		always @(posedge clk) O0_N0_S2 <=     O0_N0_S1  +  O0_N2_S1 ;
 logic signed [31:0] O0_N2_S2;		always @(posedge clk) O0_N2_S2 <=     O0_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O0_N0_S3;		always @(posedge clk) O0_N0_S3 <=     O0_N0_S2  +  O0_N2_S2 ;
 assign conv_mac_0 = O0_N0_S3;

logic signed [31:0] conv_mac_1;
logic signed [31:0] O1_N0_S0;		always @(posedge clk) O1_N0_S0 <=     O1_I1_R0_C0_SM1   +  O1_I2_R0_C0_SM1  ;
 logic signed [31:0] O1_N2_S0;		always @(posedge clk) O1_N2_S0 <=     O1_I4_R0_C0_SM1   +  O1_I5_R0_C0_SM1  ;
 logic signed [31:0] O1_N4_S0;		always @(posedge clk) O1_N4_S0 <=     O1_I6_R0_C0_SM1   +  O1_I7_R0_C0_SM1  ;
 logic signed [31:0] O1_N6_S0;		always @(posedge clk) O1_N6_S0 <=     O1_I9_R0_C0_SM1   +  O1_I11_R0_C0_SM1  ;
 logic signed [31:0] O1_N8_S0;		always @(posedge clk) O1_N8_S0 <=     O1_I12_R0_C0_SM1   +  O1_I13_R0_C0_SM1  ;
 logic signed [31:0] O1_N10_S0;		always @(posedge clk) O1_N10_S0 <=     O1_I14_R0_C0_SM1   +  O1_I15_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O1_N0_S1;		always @(posedge clk) O1_N0_S1 <=     O1_N0_S0  +  O1_N2_S0 ;
 logic signed [31:0] O1_N2_S1;		always @(posedge clk) O1_N2_S1 <=     O1_N4_S0  +  O1_N6_S0 ;
 logic signed [31:0] O1_N4_S1;		always @(posedge clk) O1_N4_S1 <=     O1_N8_S0  +  O1_N10_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O1_N0_S2;		always @(posedge clk) O1_N0_S2 <=     O1_N0_S1  +  O1_N2_S1 ;
 logic signed [31:0] O1_N2_S2;		always @(posedge clk) O1_N2_S2 <=     O1_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O1_N0_S3;		always @(posedge clk) O1_N0_S3 <=     O1_N0_S2  +  O1_N2_S2 ;
 assign conv_mac_1 = O1_N0_S3;

logic signed [31:0] conv_mac_2;
logic signed [31:0] O2_N0_S0;		always @(posedge clk) O2_N0_S0 <=     O2_I0_R0_C0_SM1   +  O2_I1_R0_C0_SM1  ;
 logic signed [31:0] O2_N2_S0;		always @(posedge clk) O2_N2_S0 <=     O2_I2_R0_C0_SM1   +  O2_I3_R0_C0_SM1  ;
 logic signed [31:0] O2_N4_S0;		always @(posedge clk) O2_N4_S0 <=     O2_I4_R0_C0_SM1   +  O2_I5_R0_C0_SM1  ;
 logic signed [31:0] O2_N6_S0;		always @(posedge clk) O2_N6_S0 <=     O2_I6_R0_C0_SM1   +  O2_I7_R0_C0_SM1  ;
 logic signed [31:0] O2_N8_S0;		always @(posedge clk) O2_N8_S0 <=     O2_I8_R0_C0_SM1   +  O2_I9_R0_C0_SM1  ;
 logic signed [31:0] O2_N10_S0;		always @(posedge clk) O2_N10_S0 <=     O2_I11_R0_C0_SM1   +  O2_I14_R0_C0_SM1  ;
 logic signed [31:0] O2_N12_S0;		always @(posedge clk) O2_N12_S0 <=     O2_I15_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O2_N0_S1;		always @(posedge clk) O2_N0_S1 <=     O2_N0_S0  +  O2_N2_S0 ;
 logic signed [31:0] O2_N2_S1;		always @(posedge clk) O2_N2_S1 <=     O2_N4_S0  +  O2_N6_S0 ;
 logic signed [31:0] O2_N4_S1;		always @(posedge clk) O2_N4_S1 <=     O2_N8_S0  +  O2_N10_S0 ;
 logic signed [31:0] O2_N6_S1;		always @(posedge clk) O2_N6_S1 <=     O2_N12_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O2_N0_S2;		always @(posedge clk) O2_N0_S2 <=     O2_N0_S1  +  O2_N2_S1 ;
 logic signed [31:0] O2_N2_S2;		always @(posedge clk) O2_N2_S2 <=     O2_N4_S1  +  O2_N6_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O2_N0_S3;		always @(posedge clk) O2_N0_S3 <=     O2_N0_S2  +  O2_N2_S2 ;
 assign conv_mac_2 = O2_N0_S3;

logic signed [31:0] conv_mac_3;
logic signed [31:0] O3_N0_S0;		always @(posedge clk) O3_N0_S0 <=     O3_I1_R0_C0_SM1   +  O3_I4_R0_C0_SM1  ;
 logic signed [31:0] O3_N2_S0;		always @(posedge clk) O3_N2_S0 <=     O3_I5_R0_C0_SM1   +  O3_I6_R0_C0_SM1  ;
 logic signed [31:0] O3_N4_S0;		always @(posedge clk) O3_N4_S0 <=     O3_I9_R0_C0_SM1   +  O3_I13_R0_C0_SM1  ;
 logic signed [31:0] O3_N6_S0;		always @(posedge clk) O3_N6_S0 <=     O3_I14_R0_C0_SM1   +  O3_I15_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O3_N0_S1;		always @(posedge clk) O3_N0_S1 <=     O3_N0_S0  +  O3_N2_S0 ;
 logic signed [31:0] O3_N2_S1;		always @(posedge clk) O3_N2_S1 <=     O3_N4_S0  +  O3_N6_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O3_N0_S2;		always @(posedge clk) O3_N0_S2 <=     O3_N0_S1  +  O3_N2_S1 ;
 assign conv_mac_3 = O3_N0_S2;

logic signed [31:0] conv_mac_4;
logic signed [31:0] O4_N0_S0;		always @(posedge clk) O4_N0_S0 <=     O4_I1_R0_C0_SM1   +  O4_I2_R0_C0_SM1  ;
 logic signed [31:0] O4_N2_S0;		always @(posedge clk) O4_N2_S0 <=     O4_I3_R0_C0_SM1   +  O4_I5_R0_C0_SM1  ;
 logic signed [31:0] O4_N4_S0;		always @(posedge clk) O4_N4_S0 <=     O4_I6_R0_C0_SM1   +  O4_I9_R0_C0_SM1  ;
 logic signed [31:0] O4_N6_S0;		always @(posedge clk) O4_N6_S0 <=     O4_I13_R0_C0_SM1   +  O4_I14_R0_C0_SM1  ;
 logic signed [31:0] O4_N8_S0;		always @(posedge clk) O4_N8_S0 <=     O4_I15_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O4_N0_S1;		always @(posedge clk) O4_N0_S1 <=     O4_N0_S0  +  O4_N2_S0 ;
 logic signed [31:0] O4_N2_S1;		always @(posedge clk) O4_N2_S1 <=     O4_N4_S0  +  O4_N6_S0 ;
 logic signed [31:0] O4_N4_S1;		always @(posedge clk) O4_N4_S1 <=     O4_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O4_N0_S2;		always @(posedge clk) O4_N0_S2 <=     O4_N0_S1  +  O4_N2_S1 ;
 logic signed [31:0] O4_N2_S2;		always @(posedge clk) O4_N2_S2 <=     O4_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O4_N0_S3;		always @(posedge clk) O4_N0_S3 <=     O4_N0_S2  +  O4_N2_S2 ;
 assign conv_mac_4 = O4_N0_S3;

logic signed [31:0] conv_mac_5;
logic signed [31:0] O5_N0_S0;		always @(posedge clk) O5_N0_S0 <=     O5_I0_R0_C0_SM1   +  O5_I3_R0_C0_SM1  ;
 logic signed [31:0] O5_N2_S0;		always @(posedge clk) O5_N2_S0 <=     O5_I4_R0_C0_SM1   +  O5_I5_R0_C0_SM1  ;
 logic signed [31:0] O5_N4_S0;		always @(posedge clk) O5_N4_S0 <=     O5_I7_R0_C0_SM1   +  O5_I10_R0_C0_SM1  ;
 logic signed [31:0] O5_N6_S0;		always @(posedge clk) O5_N6_S0 <=     O5_I13_R0_C0_SM1   +  O5_I14_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O5_N0_S1;		always @(posedge clk) O5_N0_S1 <=     O5_N0_S0  +  O5_N2_S0 ;
 logic signed [31:0] O5_N2_S1;		always @(posedge clk) O5_N2_S1 <=     O5_N4_S0  +  O5_N6_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O5_N0_S2;		always @(posedge clk) O5_N0_S2 <=     O5_N0_S1  +  O5_N2_S1 ;
 assign conv_mac_5 = O5_N0_S2;

logic signed [31:0] conv_mac_6;
logic signed [31:0] O6_N0_S0;		always @(posedge clk) O6_N0_S0 <=     O6_I0_R0_C0_SM1   +  O6_I1_R0_C0_SM1  ;
 logic signed [31:0] O6_N2_S0;		always @(posedge clk) O6_N2_S0 <=     O6_I2_R0_C0_SM1   +  O6_I6_R0_C0_SM1  ;
 logic signed [31:0] O6_N4_S0;		always @(posedge clk) O6_N4_S0 <=     O6_I8_R0_C0_SM1   +  O6_I9_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O6_N0_S1;		always @(posedge clk) O6_N0_S1 <=     O6_N0_S0  +  O6_N2_S0 ;
 logic signed [31:0] O6_N2_S1;		always @(posedge clk) O6_N2_S1 <=     O6_N4_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O6_N0_S2;		always @(posedge clk) O6_N0_S2 <=     O6_N0_S1  +  O6_N2_S1 ;
 assign conv_mac_6 = O6_N0_S2;

logic signed [31:0] conv_mac_7;
logic signed [31:0] O7_N0_S0;		always @(posedge clk) O7_N0_S0 <=     O7_I0_R0_C0_SM1   +  O7_I2_R0_C0_SM1  ;
 logic signed [31:0] O7_N2_S0;		always @(posedge clk) O7_N2_S0 <=     O7_I3_R0_C0_SM1   +  O7_I4_R0_C0_SM1  ;
 logic signed [31:0] O7_N4_S0;		always @(posedge clk) O7_N4_S0 <=     O7_I5_R0_C0_SM1   +  O7_I7_R0_C0_SM1  ;
 logic signed [31:0] O7_N6_S0;		always @(posedge clk) O7_N6_S0 <=     O7_I10_R0_C0_SM1   +  O7_I13_R0_C0_SM1  ;
 logic signed [31:0] O7_N8_S0;		always @(posedge clk) O7_N8_S0 <=     O7_I14_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O7_N0_S1;		always @(posedge clk) O7_N0_S1 <=     O7_N0_S0  +  O7_N2_S0 ;
 logic signed [31:0] O7_N2_S1;		always @(posedge clk) O7_N2_S1 <=     O7_N4_S0  +  O7_N6_S0 ;
 logic signed [31:0] O7_N4_S1;		always @(posedge clk) O7_N4_S1 <=     O7_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O7_N0_S2;		always @(posedge clk) O7_N0_S2 <=     O7_N0_S1  +  O7_N2_S1 ;
 logic signed [31:0] O7_N2_S2;		always @(posedge clk) O7_N2_S2 <=     O7_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O7_N0_S3;		always @(posedge clk) O7_N0_S3 <=     O7_N0_S2  +  O7_N2_S2 ;
 assign conv_mac_7 = O7_N0_S3;

logic signed [31:0] conv_mac_8;
logic signed [31:0] O8_N0_S0;		always @(posedge clk) O8_N0_S0 <=     O8_I1_R0_C0_SM1   +  O8_I5_R0_C0_SM1  ;
 logic signed [31:0] O8_N2_S0;		always @(posedge clk) O8_N2_S0 <=     O8_I6_R0_C0_SM1   +  O8_I9_R0_C0_SM1  ;
 logic signed [31:0] O8_N4_S0;		always @(posedge clk) O8_N4_S0 <=     O8_I12_R0_C0_SM1   +  O8_I13_R0_C0_SM1  ;
 logic signed [31:0] O8_N6_S0;		always @(posedge clk) O8_N6_S0 <=     O8_I15_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O8_N0_S1;		always @(posedge clk) O8_N0_S1 <=     O8_N0_S0  +  O8_N2_S0 ;
 logic signed [31:0] O8_N2_S1;		always @(posedge clk) O8_N2_S1 <=     O8_N4_S0  +  O8_N6_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O8_N0_S2;		always @(posedge clk) O8_N0_S2 <=     O8_N0_S1  +  O8_N2_S1 ;
 assign conv_mac_8 = O8_N0_S2;

logic signed [31:0] conv_mac_9;
logic signed [31:0] O9_N0_S0;		always @(posedge clk) O9_N0_S0 <=     O9_I3_R0_C0_SM1   +  O9_I4_R0_C0_SM1  ;
 logic signed [31:0] O9_N2_S0;		always @(posedge clk) O9_N2_S0 <=     O9_I5_R0_C0_SM1   +  O9_I10_R0_C0_SM1  ;
 logic signed [31:0] O9_N4_S0;		always @(posedge clk) O9_N4_S0 <=     O9_I13_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O9_N0_S1;		always @(posedge clk) O9_N0_S1 <=     O9_N0_S0  +  O9_N2_S0 ;
 logic signed [31:0] O9_N2_S1;		always @(posedge clk) O9_N2_S1 <=     O9_N4_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O9_N0_S2;		always @(posedge clk) O9_N0_S2 <=     O9_N0_S1  +  O9_N2_S1 ;
 assign conv_mac_9 = O9_N0_S2;

logic signed [31:0] conv_mac_10;
logic signed [31:0] O10_N0_S0;		always @(posedge clk) O10_N0_S0 <=     O10_I3_R0_C0_SM1   +  O10_I5_R0_C0_SM1  ;
 logic signed [31:0] O10_N2_S0;		always @(posedge clk) O10_N2_S0 <=     O10_I6_R0_C0_SM1   +  O10_I7_R0_C0_SM1  ;
 logic signed [31:0] O10_N4_S0;		always @(posedge clk) O10_N4_S0 <=     O10_I10_R0_C0_SM1   +  O10_I11_R0_C0_SM1  ;
 logic signed [31:0] O10_N6_S0;		always @(posedge clk) O10_N6_S0 <=     O10_I14_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O10_N0_S1;		always @(posedge clk) O10_N0_S1 <=     O10_N0_S0  +  O10_N2_S0 ;
 logic signed [31:0] O10_N2_S1;		always @(posedge clk) O10_N2_S1 <=     O10_N4_S0  +  O10_N6_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O10_N0_S2;		always @(posedge clk) O10_N0_S2 <=     O10_N0_S1  +  O10_N2_S1 ;
 assign conv_mac_10 = O10_N0_S2;

logic signed [31:0] conv_mac_11;
logic signed [31:0] O11_N0_S0;		always @(posedge clk) O11_N0_S0 <=     O11_I1_R0_C0_SM1   +  O11_I3_R0_C0_SM1  ;
 logic signed [31:0] O11_N2_S0;		always @(posedge clk) O11_N2_S0 <=     O11_I4_R0_C0_SM1   +  O11_I8_R0_C0_SM1  ;
 logic signed [31:0] O11_N4_S0;		always @(posedge clk) O11_N4_S0 <=     O11_I9_R0_C0_SM1   +  O11_I11_R0_C0_SM1  ;
 logic signed [31:0] O11_N6_S0;		always @(posedge clk) O11_N6_S0 <=     O11_I12_R0_C0_SM1   +  O11_I14_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O11_N0_S1;		always @(posedge clk) O11_N0_S1 <=     O11_N0_S0  +  O11_N2_S0 ;
 logic signed [31:0] O11_N2_S1;		always @(posedge clk) O11_N2_S1 <=     O11_N4_S0  +  O11_N6_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O11_N0_S2;		always @(posedge clk) O11_N0_S2 <=     O11_N0_S1  +  O11_N2_S1 ;
 assign conv_mac_11 = O11_N0_S2;

logic signed [31:0] conv_mac_12;
logic signed [31:0] O12_N0_S0;		always @(posedge clk) O12_N0_S0 <=     O12_I2_R0_C0_SM1   +  O12_I3_R0_C0_SM1  ;
 logic signed [31:0] O12_N2_S0;		always @(posedge clk) O12_N2_S0 <=     O12_I4_R0_C0_SM1   +  O12_I5_R0_C0_SM1  ;
 logic signed [31:0] O12_N4_S0;		always @(posedge clk) O12_N4_S0 <=     O12_I6_R0_C0_SM1   +  O12_I7_R0_C0_SM1  ;
 logic signed [31:0] O12_N6_S0;		always @(posedge clk) O12_N6_S0 <=     O12_I10_R0_C0_SM1   +  O12_I11_R0_C0_SM1  ;
 logic signed [31:0] O12_N8_S0;		always @(posedge clk) O12_N8_S0 <=     O12_I12_R0_C0_SM1   +  O12_I13_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O12_N0_S1;		always @(posedge clk) O12_N0_S1 <=     O12_N0_S0  +  O12_N2_S0 ;
 logic signed [31:0] O12_N2_S1;		always @(posedge clk) O12_N2_S1 <=     O12_N4_S0  +  O12_N6_S0 ;
 logic signed [31:0] O12_N4_S1;		always @(posedge clk) O12_N4_S1 <=     O12_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O12_N0_S2;		always @(posedge clk) O12_N0_S2 <=     O12_N0_S1  +  O12_N2_S1 ;
 logic signed [31:0] O12_N2_S2;		always @(posedge clk) O12_N2_S2 <=     O12_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O12_N0_S3;		always @(posedge clk) O12_N0_S3 <=     O12_N0_S2  +  O12_N2_S2 ;
 assign conv_mac_12 = O12_N0_S3;

logic signed [31:0] conv_mac_13;
logic signed [31:0] O13_N0_S0;		always @(posedge clk) O13_N0_S0 <=     O13_I1_R0_C0_SM1   +  O13_I2_R0_C0_SM1  ;
 logic signed [31:0] O13_N2_S0;		always @(posedge clk) O13_N2_S0 <=     O13_I4_R0_C0_SM1   +  O13_I6_R0_C0_SM1  ;
 logic signed [31:0] O13_N4_S0;		always @(posedge clk) O13_N4_S0 <=     O13_I8_R0_C0_SM1   +  O13_I11_R0_C0_SM1  ;
 logic signed [31:0] O13_N6_S0;		always @(posedge clk) O13_N6_S0 <=     O13_I12_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O13_N0_S1;		always @(posedge clk) O13_N0_S1 <=     O13_N0_S0  +  O13_N2_S0 ;
 logic signed [31:0] O13_N2_S1;		always @(posedge clk) O13_N2_S1 <=     O13_N4_S0  +  O13_N6_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O13_N0_S2;		always @(posedge clk) O13_N0_S2 <=     O13_N0_S1  +  O13_N2_S1 ;
 assign conv_mac_13 = O13_N0_S2;

logic signed [31:0] conv_mac_14;
logic signed [31:0] O14_N0_S0;		always @(posedge clk) O14_N0_S0 <=     O14_I0_R0_C0_SM1   +  O14_I1_R0_C0_SM1  ;
 logic signed [31:0] O14_N2_S0;		always @(posedge clk) O14_N2_S0 <=     O14_I2_R0_C0_SM1   +  O14_I3_R0_C0_SM1  ;
 logic signed [31:0] O14_N4_S0;		always @(posedge clk) O14_N4_S0 <=     O14_I6_R0_C0_SM1   +  O14_I7_R0_C0_SM1  ;
 logic signed [31:0] O14_N6_S0;		always @(posedge clk) O14_N6_S0 <=     O14_I9_R0_C0_SM1   +  O14_I14_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O14_N0_S1;		always @(posedge clk) O14_N0_S1 <=     O14_N0_S0  +  O14_N2_S0 ;
 logic signed [31:0] O14_N2_S1;		always @(posedge clk) O14_N2_S1 <=     O14_N4_S0  +  O14_N6_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O14_N0_S2;		always @(posedge clk) O14_N0_S2 <=     O14_N0_S1  +  O14_N2_S1 ;
 assign conv_mac_14 = O14_N0_S2;

logic signed [31:0] conv_mac_15;
logic signed [31:0] O15_N0_S0;		always @(posedge clk) O15_N0_S0 <=     O15_I0_R0_C0_SM1   +  O15_I1_R0_C0_SM1  ;
 logic signed [31:0] O15_N2_S0;		always @(posedge clk) O15_N2_S0 <=     O15_I2_R0_C0_SM1   +  O15_I3_R0_C0_SM1  ;
 logic signed [31:0] O15_N4_S0;		always @(posedge clk) O15_N4_S0 <=     O15_I4_R0_C0_SM1   +  O15_I5_R0_C0_SM1  ;
 logic signed [31:0] O15_N6_S0;		always @(posedge clk) O15_N6_S0 <=     O15_I6_R0_C0_SM1   +  O15_I7_R0_C0_SM1  ;
 logic signed [31:0] O15_N8_S0;		always @(posedge clk) O15_N8_S0 <=     O15_I8_R0_C0_SM1   +  O15_I9_R0_C0_SM1  ;
 logic signed [31:0] O15_N10_S0;		always @(posedge clk) O15_N10_S0 <=     O15_I11_R0_C0_SM1   +  O15_I12_R0_C0_SM1  ;
 logic signed [31:0] O15_N12_S0;		always @(posedge clk) O15_N12_S0 <=     O15_I13_R0_C0_SM1   +  O15_I15_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O15_N0_S1;		always @(posedge clk) O15_N0_S1 <=     O15_N0_S0  +  O15_N2_S0 ;
 logic signed [31:0] O15_N2_S1;		always @(posedge clk) O15_N2_S1 <=     O15_N4_S0  +  O15_N6_S0 ;
 logic signed [31:0] O15_N4_S1;		always @(posedge clk) O15_N4_S1 <=     O15_N8_S0  +  O15_N10_S0 ;
 logic signed [31:0] O15_N6_S1;		always @(posedge clk) O15_N6_S1 <=     O15_N12_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O15_N0_S2;		always @(posedge clk) O15_N0_S2 <=     O15_N0_S1  +  O15_N2_S1 ;
 logic signed [31:0] O15_N2_S2;		always @(posedge clk) O15_N2_S2 <=     O15_N4_S1  +  O15_N6_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O15_N0_S3;		always @(posedge clk) O15_N0_S3 <=     O15_N0_S2  +  O15_N2_S2 ;
 assign conv_mac_15 = O15_N0_S3;

logic valid_D1;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D1<= 0 ;
	else valid_D1<=valid;
end
logic valid_D2;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D2<= 0 ;
	else valid_D2<=valid_D1;
end
logic valid_D3;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D3<= 0 ;
	else valid_D3<=valid_D2;
end
logic valid_D4;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D4<= 0 ;
	else valid_D4<=valid_D3;
end
logic valid_D5;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D5<= 0 ;
	else valid_D5<=valid_D4;
end
always_ff @(posedge clk) begin
	if (rstn == 0) ready <= 0 ;
	else ready <=valid_D5;
end
logic [31:0] bias_add_0;
assign bias_add_0 = conv_mac_0 + 7'd35;
logic [31:0] bias_add_1;
assign bias_add_1 = conv_mac_1 + 7'd40;
logic [31:0] bias_add_2;
assign bias_add_2 = conv_mac_2 - 4'd5;
logic [31:0] bias_add_3;
assign bias_add_3 = conv_mac_3 - 7'd39;
logic [31:0] bias_add_4;
assign bias_add_4 = conv_mac_4 + 2'd1;
logic [31:0] bias_add_5;
assign bias_add_5 = conv_mac_5 + 7'd32;
logic [31:0] bias_add_6;
assign bias_add_6 = conv_mac_6 - 2'd1;
logic [31:0] bias_add_7;
assign bias_add_7 = conv_mac_7 + 7'd37;
logic [31:0] bias_add_8;
assign bias_add_8 = conv_mac_8 + 5'd11;
logic [31:0] bias_add_9;
assign bias_add_9 = conv_mac_9 - 5'd10;
logic [31:0] bias_add_10;
assign bias_add_10 = conv_mac_10 - 3'd3;
logic [31:0] bias_add_11;
assign bias_add_11 = conv_mac_11 + 6'd23;
logic [31:0] bias_add_12;
assign bias_add_12 = conv_mac_12 + 7'd40;
logic [31:0] bias_add_13;
assign bias_add_13 = conv_mac_13 + 5'd9;
logic [31:0] bias_add_14;
assign bias_add_14 = conv_mac_14 + 6'd25;
logic [31:0] bias_add_15;
assign bias_add_15 = conv_mac_15 + 6'd18;

logic [7:0] relu_0;
assign relu_0[7:0] = (bias_add_0[31]==0) ? ((bias_add_0<3'd6) ? {{bias_add_0[31],bias_add_0[10:4]}} :'d6) : '0;
logic [7:0] relu_1;
assign relu_1[7:0] = (bias_add_1[31]==0) ? ((bias_add_1<3'd6) ? {{bias_add_1[31],bias_add_1[10:4]}} :'d6) : '0;
logic [7:0] relu_2;
assign relu_2[7:0] = (bias_add_2[31]==0) ? ((bias_add_2<3'd6) ? {{bias_add_2[31],bias_add_2[10:4]}} :'d6) : '0;
logic [7:0] relu_3;
assign relu_3[7:0] = (bias_add_3[31]==0) ? ((bias_add_3<3'd6) ? {{bias_add_3[31],bias_add_3[10:4]}} :'d6) : '0;
logic [7:0] relu_4;
assign relu_4[7:0] = (bias_add_4[31]==0) ? ((bias_add_4<3'd6) ? {{bias_add_4[31],bias_add_4[10:4]}} :'d6) : '0;
logic [7:0] relu_5;
assign relu_5[7:0] = (bias_add_5[31]==0) ? ((bias_add_5<3'd6) ? {{bias_add_5[31],bias_add_5[10:4]}} :'d6) : '0;
logic [7:0] relu_6;
assign relu_6[7:0] = (bias_add_6[31]==0) ? ((bias_add_6<3'd6) ? {{bias_add_6[31],bias_add_6[10:4]}} :'d6) : '0;
logic [7:0] relu_7;
assign relu_7[7:0] = (bias_add_7[31]==0) ? ((bias_add_7<3'd6) ? {{bias_add_7[31],bias_add_7[10:4]}} :'d6) : '0;
logic [7:0] relu_8;
assign relu_8[7:0] = (bias_add_8[31]==0) ? ((bias_add_8<3'd6) ? {{bias_add_8[31],bias_add_8[10:4]}} :'d6) : '0;
logic [7:0] relu_9;
assign relu_9[7:0] = (bias_add_9[31]==0) ? ((bias_add_9<3'd6) ? {{bias_add_9[31],bias_add_9[10:4]}} :'d6) : '0;
logic [7:0] relu_10;
assign relu_10[7:0] = (bias_add_10[31]==0) ? ((bias_add_10<3'd6) ? {{bias_add_10[31],bias_add_10[10:4]}} :'d6) : '0;
logic [7:0] relu_11;
assign relu_11[7:0] = (bias_add_11[31]==0) ? ((bias_add_11<3'd6) ? {{bias_add_11[31],bias_add_11[10:4]}} :'d6) : '0;
logic [7:0] relu_12;
assign relu_12[7:0] = (bias_add_12[31]==0) ? ((bias_add_12<3'd6) ? {{bias_add_12[31],bias_add_12[10:4]}} :'d6) : '0;
logic [7:0] relu_13;
assign relu_13[7:0] = (bias_add_13[31]==0) ? ((bias_add_13<3'd6) ? {{bias_add_13[31],bias_add_13[10:4]}} :'d6) : '0;
logic [7:0] relu_14;
assign relu_14[7:0] = (bias_add_14[31]==0) ? ((bias_add_14<3'd6) ? {{bias_add_14[31],bias_add_14[10:4]}} :'d6) : '0;
logic [7:0] relu_15;
assign relu_15[7:0] = (bias_add_15[31]==0) ? ((bias_add_15<3'd6) ? {{bias_add_15[31],bias_add_15[10:4]}} :'d6) : '0;

assign output_act = {
	relu_15,
	relu_14,
	relu_13,
	relu_12,
	relu_11,
	relu_10,
	relu_9,
	relu_8,
	relu_7,
	relu_6,
	relu_5,
	relu_4,
	relu_3,
	relu_2,
	relu_1,
	relu_0
};

endmodule
module conv4_pw (
    input logic clk,
    input logic rstn,
    input logic valid,
    input logic [128-1:0] input_act,
    output logic [256-1:0] output_act,
    output logic ready
);
logic we;
logic [8:0] zero_number; 
assign zero_number = 9'd0; 
//1
logic [128-1:0] input_act_ff ;
always_ff @(posedge clk) begin
    if (rstn == 0) begin
        input_act_ff <= '0;
      //  ready <= '0;
    end
    else begin
        input_act_ff <= input_act;
     //   ready <= valid;
    end
end
logic [7:0] input_fmap_0;
assign input_fmap_0 = input_act_ff[7:0];
logic [7:0] input_fmap_1;
assign input_fmap_1 = input_act_ff[15:8];
logic [7:0] input_fmap_2;
assign input_fmap_2 = input_act_ff[23:16];
logic [7:0] input_fmap_3;
assign input_fmap_3 = input_act_ff[31:24];
logic [7:0] input_fmap_4;
assign input_fmap_4 = input_act_ff[39:32];
logic [7:0] input_fmap_5;
assign input_fmap_5 = input_act_ff[47:40];
logic [7:0] input_fmap_6;
assign input_fmap_6 = input_act_ff[55:48];
logic [7:0] input_fmap_7;
assign input_fmap_7 = input_act_ff[63:56];
logic [7:0] input_fmap_8;
assign input_fmap_8 = input_act_ff[71:64];
logic [7:0] input_fmap_9;
assign input_fmap_9 = input_act_ff[79:72];
logic [7:0] input_fmap_10;
assign input_fmap_10 = input_act_ff[87:80];
logic [7:0] input_fmap_11;
assign input_fmap_11 = input_act_ff[95:88];
logic [7:0] input_fmap_12;
assign input_fmap_12 = input_act_ff[103:96];
logic [7:0] input_fmap_13;
assign input_fmap_13 = input_act_ff[111:104];
logic [7:0] input_fmap_14;
assign input_fmap_14 = input_act_ff[119:112];
logic [7:0] input_fmap_15;
assign input_fmap_15 = input_act_ff[127:120];

logic [10-1:0] O0_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O0_I0_R0_C01_rom_inst (.q(O0_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O0_I0_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O0_I0_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O0_I0_R0_C01_rom_inst (.q(O0_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [10-1:0] O0_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O0_I2_R0_C01_rom_inst (.q(O0_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O0_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O0_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O0_I2_R0_C01_rom_inst (.q(O0_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [10-1:0] O0_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O0_I5_R0_C01_rom_inst (.q(O0_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I5_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O0_I5_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O0_I5_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O0_I5_R0_C01_rom_inst (.q(O0_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [10-1:0] O0_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O0_I15_R0_C01_rom_inst (.q(O0_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I15_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O0_I15_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O0_I15_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O0_I15_R0_C01_rom_inst (.q(O0_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [11-1:0] O1_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O1_I0_R0_C03_rom_inst (.q(O1_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I0_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O1_I0_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O1_I0_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O1_I0_R0_C03_rom_inst (.q(O1_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [11-1:0] O1_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O1_I1_R0_C02_rom_inst (.q(O1_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I1_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O1_I1_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O1_I1_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O1_I1_R0_C02_rom_inst (.q(O1_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [11-1:0] O1_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O1_I2_R0_C02_rom_inst (.q(O1_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I2_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O1_I2_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O1_I2_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O1_I2_R0_C02_rom_inst (.q(O1_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [11-1:0] O1_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O1_I5_R0_C02_rom_inst (.q(O1_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I5_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O1_I5_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O1_I5_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O1_I5_R0_C02_rom_inst (.q(O1_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [10-1:0] O1_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O1_I6_R0_C01_rom_inst (.q(O1_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I6_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O1_I6_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O1_I6_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O1_I6_R0_C01_rom_inst (.q(O1_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [10-1:0] O1_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O1_I7_R0_C01_rom_inst (.q(O1_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I7_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O1_I7_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O1_I7_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O1_I7_R0_C01_rom_inst (.q(O1_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [10-1:0] O1_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O1_I8_R0_C01_rom_inst (.q(O1_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I8_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O1_I8_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O1_I8_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O1_I8_R0_C01_rom_inst (.q(O1_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [10-1:0] O1_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O1_I9_R0_C01_rom_inst (.q(O1_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I9_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O1_I9_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O1_I9_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O1_I9_R0_C01_rom_inst (.q(O1_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [10-1:0] O1_I14_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O1_I14_R0_C01_rom_inst (.q(O1_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I14_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O1_I14_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O1_I14_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O1_I14_R0_C01_rom_inst (.q(O1_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clock  (clk));
logic [10-1:0] O1_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O1_I15_R0_C01_rom_inst (.q(O1_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I15_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O1_I15_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O1_I15_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O1_I15_R0_C01_rom_inst (.q(O1_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [11-1:0] O2_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O2_I1_R0_C02_rom_inst (.q(O2_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O2_I1_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O2_I1_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O2_I1_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O2_I1_R0_C02_rom_inst (.q(O2_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [10-1:0] O2_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O2_I2_R0_C01_rom_inst (.q(O2_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O2_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O2_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O2_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O2_I2_R0_C01_rom_inst (.q(O2_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [10-1:0] O2_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O2_I4_R0_C01_rom_inst (.q(O2_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O2_I4_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O2_I4_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O2_I4_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O2_I4_R0_C01_rom_inst (.q(O2_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [12-1:0] O2_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_pw_O2_I6_R0_C04_rom_inst (.q(O2_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O2_I6_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O2_I6_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O2_I6_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_pw_O2_I6_R0_C04_rom_inst (.q(O2_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [10-1:0] O2_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O2_I7_R0_C01_rom_inst (.q(O2_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O2_I7_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O2_I7_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O2_I7_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O2_I7_R0_C01_rom_inst (.q(O2_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [11-1:0] O2_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O2_I11_R0_C03_rom_inst (.q(O2_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O2_I11_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O2_I11_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O2_I11_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O2_I11_R0_C03_rom_inst (.q(O2_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [10-1:0] O2_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O2_I15_R0_C01_rom_inst (.q(O2_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O2_I15_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O2_I15_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O2_I15_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O2_I15_R0_C01_rom_inst (.q(O2_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [11-1:0] O3_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O3_I0_R0_C02_rom_inst (.q(O3_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I0_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O3_I0_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O3_I0_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O3_I0_R0_C02_rom_inst (.q(O3_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [11-1:0] O3_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O3_I2_R0_C02_rom_inst (.q(O3_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I2_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O3_I2_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O3_I2_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O3_I2_R0_C02_rom_inst (.q(O3_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [10-1:0] O3_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O3_I4_R0_C01_rom_inst (.q(O3_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I4_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O3_I4_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O3_I4_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O3_I4_R0_C01_rom_inst (.q(O3_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [11-1:0] O3_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O3_I5_R0_C02_rom_inst (.q(O3_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I5_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O3_I5_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O3_I5_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O3_I5_R0_C02_rom_inst (.q(O3_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [10-1:0] O3_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O3_I6_R0_C01_rom_inst (.q(O3_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I6_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O3_I6_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O3_I6_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O3_I6_R0_C01_rom_inst (.q(O3_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [10-1:0] O3_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O3_I7_R0_C01_rom_inst (.q(O3_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I7_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O3_I7_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O3_I7_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O3_I7_R0_C01_rom_inst (.q(O3_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [11-1:0] O3_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O3_I8_R0_C03_rom_inst (.q(O3_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I8_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O3_I8_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O3_I8_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O3_I8_R0_C03_rom_inst (.q(O3_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [11-1:0] O3_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O3_I9_R0_C03_rom_inst (.q(O3_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I9_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O3_I9_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O3_I9_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O3_I9_R0_C03_rom_inst (.q(O3_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [10-1:0] O3_I10_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O3_I10_R0_C01_rom_inst (.q(O3_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I10_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O3_I10_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O3_I10_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O3_I10_R0_C01_rom_inst (.q(O3_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clock  (clk));
logic [11-1:0] O3_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O3_I12_R0_C02_rom_inst (.q(O3_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I12_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O3_I12_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O3_I12_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O3_I12_R0_C02_rom_inst (.q(O3_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [11-1:0] O3_I14_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O3_I14_R0_C02_rom_inst (.q(O3_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I14_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O3_I14_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O3_I14_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O3_I14_R0_C02_rom_inst (.q(O3_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clock  (clk));
logic [10-1:0] O3_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O3_I15_R0_C01_rom_inst (.q(O3_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I15_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O3_I15_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O3_I15_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O3_I15_R0_C01_rom_inst (.q(O3_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [11-1:0] O4_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O4_I0_R0_C03_rom_inst (.q(O4_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I0_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O4_I0_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O4_I0_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O4_I0_R0_C03_rom_inst (.q(O4_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [12-1:0] O4_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_pw_O4_I1_R0_C05_rom_inst (.q(O4_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I1_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O4_I1_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O4_I1_R0_C05_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_pw_O4_I1_R0_C05_rom_inst (.q(O4_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [10-1:0] O4_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O4_I3_R0_C01_rom_inst (.q(O4_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I3_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I3_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O4_I3_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O4_I3_R0_C01_rom_inst (.q(O4_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [10-1:0] O4_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O4_I4_R0_C01_rom_inst (.q(O4_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I4_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O4_I4_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O4_I4_R0_C01_rom_inst (.q(O4_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [11-1:0] O4_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O4_I5_R0_C03_rom_inst (.q(O4_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I5_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O4_I5_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O4_I5_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O4_I5_R0_C03_rom_inst (.q(O4_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [11-1:0] O4_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O4_I7_R0_C02_rom_inst (.q(O4_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I7_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O4_I7_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O4_I7_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O4_I7_R0_C02_rom_inst (.q(O4_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [11-1:0] O4_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O4_I8_R0_C03_rom_inst (.q(O4_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I8_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O4_I8_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O4_I8_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O4_I8_R0_C03_rom_inst (.q(O4_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [11-1:0] O4_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O4_I9_R0_C02_rom_inst (.q(O4_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I9_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O4_I9_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O4_I9_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O4_I9_R0_C02_rom_inst (.q(O4_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [11-1:0] O4_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O4_I11_R0_C03_rom_inst (.q(O4_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I11_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O4_I11_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O4_I11_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O4_I11_R0_C03_rom_inst (.q(O4_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [11-1:0] O4_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O4_I12_R0_C02_rom_inst (.q(O4_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I12_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O4_I12_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O4_I12_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O4_I12_R0_C02_rom_inst (.q(O4_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [11-1:0] O4_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O4_I13_R0_C03_rom_inst (.q(O4_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I13_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O4_I13_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O4_I13_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O4_I13_R0_C03_rom_inst (.q(O4_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [10-1:0] O4_I14_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O4_I14_R0_C01_rom_inst (.q(O4_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I14_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I14_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O4_I14_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O4_I14_R0_C01_rom_inst (.q(O4_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clock  (clk));
logic [10-1:0] O4_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O4_I15_R0_C01_rom_inst (.q(O4_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I15_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I15_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O4_I15_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O4_I15_R0_C01_rom_inst (.q(O4_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [10-1:0] O5_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O5_I1_R0_C01_rom_inst (.q(O5_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I1_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I1_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O5_I1_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O5_I1_R0_C01_rom_inst (.q(O5_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [11-1:0] O5_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O5_I2_R0_C02_rom_inst (.q(O5_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I2_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O5_I2_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O5_I2_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O5_I2_R0_C02_rom_inst (.q(O5_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [10-1:0] O5_I10_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O5_I10_R0_C01_rom_inst (.q(O5_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I10_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I10_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O5_I10_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O5_I10_R0_C01_rom_inst (.q(O5_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clock  (clk));
logic [10-1:0] O5_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O5_I12_R0_C01_rom_inst (.q(O5_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I12_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I12_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O5_I12_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O5_I12_R0_C01_rom_inst (.q(O5_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [11-1:0] O5_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O5_I15_R0_C02_rom_inst (.q(O5_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I15_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O5_I15_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O5_I15_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O5_I15_R0_C02_rom_inst (.q(O5_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [11-1:0] O6_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O6_I0_R0_C02_rom_inst (.q(O6_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I0_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O6_I0_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O6_I0_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O6_I0_R0_C02_rom_inst (.q(O6_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [11-1:0] O6_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O6_I1_R0_C02_rom_inst (.q(O6_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I1_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O6_I1_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O6_I1_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O6_I1_R0_C02_rom_inst (.q(O6_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [10-1:0] O6_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O6_I2_R0_C01_rom_inst (.q(O6_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O6_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O6_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O6_I2_R0_C01_rom_inst (.q(O6_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [10-1:0] O6_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O6_I4_R0_C01_rom_inst (.q(O6_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I4_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O6_I4_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O6_I4_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O6_I4_R0_C01_rom_inst (.q(O6_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [11-1:0] O6_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O6_I5_R0_C02_rom_inst (.q(O6_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I5_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O6_I5_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O6_I5_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O6_I5_R0_C02_rom_inst (.q(O6_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [11-1:0] O6_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O6_I7_R0_C03_rom_inst (.q(O6_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I7_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O6_I7_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O6_I7_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O6_I7_R0_C03_rom_inst (.q(O6_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [11-1:0] O6_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O6_I8_R0_C02_rom_inst (.q(O6_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I8_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O6_I8_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O6_I8_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O6_I8_R0_C02_rom_inst (.q(O6_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [12-1:0] O6_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_pw_O6_I9_R0_C04_rom_inst (.q(O6_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I9_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O6_I9_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O6_I9_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_pw_O6_I9_R0_C04_rom_inst (.q(O6_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [11-1:0] O6_I10_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O6_I10_R0_C03_rom_inst (.q(O6_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I10_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O6_I10_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O6_I10_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O6_I10_R0_C03_rom_inst (.q(O6_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clock  (clk));
logic [10-1:0] O6_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O6_I12_R0_C01_rom_inst (.q(O6_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I12_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O6_I12_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O6_I12_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O6_I12_R0_C01_rom_inst (.q(O6_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [10-1:0] O6_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O6_I13_R0_C01_rom_inst (.q(O6_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I13_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O6_I13_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O6_I13_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O6_I13_R0_C01_rom_inst (.q(O6_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [10-1:0] O6_I14_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O6_I14_R0_C01_rom_inst (.q(O6_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I14_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O6_I14_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O6_I14_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O6_I14_R0_C01_rom_inst (.q(O6_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clock  (clk));
logic [11-1:0] O6_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O6_I15_R0_C03_rom_inst (.q(O6_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I15_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O6_I15_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O6_I15_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O6_I15_R0_C03_rom_inst (.q(O6_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [10-1:0] O7_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O7_I0_R0_C01_rom_inst (.q(O7_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I0_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O7_I0_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O7_I0_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O7_I0_R0_C01_rom_inst (.q(O7_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [10-1:0] O7_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O7_I2_R0_C01_rom_inst (.q(O7_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O7_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O7_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O7_I2_R0_C01_rom_inst (.q(O7_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [12-1:0] O7_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_pw_O7_I4_R0_C05_rom_inst (.q(O7_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I4_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O7_I4_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O7_I4_R0_C05_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_pw_O7_I4_R0_C05_rom_inst (.q(O7_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [11-1:0] O7_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O7_I5_R0_C02_rom_inst (.q(O7_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I5_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O7_I5_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O7_I5_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O7_I5_R0_C02_rom_inst (.q(O7_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [11-1:0] O7_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O7_I7_R0_C02_rom_inst (.q(O7_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I7_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O7_I7_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O7_I7_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O7_I7_R0_C02_rom_inst (.q(O7_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [10-1:0] O7_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O7_I8_R0_C01_rom_inst (.q(O7_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I8_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O7_I8_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O7_I8_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O7_I8_R0_C01_rom_inst (.q(O7_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [10-1:0] O7_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O7_I9_R0_C01_rom_inst (.q(O7_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I9_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O7_I9_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O7_I9_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O7_I9_R0_C01_rom_inst (.q(O7_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [10-1:0] O7_I10_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O7_I10_R0_C01_rom_inst (.q(O7_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I10_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O7_I10_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O7_I10_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O7_I10_R0_C01_rom_inst (.q(O7_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clock  (clk));
logic [10-1:0] O7_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O7_I11_R0_C01_rom_inst (.q(O7_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I11_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O7_I11_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O7_I11_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O7_I11_R0_C01_rom_inst (.q(O7_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [10-1:0] O7_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O7_I13_R0_C01_rom_inst (.q(O7_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I13_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O7_I13_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O7_I13_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O7_I13_R0_C01_rom_inst (.q(O7_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [11-1:0] O7_I14_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O7_I14_R0_C02_rom_inst (.q(O7_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I14_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O7_I14_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O7_I14_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O7_I14_R0_C02_rom_inst (.q(O7_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clock  (clk));
logic [10-1:0] O7_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O7_I15_R0_C01_rom_inst (.q(O7_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I15_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O7_I15_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O7_I15_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O7_I15_R0_C01_rom_inst (.q(O7_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [10-1:0] O8_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O8_I0_R0_C01_rom_inst (.q(O8_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O8_I0_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O8_I0_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O8_I0_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O8_I0_R0_C01_rom_inst (.q(O8_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [10-1:0] O8_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O8_I3_R0_C01_rom_inst (.q(O8_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O8_I3_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O8_I3_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O8_I3_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O8_I3_R0_C01_rom_inst (.q(O8_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [11-1:0] O8_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O8_I5_R0_C03_rom_inst (.q(O8_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O8_I5_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O8_I5_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O8_I5_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O8_I5_R0_C03_rom_inst (.q(O8_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [12-1:0] O8_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_pw_O8_I9_R0_C05_rom_inst (.q(O8_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O8_I9_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O8_I9_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O8_I9_R0_C05_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_pw_O8_I9_R0_C05_rom_inst (.q(O8_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [12-1:0] O8_I10_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_pw_O8_I10_R0_C06_rom_inst (.q(O8_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clk(clk),.d(0),.we(0));
//assign O8_I10_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O8_I10_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O8_I10_R0_C06_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_pw_O8_I10_R0_C06_rom_inst (.q(O8_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clock  (clk));
logic [12-1:0] O8_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_pw_O8_I12_R0_C04_rom_inst (.q(O8_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O8_I12_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O8_I12_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O8_I12_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_pw_O8_I12_R0_C04_rom_inst (.q(O8_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [10-1:0] O8_I14_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O8_I14_R0_C01_rom_inst (.q(O8_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clk(clk),.d(0),.we(0));
//assign O8_I14_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O8_I14_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O8_I14_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O8_I14_R0_C01_rom_inst (.q(O8_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clock  (clk));
logic [11-1:0] O8_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O8_I15_R0_C02_rom_inst (.q(O8_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O8_I15_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O8_I15_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O8_I15_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O8_I15_R0_C02_rom_inst (.q(O8_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [10-1:0] O9_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O9_I1_R0_C01_rom_inst (.q(O9_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O9_I1_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O9_I1_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O9_I1_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O9_I1_R0_C01_rom_inst (.q(O9_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [10-1:0] O9_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O9_I2_R0_C01_rom_inst (.q(O9_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O9_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O9_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O9_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O9_I2_R0_C01_rom_inst (.q(O9_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [11-1:0] O9_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O9_I3_R0_C03_rom_inst (.q(O9_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O9_I3_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O9_I3_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O9_I3_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O9_I3_R0_C03_rom_inst (.q(O9_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [10-1:0] O9_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O9_I6_R0_C01_rom_inst (.q(O9_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O9_I6_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O9_I6_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O9_I6_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O9_I6_R0_C01_rom_inst (.q(O9_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [10-1:0] O9_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O9_I8_R0_C01_rom_inst (.q(O9_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O9_I8_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O9_I8_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O9_I8_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O9_I8_R0_C01_rom_inst (.q(O9_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [10-1:0] O9_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O9_I11_R0_C01_rom_inst (.q(O9_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O9_I11_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O9_I11_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O9_I11_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O9_I11_R0_C01_rom_inst (.q(O9_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [10-1:0] O9_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O9_I13_R0_C01_rom_inst (.q(O9_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O9_I13_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O9_I13_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O9_I13_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O9_I13_R0_C01_rom_inst (.q(O9_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [10-1:0] O9_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O9_I15_R0_C01_rom_inst (.q(O9_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O9_I15_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O9_I15_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O9_I15_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O9_I15_R0_C01_rom_inst (.q(O9_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [11-1:0] O10_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O10_I0_R0_C02_rom_inst (.q(O10_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O10_I0_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O10_I0_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O10_I0_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O10_I0_R0_C02_rom_inst (.q(O10_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [11-1:0] O10_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O10_I1_R0_C03_rom_inst (.q(O10_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O10_I1_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O10_I1_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O10_I1_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O10_I1_R0_C03_rom_inst (.q(O10_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [10-1:0] O10_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O10_I2_R0_C01_rom_inst (.q(O10_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O10_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O10_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O10_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O10_I2_R0_C01_rom_inst (.q(O10_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [10-1:0] O10_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O10_I3_R0_C01_rom_inst (.q(O10_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O10_I3_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O10_I3_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O10_I3_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O10_I3_R0_C01_rom_inst (.q(O10_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [12-1:0] O10_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_pw_O10_I5_R0_C06_rom_inst (.q(O10_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O10_I5_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O10_I5_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O10_I5_R0_C06_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_pw_O10_I5_R0_C06_rom_inst (.q(O10_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [12-1:0] O10_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_pw_O10_I7_R0_C04_rom_inst (.q(O10_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O10_I7_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O10_I7_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O10_I7_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_pw_O10_I7_R0_C04_rom_inst (.q(O10_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [11-1:0] O10_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O10_I8_R0_C02_rom_inst (.q(O10_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O10_I8_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O10_I8_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O10_I8_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O10_I8_R0_C02_rom_inst (.q(O10_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [12-1:0] O10_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_pw_O10_I9_R0_C05_rom_inst (.q(O10_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O10_I9_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O10_I9_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O10_I9_R0_C05_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_pw_O10_I9_R0_C05_rom_inst (.q(O10_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [11-1:0] O10_I10_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O10_I10_R0_C03_rom_inst (.q(O10_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clk(clk),.d(0),.we(0));
//assign O10_I10_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O10_I10_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O10_I10_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O10_I10_R0_C03_rom_inst (.q(O10_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clock  (clk));
logic [10-1:0] O10_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O10_I11_R0_C01_rom_inst (.q(O10_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O10_I11_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O10_I11_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O10_I11_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O10_I11_R0_C01_rom_inst (.q(O10_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [12-1:0] O10_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_pw_O10_I12_R0_C05_rom_inst (.q(O10_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O10_I12_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O10_I12_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O10_I12_R0_C05_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_pw_O10_I12_R0_C05_rom_inst (.q(O10_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [10-1:0] O10_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O10_I15_R0_C01_rom_inst (.q(O10_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O10_I15_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O10_I15_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O10_I15_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O10_I15_R0_C01_rom_inst (.q(O10_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [10-1:0] O11_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O11_I1_R0_C01_rom_inst (.q(O11_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I1_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O11_I1_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O11_I1_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O11_I1_R0_C01_rom_inst (.q(O11_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [10-1:0] O11_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O11_I3_R0_C01_rom_inst (.q(O11_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I3_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O11_I3_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O11_I3_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O11_I3_R0_C01_rom_inst (.q(O11_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [10-1:0] O11_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O11_I4_R0_C01_rom_inst (.q(O11_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I4_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O11_I4_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O11_I4_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O11_I4_R0_C01_rom_inst (.q(O11_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [10-1:0] O11_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O11_I5_R0_C01_rom_inst (.q(O11_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I5_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O11_I5_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O11_I5_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O11_I5_R0_C01_rom_inst (.q(O11_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [10-1:0] O11_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O11_I7_R0_C01_rom_inst (.q(O11_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I7_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O11_I7_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O11_I7_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O11_I7_R0_C01_rom_inst (.q(O11_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [10-1:0] O11_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O11_I8_R0_C01_rom_inst (.q(O11_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I8_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O11_I8_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O11_I8_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O11_I8_R0_C01_rom_inst (.q(O11_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [10-1:0] O11_I10_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O11_I10_R0_C01_rom_inst (.q(O11_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I10_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O11_I10_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O11_I10_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O11_I10_R0_C01_rom_inst (.q(O11_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clock  (clk));
logic [10-1:0] O11_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O11_I11_R0_C01_rom_inst (.q(O11_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I11_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O11_I11_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O11_I11_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O11_I11_R0_C01_rom_inst (.q(O11_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [10-1:0] O11_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O11_I12_R0_C01_rom_inst (.q(O11_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I12_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O11_I12_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O11_I12_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O11_I12_R0_C01_rom_inst (.q(O11_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [11-1:0] O11_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O11_I13_R0_C02_rom_inst (.q(O11_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I13_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O11_I13_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O11_I13_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O11_I13_R0_C02_rom_inst (.q(O11_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [12-1:0] O11_I14_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_pw_O11_I14_R0_C06_rom_inst (.q(O11_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I14_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O11_I14_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O11_I14_R0_C06_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_pw_O11_I14_R0_C06_rom_inst (.q(O11_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clock  (clk));
logic [10-1:0] O12_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O12_I1_R0_C01_rom_inst (.q(O12_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I1_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O12_I1_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O12_I1_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O12_I1_R0_C01_rom_inst (.q(O12_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [10-1:0] O12_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O12_I2_R0_C01_rom_inst (.q(O12_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O12_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O12_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O12_I2_R0_C01_rom_inst (.q(O12_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [10-1:0] O12_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O12_I5_R0_C01_rom_inst (.q(O12_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I5_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O12_I5_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O12_I5_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O12_I5_R0_C01_rom_inst (.q(O12_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [12-1:0] O12_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_pw_O12_I6_R0_C05_rom_inst (.q(O12_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I6_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O12_I6_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O12_I6_R0_C05_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_pw_O12_I6_R0_C05_rom_inst (.q(O12_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [10-1:0] O12_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O12_I8_R0_C01_rom_inst (.q(O12_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I8_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O12_I8_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O12_I8_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O12_I8_R0_C01_rom_inst (.q(O12_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [10-1:0] O12_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O12_I12_R0_C01_rom_inst (.q(O12_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I12_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O12_I12_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O12_I12_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O12_I12_R0_C01_rom_inst (.q(O12_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [10-1:0] O12_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O12_I13_R0_C01_rom_inst (.q(O12_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I13_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O12_I13_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O12_I13_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O12_I13_R0_C01_rom_inst (.q(O12_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [11-1:0] O13_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O13_I0_R0_C02_rom_inst (.q(O13_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O13_I0_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O13_I0_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O13_I0_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O13_I0_R0_C02_rom_inst (.q(O13_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [10-1:0] O13_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O13_I2_R0_C01_rom_inst (.q(O13_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O13_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O13_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O13_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O13_I2_R0_C01_rom_inst (.q(O13_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [11-1:0] O13_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O13_I5_R0_C02_rom_inst (.q(O13_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O13_I5_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O13_I5_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O13_I5_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O13_I5_R0_C02_rom_inst (.q(O13_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [10-1:0] O13_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O13_I12_R0_C01_rom_inst (.q(O13_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O13_I12_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O13_I12_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O13_I12_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O13_I12_R0_C01_rom_inst (.q(O13_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [10-1:0] O13_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O13_I15_R0_C01_rom_inst (.q(O13_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O13_I15_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O13_I15_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O13_I15_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O13_I15_R0_C01_rom_inst (.q(O13_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [11-1:0] O14_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O14_I0_R0_C02_rom_inst (.q(O14_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I0_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O14_I0_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O14_I0_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O14_I0_R0_C02_rom_inst (.q(O14_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [11-1:0] O14_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O14_I5_R0_C03_rom_inst (.q(O14_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I5_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O14_I5_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O14_I5_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O14_I5_R0_C03_rom_inst (.q(O14_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [12-1:0] O14_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_pw_O14_I7_R0_C05_rom_inst (.q(O14_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I7_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O14_I7_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O14_I7_R0_C05_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_pw_O14_I7_R0_C05_rom_inst (.q(O14_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [12-1:0] O14_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_pw_O14_I9_R0_C04_rom_inst (.q(O14_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I9_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O14_I9_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O14_I9_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_pw_O14_I9_R0_C04_rom_inst (.q(O14_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [10-1:0] O14_I10_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O14_I10_R0_C01_rom_inst (.q(O14_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I10_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O14_I10_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O14_I10_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O14_I10_R0_C01_rom_inst (.q(O14_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clock  (clk));
logic [10-1:0] O14_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O14_I11_R0_C01_rom_inst (.q(O14_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I11_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O14_I11_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O14_I11_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O14_I11_R0_C01_rom_inst (.q(O14_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [12-1:0] O14_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_pw_O14_I12_R0_C04_rom_inst (.q(O14_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I12_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O14_I12_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O14_I12_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_pw_O14_I12_R0_C04_rom_inst (.q(O14_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [10-1:0] O14_I14_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O14_I14_R0_C01_rom_inst (.q(O14_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I14_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O14_I14_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O14_I14_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O14_I14_R0_C01_rom_inst (.q(O14_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clock  (clk));
logic [10-1:0] O15_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O15_I0_R0_C01_rom_inst (.q(O15_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I0_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O15_I0_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O15_I0_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O15_I0_R0_C01_rom_inst (.q(O15_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [10-1:0] O15_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O15_I1_R0_C01_rom_inst (.q(O15_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I1_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O15_I1_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O15_I1_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O15_I1_R0_C01_rom_inst (.q(O15_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [10-1:0] O15_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O15_I4_R0_C01_rom_inst (.q(O15_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I4_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O15_I4_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O15_I4_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O15_I4_R0_C01_rom_inst (.q(O15_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [10-1:0] O15_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O15_I6_R0_C01_rom_inst (.q(O15_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I6_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O15_I6_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O15_I6_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O15_I6_R0_C01_rom_inst (.q(O15_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [12-1:0] O15_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_pw_O15_I7_R0_C04_rom_inst (.q(O15_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I7_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O15_I7_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O15_I7_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_pw_O15_I7_R0_C04_rom_inst (.q(O15_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [10-1:0] O15_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O15_I9_R0_C01_rom_inst (.q(O15_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I9_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O15_I9_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O15_I9_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O15_I9_R0_C01_rom_inst (.q(O15_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [10-1:0] O15_I10_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O15_I10_R0_C01_rom_inst (.q(O15_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I10_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O15_I10_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O15_I10_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O15_I10_R0_C01_rom_inst (.q(O15_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clock  (clk));
logic [10-1:0] O15_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O15_I11_R0_C01_rom_inst (.q(O15_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I11_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O15_I11_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O15_I11_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O15_I11_R0_C01_rom_inst (.q(O15_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [10-1:0] O15_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O15_I12_R0_C01_rom_inst (.q(O15_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I12_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O15_I12_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O15_I12_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O15_I12_R0_C01_rom_inst (.q(O15_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [10-1:0] O15_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O15_I15_R0_C01_rom_inst (.q(O15_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I15_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O15_I15_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O15_I15_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O15_I15_R0_C01_rom_inst (.q(O15_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [10-1:0] O16_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O16_I1_R0_C01_rom_inst (.q(O16_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O16_I1_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O16_I1_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O16_I1_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O16_I1_R0_C01_rom_inst (.q(O16_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [10-1:0] O16_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O16_I4_R0_C01_rom_inst (.q(O16_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O16_I4_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O16_I4_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O16_I4_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O16_I4_R0_C01_rom_inst (.q(O16_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [10-1:0] O16_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O16_I8_R0_C01_rom_inst (.q(O16_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O16_I8_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O16_I8_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O16_I8_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O16_I8_R0_C01_rom_inst (.q(O16_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [11-1:0] O16_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O16_I11_R0_C02_rom_inst (.q(O16_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O16_I11_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O16_I11_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O16_I11_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O16_I11_R0_C02_rom_inst (.q(O16_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [11-1:0] O16_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O16_I13_R0_C03_rom_inst (.q(O16_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O16_I13_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O16_I13_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O16_I13_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O16_I13_R0_C03_rom_inst (.q(O16_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [11-1:0] O16_I14_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O16_I14_R0_C03_rom_inst (.q(O16_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clk(clk),.d(0),.we(0));
//assign O16_I14_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O16_I14_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O16_I14_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O16_I14_R0_C03_rom_inst (.q(O16_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clock  (clk));
logic [10-1:0] O17_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O17_I0_R0_C01_rom_inst (.q(O17_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O17_I0_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O17_I0_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O17_I0_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O17_I0_R0_C01_rom_inst (.q(O17_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [12-1:0] O17_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_pw_O17_I2_R0_C04_rom_inst (.q(O17_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O17_I2_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O17_I2_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O17_I2_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_pw_O17_I2_R0_C04_rom_inst (.q(O17_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [11-1:0] O17_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O17_I4_R0_C02_rom_inst (.q(O17_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O17_I4_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O17_I4_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O17_I4_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O17_I4_R0_C02_rom_inst (.q(O17_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [10-1:0] O17_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O17_I5_R0_C01_rom_inst (.q(O17_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O17_I5_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O17_I5_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O17_I5_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O17_I5_R0_C01_rom_inst (.q(O17_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [10-1:0] O17_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O17_I6_R0_C01_rom_inst (.q(O17_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O17_I6_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O17_I6_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O17_I6_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O17_I6_R0_C01_rom_inst (.q(O17_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [10-1:0] O17_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O17_I9_R0_C01_rom_inst (.q(O17_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O17_I9_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O17_I9_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O17_I9_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O17_I9_R0_C01_rom_inst (.q(O17_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [10-1:0] O17_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O17_I11_R0_C01_rom_inst (.q(O17_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O17_I11_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O17_I11_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O17_I11_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O17_I11_R0_C01_rom_inst (.q(O17_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [10-1:0] O17_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O17_I12_R0_C01_rom_inst (.q(O17_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O17_I12_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O17_I12_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O17_I12_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O17_I12_R0_C01_rom_inst (.q(O17_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [11-1:0] O17_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O17_I15_R0_C02_rom_inst (.q(O17_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O17_I15_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O17_I15_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O17_I15_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O17_I15_R0_C02_rom_inst (.q(O17_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [10-1:0] O18_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O18_I0_R0_C01_rom_inst (.q(O18_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O18_I0_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O18_I0_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O18_I0_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O18_I0_R0_C01_rom_inst (.q(O18_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [11-1:0] O18_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O18_I5_R0_C02_rom_inst (.q(O18_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O18_I5_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O18_I5_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O18_I5_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O18_I5_R0_C02_rom_inst (.q(O18_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [12-1:0] O18_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_pw_O18_I9_R0_C04_rom_inst (.q(O18_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O18_I9_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O18_I9_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O18_I9_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_pw_O18_I9_R0_C04_rom_inst (.q(O18_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [11-1:0] O18_I10_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O18_I10_R0_C02_rom_inst (.q(O18_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clk(clk),.d(0),.we(0));
//assign O18_I10_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O18_I10_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O18_I10_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O18_I10_R0_C02_rom_inst (.q(O18_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clock  (clk));
logic [10-1:0] O19_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O19_I0_R0_C01_rom_inst (.q(O19_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O19_I0_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O19_I0_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O19_I0_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O19_I0_R0_C01_rom_inst (.q(O19_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [10-1:0] O19_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O19_I6_R0_C01_rom_inst (.q(O19_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O19_I6_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O19_I6_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O19_I6_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O19_I6_R0_C01_rom_inst (.q(O19_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [11-1:0] O19_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O19_I11_R0_C03_rom_inst (.q(O19_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O19_I11_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O19_I11_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O19_I11_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O19_I11_R0_C03_rom_inst (.q(O19_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [10-1:0] O19_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O19_I13_R0_C01_rom_inst (.q(O19_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O19_I13_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O19_I13_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O19_I13_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O19_I13_R0_C01_rom_inst (.q(O19_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [11-1:0] O20_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O20_I11_R0_C02_rom_inst (.q(O20_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O20_I11_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O20_I11_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O20_I11_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O20_I11_R0_C02_rom_inst (.q(O20_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [10-1:0] O20_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O20_I13_R0_C01_rom_inst (.q(O20_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O20_I13_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O20_I13_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O20_I13_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O20_I13_R0_C01_rom_inst (.q(O20_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [12-1:0] O21_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_pw_O21_I2_R0_C04_rom_inst (.q(O21_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O21_I2_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O21_I2_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O21_I2_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_pw_O21_I2_R0_C04_rom_inst (.q(O21_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [10-1:0] O21_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O21_I3_R0_C01_rom_inst (.q(O21_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O21_I3_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O21_I3_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O21_I3_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O21_I3_R0_C01_rom_inst (.q(O21_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [11-1:0] O21_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O21_I5_R0_C02_rom_inst (.q(O21_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O21_I5_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O21_I5_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O21_I5_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O21_I5_R0_C02_rom_inst (.q(O21_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [10-1:0] O21_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O21_I6_R0_C01_rom_inst (.q(O21_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O21_I6_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O21_I6_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O21_I6_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O21_I6_R0_C01_rom_inst (.q(O21_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [12-1:0] O21_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_pw_O21_I7_R0_C05_rom_inst (.q(O21_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O21_I7_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O21_I7_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O21_I7_R0_C05_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_pw_O21_I7_R0_C05_rom_inst (.q(O21_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [10-1:0] O21_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O21_I8_R0_C01_rom_inst (.q(O21_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O21_I8_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O21_I8_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O21_I8_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O21_I8_R0_C01_rom_inst (.q(O21_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [11-1:0] O21_I10_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O21_I10_R0_C03_rom_inst (.q(O21_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clk(clk),.d(0),.we(0));
//assign O21_I10_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O21_I10_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O21_I10_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O21_I10_R0_C03_rom_inst (.q(O21_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clock  (clk));
logic [10-1:0] O21_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O21_I11_R0_C01_rom_inst (.q(O21_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O21_I11_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O21_I11_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O21_I11_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O21_I11_R0_C01_rom_inst (.q(O21_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [10-1:0] O21_I14_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O21_I14_R0_C01_rom_inst (.q(O21_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clk(clk),.d(0),.we(0));
//assign O21_I14_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O21_I14_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O21_I14_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O21_I14_R0_C01_rom_inst (.q(O21_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clock  (clk));
logic [10-1:0] O21_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O21_I15_R0_C01_rom_inst (.q(O21_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O21_I15_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O21_I15_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O21_I15_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O21_I15_R0_C01_rom_inst (.q(O21_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [11-1:0] O22_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O22_I0_R0_C03_rom_inst (.q(O22_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O22_I0_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O22_I0_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O22_I0_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O22_I0_R0_C03_rom_inst (.q(O22_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [10-1:0] O22_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O22_I2_R0_C01_rom_inst (.q(O22_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O22_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O22_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O22_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O22_I2_R0_C01_rom_inst (.q(O22_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [11-1:0] O22_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O22_I5_R0_C02_rom_inst (.q(O22_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O22_I5_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O22_I5_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O22_I5_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O22_I5_R0_C02_rom_inst (.q(O22_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [10-1:0] O22_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O22_I8_R0_C01_rom_inst (.q(O22_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O22_I8_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O22_I8_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O22_I8_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O22_I8_R0_C01_rom_inst (.q(O22_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [10-1:0] O22_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O22_I9_R0_C01_rom_inst (.q(O22_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O22_I9_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O22_I9_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O22_I9_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O22_I9_R0_C01_rom_inst (.q(O22_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [10-1:0] O22_I10_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O22_I10_R0_C01_rom_inst (.q(O22_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clk(clk),.d(0),.we(0));
//assign O22_I10_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O22_I10_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O22_I10_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O22_I10_R0_C01_rom_inst (.q(O22_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clock  (clk));
logic [10-1:0] O22_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O22_I11_R0_C01_rom_inst (.q(O22_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O22_I11_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O22_I11_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O22_I11_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O22_I11_R0_C01_rom_inst (.q(O22_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [10-1:0] O22_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O22_I12_R0_C01_rom_inst (.q(O22_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O22_I12_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O22_I12_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O22_I12_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O22_I12_R0_C01_rom_inst (.q(O22_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [11-1:0] O22_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O22_I15_R0_C03_rom_inst (.q(O22_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O22_I15_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O22_I15_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O22_I15_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O22_I15_R0_C03_rom_inst (.q(O22_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [10-1:0] O23_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O23_I1_R0_C01_rom_inst (.q(O23_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O23_I1_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O23_I1_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O23_I1_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O23_I1_R0_C01_rom_inst (.q(O23_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [12-1:0] O23_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_pw_O23_I3_R0_C05_rom_inst (.q(O23_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O23_I3_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O23_I3_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O23_I3_R0_C05_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_pw_O23_I3_R0_C05_rom_inst (.q(O23_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [12-1:0] O23_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_pw_O23_I4_R0_C04_rom_inst (.q(O23_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O23_I4_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O23_I4_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O23_I4_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_pw_O23_I4_R0_C04_rom_inst (.q(O23_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [10-1:0] O23_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O23_I5_R0_C01_rom_inst (.q(O23_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O23_I5_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O23_I5_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O23_I5_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O23_I5_R0_C01_rom_inst (.q(O23_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [12-1:0] O23_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_pw_O23_I8_R0_C05_rom_inst (.q(O23_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O23_I8_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O23_I8_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O23_I8_R0_C05_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_pw_O23_I8_R0_C05_rom_inst (.q(O23_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [10-1:0] O23_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O23_I11_R0_C01_rom_inst (.q(O23_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O23_I11_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O23_I11_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O23_I11_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O23_I11_R0_C01_rom_inst (.q(O23_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [10-1:0] O23_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O23_I12_R0_C01_rom_inst (.q(O23_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O23_I12_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O23_I12_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O23_I12_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O23_I12_R0_C01_rom_inst (.q(O23_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [10-1:0] O23_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O23_I13_R0_C01_rom_inst (.q(O23_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O23_I13_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O23_I13_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O23_I13_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O23_I13_R0_C01_rom_inst (.q(O23_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [10-1:0] O23_I14_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O23_I14_R0_C01_rom_inst (.q(O23_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clk(clk),.d(0),.we(0));
//assign O23_I14_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O23_I14_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O23_I14_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O23_I14_R0_C01_rom_inst (.q(O23_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clock  (clk));
logic [11-1:0] O24_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O24_I0_R0_C03_rom_inst (.q(O24_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O24_I0_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O24_I0_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O24_I0_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O24_I0_R0_C03_rom_inst (.q(O24_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [11-1:0] O24_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O24_I1_R0_C02_rom_inst (.q(O24_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O24_I1_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O24_I1_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O24_I1_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O24_I1_R0_C02_rom_inst (.q(O24_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [10-1:0] O24_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O24_I2_R0_C01_rom_inst (.q(O24_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O24_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O24_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O24_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O24_I2_R0_C01_rom_inst (.q(O24_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [12-1:0] O24_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_pw_O24_I3_R0_C06_rom_inst (.q(O24_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O24_I3_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O24_I3_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O24_I3_R0_C06_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_pw_O24_I3_R0_C06_rom_inst (.q(O24_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [12-1:0] O24_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_pw_O24_I4_R0_C04_rom_inst (.q(O24_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O24_I4_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O24_I4_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O24_I4_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_pw_O24_I4_R0_C04_rom_inst (.q(O24_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [10-1:0] O24_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O24_I5_R0_C01_rom_inst (.q(O24_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O24_I5_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O24_I5_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O24_I5_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O24_I5_R0_C01_rom_inst (.q(O24_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [11-1:0] O24_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O24_I6_R0_C02_rom_inst (.q(O24_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O24_I6_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O24_I6_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O24_I6_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O24_I6_R0_C02_rom_inst (.q(O24_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [11-1:0] O24_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O24_I7_R0_C03_rom_inst (.q(O24_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O24_I7_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O24_I7_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O24_I7_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O24_I7_R0_C03_rom_inst (.q(O24_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [13-1:0] O24_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv4_pw_O24_I8_R0_C09_rom_inst (.q(O24_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O24_I8_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O24_I8_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O24_I8_R0_C09_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv4_pw_O24_I8_R0_C09_rom_inst (.q(O24_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [10-1:0] O24_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O24_I9_R0_C01_rom_inst (.q(O24_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O24_I9_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O24_I9_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O24_I9_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O24_I9_R0_C01_rom_inst (.q(O24_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [11-1:0] O24_I10_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O24_I10_R0_C02_rom_inst (.q(O24_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clk(clk),.d(0),.we(0));
//assign O24_I10_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O24_I10_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O24_I10_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O24_I10_R0_C02_rom_inst (.q(O24_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clock  (clk));
logic [12-1:0] O24_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_pw_O24_I11_R0_C04_rom_inst (.q(O24_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O24_I11_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O24_I11_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O24_I11_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_pw_O24_I11_R0_C04_rom_inst (.q(O24_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [12-1:0] O24_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_pw_O24_I13_R0_C04_rom_inst (.q(O24_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O24_I13_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O24_I13_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O24_I13_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_pw_O24_I13_R0_C04_rom_inst (.q(O24_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [11-1:0] O24_I14_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O24_I14_R0_C03_rom_inst (.q(O24_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clk(clk),.d(0),.we(0));
//assign O24_I14_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O24_I14_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O24_I14_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O24_I14_R0_C03_rom_inst (.q(O24_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clock  (clk));
logic [10-1:0] O24_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O24_I15_R0_C01_rom_inst (.q(O24_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O24_I15_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O24_I15_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O24_I15_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O24_I15_R0_C01_rom_inst (.q(O24_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [11-1:0] O25_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O25_I1_R0_C02_rom_inst (.q(O25_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O25_I1_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O25_I1_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O25_I1_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O25_I1_R0_C02_rom_inst (.q(O25_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [10-1:0] O25_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O25_I3_R0_C01_rom_inst (.q(O25_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O25_I3_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O25_I3_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O25_I3_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O25_I3_R0_C01_rom_inst (.q(O25_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [10-1:0] O25_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O25_I5_R0_C01_rom_inst (.q(O25_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O25_I5_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O25_I5_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O25_I5_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O25_I5_R0_C01_rom_inst (.q(O25_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [10-1:0] O25_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O25_I6_R0_C01_rom_inst (.q(O25_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O25_I6_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O25_I6_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O25_I6_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O25_I6_R0_C01_rom_inst (.q(O25_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [10-1:0] O25_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O25_I7_R0_C01_rom_inst (.q(O25_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O25_I7_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O25_I7_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O25_I7_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O25_I7_R0_C01_rom_inst (.q(O25_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [10-1:0] O25_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O25_I8_R0_C01_rom_inst (.q(O25_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O25_I8_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O25_I8_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O25_I8_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O25_I8_R0_C01_rom_inst (.q(O25_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [10-1:0] O25_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O25_I9_R0_C01_rom_inst (.q(O25_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O25_I9_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O25_I9_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O25_I9_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O25_I9_R0_C01_rom_inst (.q(O25_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [10-1:0] O25_I10_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O25_I10_R0_C01_rom_inst (.q(O25_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clk(clk),.d(0),.we(0));
//assign O25_I10_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O25_I10_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O25_I10_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O25_I10_R0_C01_rom_inst (.q(O25_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clock  (clk));
logic [11-1:0] O25_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O25_I11_R0_C02_rom_inst (.q(O25_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O25_I11_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O25_I11_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O25_I11_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O25_I11_R0_C02_rom_inst (.q(O25_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [10-1:0] O25_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O25_I12_R0_C01_rom_inst (.q(O25_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O25_I12_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O25_I12_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O25_I12_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O25_I12_R0_C01_rom_inst (.q(O25_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [10-1:0] O25_I14_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O25_I14_R0_C01_rom_inst (.q(O25_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clk(clk),.d(0),.we(0));
//assign O25_I14_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O25_I14_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O25_I14_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O25_I14_R0_C01_rom_inst (.q(O25_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clock  (clk));
logic [10-1:0] O26_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O26_I1_R0_C01_rom_inst (.q(O26_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O26_I1_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O26_I1_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O26_I1_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O26_I1_R0_C01_rom_inst (.q(O26_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [10-1:0] O26_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O26_I2_R0_C01_rom_inst (.q(O26_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O26_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O26_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O26_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O26_I2_R0_C01_rom_inst (.q(O26_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [10-1:0] O26_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O26_I3_R0_C01_rom_inst (.q(O26_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O26_I3_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O26_I3_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O26_I3_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O26_I3_R0_C01_rom_inst (.q(O26_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [11-1:0] O26_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O26_I4_R0_C02_rom_inst (.q(O26_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O26_I4_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O26_I4_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O26_I4_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O26_I4_R0_C02_rom_inst (.q(O26_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [10-1:0] O26_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O26_I6_R0_C01_rom_inst (.q(O26_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O26_I6_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O26_I6_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O26_I6_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O26_I6_R0_C01_rom_inst (.q(O26_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [10-1:0] O26_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O26_I8_R0_C01_rom_inst (.q(O26_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O26_I8_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O26_I8_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O26_I8_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O26_I8_R0_C01_rom_inst (.q(O26_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [10-1:0] O26_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O26_I11_R0_C01_rom_inst (.q(O26_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O26_I11_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O26_I11_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O26_I11_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O26_I11_R0_C01_rom_inst (.q(O26_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [11-1:0] O26_I14_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O26_I14_R0_C02_rom_inst (.q(O26_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clk(clk),.d(0),.we(0));
//assign O26_I14_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O26_I14_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O26_I14_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O26_I14_R0_C02_rom_inst (.q(O26_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clock  (clk));
logic [11-1:0] O27_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O27_I0_R0_C02_rom_inst (.q(O27_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O27_I0_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O27_I0_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O27_I0_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O27_I0_R0_C02_rom_inst (.q(O27_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [11-1:0] O27_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O27_I5_R0_C02_rom_inst (.q(O27_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O27_I5_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O27_I5_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O27_I5_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O27_I5_R0_C02_rom_inst (.q(O27_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [11-1:0] O27_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O27_I12_R0_C02_rom_inst (.q(O27_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O27_I12_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O27_I12_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O27_I12_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O27_I12_R0_C02_rom_inst (.q(O27_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [11-1:0] O27_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O27_I15_R0_C02_rom_inst (.q(O27_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O27_I15_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O27_I15_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O27_I15_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O27_I15_R0_C02_rom_inst (.q(O27_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [11-1:0] O28_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O28_I0_R0_C02_rom_inst (.q(O28_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O28_I0_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O28_I0_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O28_I0_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O28_I0_R0_C02_rom_inst (.q(O28_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [10-1:0] O28_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O28_I1_R0_C01_rom_inst (.q(O28_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O28_I1_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O28_I1_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O28_I1_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O28_I1_R0_C01_rom_inst (.q(O28_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [10-1:0] O28_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O28_I3_R0_C01_rom_inst (.q(O28_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O28_I3_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O28_I3_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O28_I3_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O28_I3_R0_C01_rom_inst (.q(O28_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [11-1:0] O28_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O28_I4_R0_C02_rom_inst (.q(O28_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O28_I4_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O28_I4_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O28_I4_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O28_I4_R0_C02_rom_inst (.q(O28_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [11-1:0] O28_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O28_I5_R0_C02_rom_inst (.q(O28_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O28_I5_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O28_I5_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O28_I5_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O28_I5_R0_C02_rom_inst (.q(O28_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [11-1:0] O28_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O28_I6_R0_C02_rom_inst (.q(O28_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O28_I6_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O28_I6_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O28_I6_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O28_I6_R0_C02_rom_inst (.q(O28_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [11-1:0] O28_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O28_I7_R0_C02_rom_inst (.q(O28_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O28_I7_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O28_I7_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O28_I7_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O28_I7_R0_C02_rom_inst (.q(O28_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [11-1:0] O28_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O28_I8_R0_C02_rom_inst (.q(O28_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O28_I8_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O28_I8_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O28_I8_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O28_I8_R0_C02_rom_inst (.q(O28_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [10-1:0] O28_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O28_I9_R0_C01_rom_inst (.q(O28_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O28_I9_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O28_I9_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O28_I9_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O28_I9_R0_C01_rom_inst (.q(O28_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [10-1:0] O28_I10_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O28_I10_R0_C01_rom_inst (.q(O28_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clk(clk),.d(0),.we(0));
//assign O28_I10_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O28_I10_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O28_I10_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O28_I10_R0_C01_rom_inst (.q(O28_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clock  (clk));
logic [10-1:0] O28_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O28_I12_R0_C01_rom_inst (.q(O28_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O28_I12_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O28_I12_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O28_I12_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O28_I12_R0_C01_rom_inst (.q(O28_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [11-1:0] O28_I14_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O28_I14_R0_C02_rom_inst (.q(O28_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clk(clk),.d(0),.we(0));
//assign O28_I14_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O28_I14_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O28_I14_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O28_I14_R0_C02_rom_inst (.q(O28_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clock  (clk));
logic [10-1:0] O28_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O28_I15_R0_C01_rom_inst (.q(O28_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O28_I15_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O28_I15_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O28_I15_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O28_I15_R0_C01_rom_inst (.q(O28_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [11-1:0] O29_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O29_I0_R0_C02_rom_inst (.q(O29_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O29_I0_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O29_I0_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O29_I0_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O29_I0_R0_C02_rom_inst (.q(O29_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [10-1:0] O29_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O29_I1_R0_C01_rom_inst (.q(O29_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O29_I1_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O29_I1_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O29_I1_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O29_I1_R0_C01_rom_inst (.q(O29_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [12-1:0] O29_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_pw_O29_I5_R0_C05_rom_inst (.q(O29_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O29_I5_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O29_I5_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O29_I5_R0_C05_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_pw_O29_I5_R0_C05_rom_inst (.q(O29_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [10-1:0] O29_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O29_I7_R0_C01_rom_inst (.q(O29_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O29_I7_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O29_I7_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O29_I7_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O29_I7_R0_C01_rom_inst (.q(O29_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [10-1:0] O29_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O29_I9_R0_C01_rom_inst (.q(O29_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O29_I9_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O29_I9_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O29_I9_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O29_I9_R0_C01_rom_inst (.q(O29_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [12-1:0] O29_I10_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_pw_O29_I10_R0_C04_rom_inst (.q(O29_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clk(clk),.d(0),.we(0));
//assign O29_I10_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O29_I10_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O29_I10_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_pw_O29_I10_R0_C04_rom_inst (.q(O29_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clock  (clk));
logic [12-1:0] O29_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_pw_O29_I12_R0_C06_rom_inst (.q(O29_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O29_I12_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O29_I12_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O29_I12_R0_C06_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_pw_O29_I12_R0_C06_rom_inst (.q(O29_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [10-1:0] O29_I14_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O29_I14_R0_C01_rom_inst (.q(O29_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clk(clk),.d(0),.we(0));
//assign O29_I14_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O29_I14_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O29_I14_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O29_I14_R0_C01_rom_inst (.q(O29_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clock  (clk));
logic [11-1:0] O29_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O29_I15_R0_C02_rom_inst (.q(O29_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O29_I15_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O29_I15_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O29_I15_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O29_I15_R0_C02_rom_inst (.q(O29_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [10-1:0] O30_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O30_I0_R0_C01_rom_inst (.q(O30_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O30_I0_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O30_I0_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O30_I0_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O30_I0_R0_C01_rom_inst (.q(O30_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [10-1:0] O30_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O30_I1_R0_C01_rom_inst (.q(O30_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O30_I1_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O30_I1_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O30_I1_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O30_I1_R0_C01_rom_inst (.q(O30_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [11-1:0] O30_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O30_I2_R0_C02_rom_inst (.q(O30_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O30_I2_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O30_I2_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O30_I2_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O30_I2_R0_C02_rom_inst (.q(O30_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [11-1:0] O30_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O30_I3_R0_C02_rom_inst (.q(O30_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O30_I3_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O30_I3_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O30_I3_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O30_I3_R0_C02_rom_inst (.q(O30_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [10-1:0] O30_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O30_I6_R0_C01_rom_inst (.q(O30_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O30_I6_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O30_I6_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O30_I6_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O30_I6_R0_C01_rom_inst (.q(O30_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [10-1:0] O30_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O30_I8_R0_C01_rom_inst (.q(O30_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O30_I8_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O30_I8_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O30_I8_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O30_I8_R0_C01_rom_inst (.q(O30_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [10-1:0] O30_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O30_I11_R0_C01_rom_inst (.q(O30_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O30_I11_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O30_I11_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O30_I11_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O30_I11_R0_C01_rom_inst (.q(O30_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [10-1:0] O30_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O30_I12_R0_C01_rom_inst (.q(O30_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O30_I12_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O30_I12_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O30_I12_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O30_I12_R0_C01_rom_inst (.q(O30_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [10-1:0] O30_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O30_I13_R0_C01_rom_inst (.q(O30_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O30_I13_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O30_I13_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O30_I13_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O30_I13_R0_C01_rom_inst (.q(O30_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [12-1:0] O30_I14_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv4_pw_O30_I14_R0_C05_rom_inst (.q(O30_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clk(clk),.d(0),.we(0));
//assign O30_I14_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O30_I14_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O30_I14_R0_C05_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv4_pw_O30_I14_R0_C05_rom_inst (.q(O30_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clock  (clk));
logic [10-1:0] O30_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O30_I15_R0_C01_rom_inst (.q(O30_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O30_I15_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O30_I15_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O30_I15_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O30_I15_R0_C01_rom_inst (.q(O30_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [10-1:0] O31_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O31_I0_R0_C01_rom_inst (.q(O31_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O31_I0_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O31_I0_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O31_I0_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O31_I0_R0_C01_rom_inst (.q(O31_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [10-1:0] O31_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O31_I1_R0_C01_rom_inst (.q(O31_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O31_I1_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O31_I1_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O31_I1_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O31_I1_R0_C01_rom_inst (.q(O31_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [10-1:0] O31_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O31_I2_R0_C01_rom_inst (.q(O31_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O31_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O31_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O31_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O31_I2_R0_C01_rom_inst (.q(O31_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [10-1:0] O31_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O31_I3_R0_C01_rom_inst (.q(O31_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O31_I3_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O31_I3_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O31_I3_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O31_I3_R0_C01_rom_inst (.q(O31_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [11-1:0] O31_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O31_I4_R0_C02_rom_inst (.q(O31_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O31_I4_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O31_I4_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O31_I4_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O31_I4_R0_C02_rom_inst (.q(O31_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [10-1:0] O31_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O31_I8_R0_C01_rom_inst (.q(O31_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O31_I8_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O31_I8_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O31_I8_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O31_I8_R0_C01_rom_inst (.q(O31_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [10-1:0] O31_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O31_I11_R0_C01_rom_inst (.q(O31_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O31_I11_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O31_I11_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O31_I11_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O31_I11_R0_C01_rom_inst (.q(O31_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [10-1:0] O31_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O31_I12_R0_C01_rom_inst (.q(O31_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O31_I12_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O31_I12_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O31_I12_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O31_I12_R0_C01_rom_inst (.q(O31_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [10-1:0] O31_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv4_pw_O31_I13_R0_C01_rom_inst (.q(O31_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O31_I13_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O31_I13_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O31_I13_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv4_pw_O31_I13_R0_C01_rom_inst (.q(O31_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [11-1:0] O31_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv4_pw_O31_I15_R0_C02_rom_inst (.q(O31_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O31_I15_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O31_I15_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv4_pw_O31_I15_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv4_pw_O31_I15_R0_C02_rom_inst (.q(O31_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic signed [31:0] conv_mac_0;
logic signed [31:0] O0_N0_S0;		always @(posedge clk) O0_N0_S0 <=     O0_I0_R0_C0_SM1   +  O0_I2_R0_C0_SM1  ;
 logic signed [31:0] O0_N2_S0;		always @(posedge clk) O0_N2_S0 <=     O0_I5_R0_C0_SM1   +  O0_I15_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O0_N0_S1;		always @(posedge clk) O0_N0_S1 <=     O0_N0_S0  +  O0_N2_S0 ;
 assign conv_mac_0 = O0_N0_S1;

logic signed [31:0] conv_mac_1;
logic signed [31:0] O1_N0_S0;		always @(posedge clk) O1_N0_S0 <=     O1_I0_R0_C0_SM1   +  O1_I1_R0_C0_SM1  ;
 logic signed [31:0] O1_N2_S0;		always @(posedge clk) O1_N2_S0 <=     O1_I2_R0_C0_SM1   +  O1_I5_R0_C0_SM1  ;
 logic signed [31:0] O1_N4_S0;		always @(posedge clk) O1_N4_S0 <=     O1_I6_R0_C0_SM1   +  O1_I7_R0_C0_SM1  ;
 logic signed [31:0] O1_N6_S0;		always @(posedge clk) O1_N6_S0 <=     O1_I8_R0_C0_SM1   +  O1_I9_R0_C0_SM1  ;
 logic signed [31:0] O1_N8_S0;		always @(posedge clk) O1_N8_S0 <=     O1_I14_R0_C0_SM1   +  O1_I15_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O1_N0_S1;		always @(posedge clk) O1_N0_S1 <=     O1_N0_S0  +  O1_N2_S0 ;
 logic signed [31:0] O1_N2_S1;		always @(posedge clk) O1_N2_S1 <=     O1_N4_S0  +  O1_N6_S0 ;
 logic signed [31:0] O1_N4_S1;		always @(posedge clk) O1_N4_S1 <=     O1_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O1_N0_S2;		always @(posedge clk) O1_N0_S2 <=     O1_N0_S1  +  O1_N2_S1 ;
 logic signed [31:0] O1_N2_S2;		always @(posedge clk) O1_N2_S2 <=     O1_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O1_N0_S3;		always @(posedge clk) O1_N0_S3 <=     O1_N0_S2  +  O1_N2_S2 ;
 assign conv_mac_1 = O1_N0_S3;

logic signed [31:0] conv_mac_2;
logic signed [31:0] O2_N0_S0;		always @(posedge clk) O2_N0_S0 <=     O2_I1_R0_C0_SM1   +  O2_I2_R0_C0_SM1  ;
 logic signed [31:0] O2_N2_S0;		always @(posedge clk) O2_N2_S0 <=     O2_I4_R0_C0_SM1   +  O2_I6_R0_C0_SM1  ;
 logic signed [31:0] O2_N4_S0;		always @(posedge clk) O2_N4_S0 <=     O2_I7_R0_C0_SM1   +  O2_I11_R0_C0_SM1  ;
 logic signed [31:0] O2_N6_S0;		always @(posedge clk) O2_N6_S0 <=     O2_I15_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O2_N0_S1;		always @(posedge clk) O2_N0_S1 <=     O2_N0_S0  +  O2_N2_S0 ;
 logic signed [31:0] O2_N2_S1;		always @(posedge clk) O2_N2_S1 <=     O2_N4_S0  +  O2_N6_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O2_N0_S2;		always @(posedge clk) O2_N0_S2 <=     O2_N0_S1  +  O2_N2_S1 ;
 assign conv_mac_2 = O2_N0_S2;

logic signed [31:0] conv_mac_3;
logic signed [31:0] O3_N0_S0;		always @(posedge clk) O3_N0_S0 <=     O3_I0_R0_C0_SM1   +  O3_I2_R0_C0_SM1  ;
 logic signed [31:0] O3_N2_S0;		always @(posedge clk) O3_N2_S0 <=     O3_I4_R0_C0_SM1   +  O3_I5_R0_C0_SM1  ;
 logic signed [31:0] O3_N4_S0;		always @(posedge clk) O3_N4_S0 <=     O3_I6_R0_C0_SM1   +  O3_I7_R0_C0_SM1  ;
 logic signed [31:0] O3_N6_S0;		always @(posedge clk) O3_N6_S0 <=     O3_I8_R0_C0_SM1   +  O3_I9_R0_C0_SM1  ;
 logic signed [31:0] O3_N8_S0;		always @(posedge clk) O3_N8_S0 <=     O3_I10_R0_C0_SM1   +  O3_I12_R0_C0_SM1  ;
 logic signed [31:0] O3_N10_S0;		always @(posedge clk) O3_N10_S0 <=     O3_I14_R0_C0_SM1   +  O3_I15_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O3_N0_S1;		always @(posedge clk) O3_N0_S1 <=     O3_N0_S0  +  O3_N2_S0 ;
 logic signed [31:0] O3_N2_S1;		always @(posedge clk) O3_N2_S1 <=     O3_N4_S0  +  O3_N6_S0 ;
 logic signed [31:0] O3_N4_S1;		always @(posedge clk) O3_N4_S1 <=     O3_N8_S0  +  O3_N10_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O3_N0_S2;		always @(posedge clk) O3_N0_S2 <=     O3_N0_S1  +  O3_N2_S1 ;
 logic signed [31:0] O3_N2_S2;		always @(posedge clk) O3_N2_S2 <=     O3_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O3_N0_S3;		always @(posedge clk) O3_N0_S3 <=     O3_N0_S2  +  O3_N2_S2 ;
 assign conv_mac_3 = O3_N0_S3;

logic signed [31:0] conv_mac_4;
logic signed [31:0] O4_N0_S0;		always @(posedge clk) O4_N0_S0 <=     O4_I0_R0_C0_SM1   +  O4_I1_R0_C0_SM1  ;
 logic signed [31:0] O4_N2_S0;		always @(posedge clk) O4_N2_S0 <=     O4_I3_R0_C0_SM1   +  O4_I4_R0_C0_SM1  ;
 logic signed [31:0] O4_N4_S0;		always @(posedge clk) O4_N4_S0 <=     O4_I5_R0_C0_SM1   +  O4_I7_R0_C0_SM1  ;
 logic signed [31:0] O4_N6_S0;		always @(posedge clk) O4_N6_S0 <=     O4_I8_R0_C0_SM1   +  O4_I9_R0_C0_SM1  ;
 logic signed [31:0] O4_N8_S0;		always @(posedge clk) O4_N8_S0 <=     O4_I11_R0_C0_SM1   +  O4_I12_R0_C0_SM1  ;
 logic signed [31:0] O4_N10_S0;		always @(posedge clk) O4_N10_S0 <=     O4_I13_R0_C0_SM1   +  O4_I14_R0_C0_SM1  ;
 logic signed [31:0] O4_N12_S0;		always @(posedge clk) O4_N12_S0 <=     O4_I15_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O4_N0_S1;		always @(posedge clk) O4_N0_S1 <=     O4_N0_S0  +  O4_N2_S0 ;
 logic signed [31:0] O4_N2_S1;		always @(posedge clk) O4_N2_S1 <=     O4_N4_S0  +  O4_N6_S0 ;
 logic signed [31:0] O4_N4_S1;		always @(posedge clk) O4_N4_S1 <=     O4_N8_S0  +  O4_N10_S0 ;
 logic signed [31:0] O4_N6_S1;		always @(posedge clk) O4_N6_S1 <=     O4_N12_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O4_N0_S2;		always @(posedge clk) O4_N0_S2 <=     O4_N0_S1  +  O4_N2_S1 ;
 logic signed [31:0] O4_N2_S2;		always @(posedge clk) O4_N2_S2 <=     O4_N4_S1  +  O4_N6_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O4_N0_S3;		always @(posedge clk) O4_N0_S3 <=     O4_N0_S2  +  O4_N2_S2 ;
 assign conv_mac_4 = O4_N0_S3;

logic signed [31:0] conv_mac_5;
logic signed [31:0] O5_N0_S0;		always @(posedge clk) O5_N0_S0 <=     O5_I1_R0_C0_SM1   +  O5_I2_R0_C0_SM1  ;
 logic signed [31:0] O5_N2_S0;		always @(posedge clk) O5_N2_S0 <=     O5_I10_R0_C0_SM1   +  O5_I12_R0_C0_SM1  ;
 logic signed [31:0] O5_N4_S0;		always @(posedge clk) O5_N4_S0 <=     O5_I15_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O5_N0_S1;		always @(posedge clk) O5_N0_S1 <=     O5_N0_S0  +  O5_N2_S0 ;
 logic signed [31:0] O5_N2_S1;		always @(posedge clk) O5_N2_S1 <=     O5_N4_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O5_N0_S2;		always @(posedge clk) O5_N0_S2 <=     O5_N0_S1  +  O5_N2_S1 ;
 assign conv_mac_5 = O5_N0_S2;

logic signed [31:0] conv_mac_6;
logic signed [31:0] O6_N0_S0;		always @(posedge clk) O6_N0_S0 <=     O6_I0_R0_C0_SM1   +  O6_I1_R0_C0_SM1  ;
 logic signed [31:0] O6_N2_S0;		always @(posedge clk) O6_N2_S0 <=     O6_I2_R0_C0_SM1   +  O6_I4_R0_C0_SM1  ;
 logic signed [31:0] O6_N4_S0;		always @(posedge clk) O6_N4_S0 <=     O6_I5_R0_C0_SM1   +  O6_I7_R0_C0_SM1  ;
 logic signed [31:0] O6_N6_S0;		always @(posedge clk) O6_N6_S0 <=     O6_I8_R0_C0_SM1   +  O6_I9_R0_C0_SM1  ;
 logic signed [31:0] O6_N8_S0;		always @(posedge clk) O6_N8_S0 <=     O6_I10_R0_C0_SM1   +  O6_I12_R0_C0_SM1  ;
 logic signed [31:0] O6_N10_S0;		always @(posedge clk) O6_N10_S0 <=     O6_I13_R0_C0_SM1   +  O6_I14_R0_C0_SM1  ;
 logic signed [31:0] O6_N12_S0;		always @(posedge clk) O6_N12_S0 <=     O6_I15_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O6_N0_S1;		always @(posedge clk) O6_N0_S1 <=     O6_N0_S0  +  O6_N2_S0 ;
 logic signed [31:0] O6_N2_S1;		always @(posedge clk) O6_N2_S1 <=     O6_N4_S0  +  O6_N6_S0 ;
 logic signed [31:0] O6_N4_S1;		always @(posedge clk) O6_N4_S1 <=     O6_N8_S0  +  O6_N10_S0 ;
 logic signed [31:0] O6_N6_S1;		always @(posedge clk) O6_N6_S1 <=     O6_N12_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O6_N0_S2;		always @(posedge clk) O6_N0_S2 <=     O6_N0_S1  +  O6_N2_S1 ;
 logic signed [31:0] O6_N2_S2;		always @(posedge clk) O6_N2_S2 <=     O6_N4_S1  +  O6_N6_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O6_N0_S3;		always @(posedge clk) O6_N0_S3 <=     O6_N0_S2  +  O6_N2_S2 ;
 assign conv_mac_6 = O6_N0_S3;

logic signed [31:0] conv_mac_7;
logic signed [31:0] O7_N0_S0;		always @(posedge clk) O7_N0_S0 <=     O7_I0_R0_C0_SM1   +  O7_I2_R0_C0_SM1  ;
 logic signed [31:0] O7_N2_S0;		always @(posedge clk) O7_N2_S0 <=     O7_I4_R0_C0_SM1   +  O7_I5_R0_C0_SM1  ;
 logic signed [31:0] O7_N4_S0;		always @(posedge clk) O7_N4_S0 <=     O7_I7_R0_C0_SM1   +  O7_I8_R0_C0_SM1  ;
 logic signed [31:0] O7_N6_S0;		always @(posedge clk) O7_N6_S0 <=     O7_I9_R0_C0_SM1   +  O7_I10_R0_C0_SM1  ;
 logic signed [31:0] O7_N8_S0;		always @(posedge clk) O7_N8_S0 <=     O7_I11_R0_C0_SM1   +  O7_I13_R0_C0_SM1  ;
 logic signed [31:0] O7_N10_S0;		always @(posedge clk) O7_N10_S0 <=     O7_I14_R0_C0_SM1   +  O7_I15_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O7_N0_S1;		always @(posedge clk) O7_N0_S1 <=     O7_N0_S0  +  O7_N2_S0 ;
 logic signed [31:0] O7_N2_S1;		always @(posedge clk) O7_N2_S1 <=     O7_N4_S0  +  O7_N6_S0 ;
 logic signed [31:0] O7_N4_S1;		always @(posedge clk) O7_N4_S1 <=     O7_N8_S0  +  O7_N10_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O7_N0_S2;		always @(posedge clk) O7_N0_S2 <=     O7_N0_S1  +  O7_N2_S1 ;
 logic signed [31:0] O7_N2_S2;		always @(posedge clk) O7_N2_S2 <=     O7_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O7_N0_S3;		always @(posedge clk) O7_N0_S3 <=     O7_N0_S2  +  O7_N2_S2 ;
 assign conv_mac_7 = O7_N0_S3;

logic signed [31:0] conv_mac_8;
logic signed [31:0] O8_N0_S0;		always @(posedge clk) O8_N0_S0 <=     O8_I0_R0_C0_SM1   +  O8_I3_R0_C0_SM1  ;
 logic signed [31:0] O8_N2_S0;		always @(posedge clk) O8_N2_S0 <=     O8_I5_R0_C0_SM1   +  O8_I9_R0_C0_SM1  ;
 logic signed [31:0] O8_N4_S0;		always @(posedge clk) O8_N4_S0 <=     O8_I10_R0_C0_SM1   +  O8_I12_R0_C0_SM1  ;
 logic signed [31:0] O8_N6_S0;		always @(posedge clk) O8_N6_S0 <=     O8_I14_R0_C0_SM1   +  O8_I15_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O8_N0_S1;		always @(posedge clk) O8_N0_S1 <=     O8_N0_S0  +  O8_N2_S0 ;
 logic signed [31:0] O8_N2_S1;		always @(posedge clk) O8_N2_S1 <=     O8_N4_S0  +  O8_N6_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O8_N0_S2;		always @(posedge clk) O8_N0_S2 <=     O8_N0_S1  +  O8_N2_S1 ;
 assign conv_mac_8 = O8_N0_S2;

logic signed [31:0] conv_mac_9;
logic signed [31:0] O9_N0_S0;		always @(posedge clk) O9_N0_S0 <=     O9_I1_R0_C0_SM1   +  O9_I2_R0_C0_SM1  ;
 logic signed [31:0] O9_N2_S0;		always @(posedge clk) O9_N2_S0 <=     O9_I3_R0_C0_SM1   +  O9_I6_R0_C0_SM1  ;
 logic signed [31:0] O9_N4_S0;		always @(posedge clk) O9_N4_S0 <=     O9_I8_R0_C0_SM1   +  O9_I11_R0_C0_SM1  ;
 logic signed [31:0] O9_N6_S0;		always @(posedge clk) O9_N6_S0 <=     O9_I13_R0_C0_SM1   +  O9_I15_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O9_N0_S1;		always @(posedge clk) O9_N0_S1 <=     O9_N0_S0  +  O9_N2_S0 ;
 logic signed [31:0] O9_N2_S1;		always @(posedge clk) O9_N2_S1 <=     O9_N4_S0  +  O9_N6_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O9_N0_S2;		always @(posedge clk) O9_N0_S2 <=     O9_N0_S1  +  O9_N2_S1 ;
 assign conv_mac_9 = O9_N0_S2;

logic signed [31:0] conv_mac_10;
logic signed [31:0] O10_N0_S0;		always @(posedge clk) O10_N0_S0 <=     O10_I0_R0_C0_SM1   +  O10_I1_R0_C0_SM1  ;
 logic signed [31:0] O10_N2_S0;		always @(posedge clk) O10_N2_S0 <=     O10_I2_R0_C0_SM1   +  O10_I3_R0_C0_SM1  ;
 logic signed [31:0] O10_N4_S0;		always @(posedge clk) O10_N4_S0 <=     O10_I5_R0_C0_SM1   +  O10_I7_R0_C0_SM1  ;
 logic signed [31:0] O10_N6_S0;		always @(posedge clk) O10_N6_S0 <=     O10_I8_R0_C0_SM1   +  O10_I9_R0_C0_SM1  ;
 logic signed [31:0] O10_N8_S0;		always @(posedge clk) O10_N8_S0 <=     O10_I10_R0_C0_SM1   +  O10_I11_R0_C0_SM1  ;
 logic signed [31:0] O10_N10_S0;		always @(posedge clk) O10_N10_S0 <=     O10_I12_R0_C0_SM1   +  O10_I15_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O10_N0_S1;		always @(posedge clk) O10_N0_S1 <=     O10_N0_S0  +  O10_N2_S0 ;
 logic signed [31:0] O10_N2_S1;		always @(posedge clk) O10_N2_S1 <=     O10_N4_S0  +  O10_N6_S0 ;
 logic signed [31:0] O10_N4_S1;		always @(posedge clk) O10_N4_S1 <=     O10_N8_S0  +  O10_N10_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O10_N0_S2;		always @(posedge clk) O10_N0_S2 <=     O10_N0_S1  +  O10_N2_S1 ;
 logic signed [31:0] O10_N2_S2;		always @(posedge clk) O10_N2_S2 <=     O10_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O10_N0_S3;		always @(posedge clk) O10_N0_S3 <=     O10_N0_S2  +  O10_N2_S2 ;
 assign conv_mac_10 = O10_N0_S3;

logic signed [31:0] conv_mac_11;
logic signed [31:0] O11_N0_S0;		always @(posedge clk) O11_N0_S0 <=     O11_I1_R0_C0_SM1   +  O11_I3_R0_C0_SM1  ;
 logic signed [31:0] O11_N2_S0;		always @(posedge clk) O11_N2_S0 <=     O11_I4_R0_C0_SM1   +  O11_I5_R0_C0_SM1  ;
 logic signed [31:0] O11_N4_S0;		always @(posedge clk) O11_N4_S0 <=     O11_I7_R0_C0_SM1   +  O11_I8_R0_C0_SM1  ;
 logic signed [31:0] O11_N6_S0;		always @(posedge clk) O11_N6_S0 <=     O11_I10_R0_C0_SM1   +  O11_I11_R0_C0_SM1  ;
 logic signed [31:0] O11_N8_S0;		always @(posedge clk) O11_N8_S0 <=     O11_I12_R0_C0_SM1   +  O11_I13_R0_C0_SM1  ;
 logic signed [31:0] O11_N10_S0;		always @(posedge clk) O11_N10_S0 <=     O11_I14_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O11_N0_S1;		always @(posedge clk) O11_N0_S1 <=     O11_N0_S0  +  O11_N2_S0 ;
 logic signed [31:0] O11_N2_S1;		always @(posedge clk) O11_N2_S1 <=     O11_N4_S0  +  O11_N6_S0 ;
 logic signed [31:0] O11_N4_S1;		always @(posedge clk) O11_N4_S1 <=     O11_N8_S0  +  O11_N10_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O11_N0_S2;		always @(posedge clk) O11_N0_S2 <=     O11_N0_S1  +  O11_N2_S1 ;
 logic signed [31:0] O11_N2_S2;		always @(posedge clk) O11_N2_S2 <=     O11_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O11_N0_S3;		always @(posedge clk) O11_N0_S3 <=     O11_N0_S2  +  O11_N2_S2 ;
 assign conv_mac_11 = O11_N0_S3;

logic signed [31:0] conv_mac_12;
logic signed [31:0] O12_N0_S0;		always @(posedge clk) O12_N0_S0 <=     O12_I1_R0_C0_SM1   +  O12_I2_R0_C0_SM1  ;
 logic signed [31:0] O12_N2_S0;		always @(posedge clk) O12_N2_S0 <=     O12_I5_R0_C0_SM1   +  O12_I6_R0_C0_SM1  ;
 logic signed [31:0] O12_N4_S0;		always @(posedge clk) O12_N4_S0 <=     O12_I8_R0_C0_SM1   +  O12_I12_R0_C0_SM1  ;
 logic signed [31:0] O12_N6_S0;		always @(posedge clk) O12_N6_S0 <=     O12_I13_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O12_N0_S1;		always @(posedge clk) O12_N0_S1 <=     O12_N0_S0  +  O12_N2_S0 ;
 logic signed [31:0] O12_N2_S1;		always @(posedge clk) O12_N2_S1 <=     O12_N4_S0  +  O12_N6_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O12_N0_S2;		always @(posedge clk) O12_N0_S2 <=     O12_N0_S1  +  O12_N2_S1 ;
 assign conv_mac_12 = O12_N0_S2;

logic signed [31:0] conv_mac_13;
logic signed [31:0] O13_N0_S0;		always @(posedge clk) O13_N0_S0 <=     O13_I0_R0_C0_SM1   +  O13_I2_R0_C0_SM1  ;
 logic signed [31:0] O13_N2_S0;		always @(posedge clk) O13_N2_S0 <=     O13_I5_R0_C0_SM1   +  O13_I12_R0_C0_SM1  ;
 logic signed [31:0] O13_N4_S0;		always @(posedge clk) O13_N4_S0 <=     O13_I15_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O13_N0_S1;		always @(posedge clk) O13_N0_S1 <=     O13_N0_S0  +  O13_N2_S0 ;
 logic signed [31:0] O13_N2_S1;		always @(posedge clk) O13_N2_S1 <=     O13_N4_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O13_N0_S2;		always @(posedge clk) O13_N0_S2 <=     O13_N0_S1  +  O13_N2_S1 ;
 assign conv_mac_13 = O13_N0_S2;

logic signed [31:0] conv_mac_14;
logic signed [31:0] O14_N0_S0;		always @(posedge clk) O14_N0_S0 <=     O14_I0_R0_C0_SM1   +  O14_I5_R0_C0_SM1  ;
 logic signed [31:0] O14_N2_S0;		always @(posedge clk) O14_N2_S0 <=     O14_I7_R0_C0_SM1   +  O14_I9_R0_C0_SM1  ;
 logic signed [31:0] O14_N4_S0;		always @(posedge clk) O14_N4_S0 <=     O14_I10_R0_C0_SM1   +  O14_I11_R0_C0_SM1  ;
 logic signed [31:0] O14_N6_S0;		always @(posedge clk) O14_N6_S0 <=     O14_I12_R0_C0_SM1   +  O14_I14_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O14_N0_S1;		always @(posedge clk) O14_N0_S1 <=     O14_N0_S0  +  O14_N2_S0 ;
 logic signed [31:0] O14_N2_S1;		always @(posedge clk) O14_N2_S1 <=     O14_N4_S0  +  O14_N6_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O14_N0_S2;		always @(posedge clk) O14_N0_S2 <=     O14_N0_S1  +  O14_N2_S1 ;
 assign conv_mac_14 = O14_N0_S2;

logic signed [31:0] conv_mac_15;
logic signed [31:0] O15_N0_S0;		always @(posedge clk) O15_N0_S0 <=     O15_I0_R0_C0_SM1   +  O15_I1_R0_C0_SM1  ;
 logic signed [31:0] O15_N2_S0;		always @(posedge clk) O15_N2_S0 <=     O15_I4_R0_C0_SM1   +  O15_I6_R0_C0_SM1  ;
 logic signed [31:0] O15_N4_S0;		always @(posedge clk) O15_N4_S0 <=     O15_I7_R0_C0_SM1   +  O15_I9_R0_C0_SM1  ;
 logic signed [31:0] O15_N6_S0;		always @(posedge clk) O15_N6_S0 <=     O15_I10_R0_C0_SM1   +  O15_I11_R0_C0_SM1  ;
 logic signed [31:0] O15_N8_S0;		always @(posedge clk) O15_N8_S0 <=     O15_I12_R0_C0_SM1   +  O15_I15_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O15_N0_S1;		always @(posedge clk) O15_N0_S1 <=     O15_N0_S0  +  O15_N2_S0 ;
 logic signed [31:0] O15_N2_S1;		always @(posedge clk) O15_N2_S1 <=     O15_N4_S0  +  O15_N6_S0 ;
 logic signed [31:0] O15_N4_S1;		always @(posedge clk) O15_N4_S1 <=     O15_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O15_N0_S2;		always @(posedge clk) O15_N0_S2 <=     O15_N0_S1  +  O15_N2_S1 ;
 logic signed [31:0] O15_N2_S2;		always @(posedge clk) O15_N2_S2 <=     O15_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O15_N0_S3;		always @(posedge clk) O15_N0_S3 <=     O15_N0_S2  +  O15_N2_S2 ;
 assign conv_mac_15 = O15_N0_S3;

logic signed [31:0] conv_mac_16;
logic signed [31:0] O16_N0_S0;		always @(posedge clk) O16_N0_S0 <=     O16_I1_R0_C0_SM1   +  O16_I4_R0_C0_SM1  ;
 logic signed [31:0] O16_N2_S0;		always @(posedge clk) O16_N2_S0 <=     O16_I8_R0_C0_SM1   +  O16_I11_R0_C0_SM1  ;
 logic signed [31:0] O16_N4_S0;		always @(posedge clk) O16_N4_S0 <=     O16_I13_R0_C0_SM1   +  O16_I14_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O16_N0_S1;		always @(posedge clk) O16_N0_S1 <=     O16_N0_S0  +  O16_N2_S0 ;
 logic signed [31:0] O16_N2_S1;		always @(posedge clk) O16_N2_S1 <=     O16_N4_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O16_N0_S2;		always @(posedge clk) O16_N0_S2 <=     O16_N0_S1  +  O16_N2_S1 ;
 assign conv_mac_16 = O16_N0_S2;

logic signed [31:0] conv_mac_17;
logic signed [31:0] O17_N0_S0;		always @(posedge clk) O17_N0_S0 <=     O17_I0_R0_C0_SM1   +  O17_I2_R0_C0_SM1  ;
 logic signed [31:0] O17_N2_S0;		always @(posedge clk) O17_N2_S0 <=     O17_I4_R0_C0_SM1   +  O17_I5_R0_C0_SM1  ;
 logic signed [31:0] O17_N4_S0;		always @(posedge clk) O17_N4_S0 <=     O17_I6_R0_C0_SM1   +  O17_I9_R0_C0_SM1  ;
 logic signed [31:0] O17_N6_S0;		always @(posedge clk) O17_N6_S0 <=     O17_I11_R0_C0_SM1   +  O17_I12_R0_C0_SM1  ;
 logic signed [31:0] O17_N8_S0;		always @(posedge clk) O17_N8_S0 <=     O17_I15_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O17_N0_S1;		always @(posedge clk) O17_N0_S1 <=     O17_N0_S0  +  O17_N2_S0 ;
 logic signed [31:0] O17_N2_S1;		always @(posedge clk) O17_N2_S1 <=     O17_N4_S0  +  O17_N6_S0 ;
 logic signed [31:0] O17_N4_S1;		always @(posedge clk) O17_N4_S1 <=     O17_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O17_N0_S2;		always @(posedge clk) O17_N0_S2 <=     O17_N0_S1  +  O17_N2_S1 ;
 logic signed [31:0] O17_N2_S2;		always @(posedge clk) O17_N2_S2 <=     O17_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O17_N0_S3;		always @(posedge clk) O17_N0_S3 <=     O17_N0_S2  +  O17_N2_S2 ;
 assign conv_mac_17 = O17_N0_S3;

logic signed [31:0] conv_mac_18;
logic signed [31:0] O18_N0_S0;		always @(posedge clk) O18_N0_S0 <=     O18_I0_R0_C0_SM1   +  O18_I5_R0_C0_SM1  ;
 logic signed [31:0] O18_N2_S0;		always @(posedge clk) O18_N2_S0 <=     O18_I9_R0_C0_SM1   +  O18_I10_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O18_N0_S1;		always @(posedge clk) O18_N0_S1 <=     O18_N0_S0  +  O18_N2_S0 ;
 assign conv_mac_18 = O18_N0_S1;

logic signed [31:0] conv_mac_19;
logic signed [31:0] O19_N0_S0;		always @(posedge clk) O19_N0_S0 <=     O19_I0_R0_C0_SM1   +  O19_I6_R0_C0_SM1  ;
 logic signed [31:0] O19_N2_S0;		always @(posedge clk) O19_N2_S0 <=     O19_I11_R0_C0_SM1   +  O19_I13_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O19_N0_S1;		always @(posedge clk) O19_N0_S1 <=     O19_N0_S0  +  O19_N2_S0 ;
 assign conv_mac_19 = O19_N0_S1;

logic signed [31:0] conv_mac_20;
logic signed [31:0] O20_N0_S0;		always @(posedge clk) O20_N0_S0 <=     O20_I11_R0_C0_SM1   +  O20_I13_R0_C0_SM1  ;
 assign conv_mac_20 = O20_N0_S0;

logic signed [31:0] conv_mac_21;
logic signed [31:0] O21_N0_S0;		always @(posedge clk) O21_N0_S0 <=     O21_I2_R0_C0_SM1   +  O21_I3_R0_C0_SM1  ;
 logic signed [31:0] O21_N2_S0;		always @(posedge clk) O21_N2_S0 <=     O21_I5_R0_C0_SM1   +  O21_I6_R0_C0_SM1  ;
 logic signed [31:0] O21_N4_S0;		always @(posedge clk) O21_N4_S0 <=     O21_I7_R0_C0_SM1   +  O21_I8_R0_C0_SM1  ;
 logic signed [31:0] O21_N6_S0;		always @(posedge clk) O21_N6_S0 <=     O21_I10_R0_C0_SM1   +  O21_I11_R0_C0_SM1  ;
 logic signed [31:0] O21_N8_S0;		always @(posedge clk) O21_N8_S0 <=     O21_I14_R0_C0_SM1   +  O21_I15_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O21_N0_S1;		always @(posedge clk) O21_N0_S1 <=     O21_N0_S0  +  O21_N2_S0 ;
 logic signed [31:0] O21_N2_S1;		always @(posedge clk) O21_N2_S1 <=     O21_N4_S0  +  O21_N6_S0 ;
 logic signed [31:0] O21_N4_S1;		always @(posedge clk) O21_N4_S1 <=     O21_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O21_N0_S2;		always @(posedge clk) O21_N0_S2 <=     O21_N0_S1  +  O21_N2_S1 ;
 logic signed [31:0] O21_N2_S2;		always @(posedge clk) O21_N2_S2 <=     O21_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O21_N0_S3;		always @(posedge clk) O21_N0_S3 <=     O21_N0_S2  +  O21_N2_S2 ;
 assign conv_mac_21 = O21_N0_S3;

logic signed [31:0] conv_mac_22;
logic signed [31:0] O22_N0_S0;		always @(posedge clk) O22_N0_S0 <=     O22_I0_R0_C0_SM1   +  O22_I2_R0_C0_SM1  ;
 logic signed [31:0] O22_N2_S0;		always @(posedge clk) O22_N2_S0 <=     O22_I5_R0_C0_SM1   +  O22_I8_R0_C0_SM1  ;
 logic signed [31:0] O22_N4_S0;		always @(posedge clk) O22_N4_S0 <=     O22_I9_R0_C0_SM1   +  O22_I10_R0_C0_SM1  ;
 logic signed [31:0] O22_N6_S0;		always @(posedge clk) O22_N6_S0 <=     O22_I11_R0_C0_SM1   +  O22_I12_R0_C0_SM1  ;
 logic signed [31:0] O22_N8_S0;		always @(posedge clk) O22_N8_S0 <=     O22_I15_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O22_N0_S1;		always @(posedge clk) O22_N0_S1 <=     O22_N0_S0  +  O22_N2_S0 ;
 logic signed [31:0] O22_N2_S1;		always @(posedge clk) O22_N2_S1 <=     O22_N4_S0  +  O22_N6_S0 ;
 logic signed [31:0] O22_N4_S1;		always @(posedge clk) O22_N4_S1 <=     O22_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O22_N0_S2;		always @(posedge clk) O22_N0_S2 <=     O22_N0_S1  +  O22_N2_S1 ;
 logic signed [31:0] O22_N2_S2;		always @(posedge clk) O22_N2_S2 <=     O22_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O22_N0_S3;		always @(posedge clk) O22_N0_S3 <=     O22_N0_S2  +  O22_N2_S2 ;
 assign conv_mac_22 = O22_N0_S3;

logic signed [31:0] conv_mac_23;
logic signed [31:0] O23_N0_S0;		always @(posedge clk) O23_N0_S0 <=     O23_I1_R0_C0_SM1   +  O23_I3_R0_C0_SM1  ;
 logic signed [31:0] O23_N2_S0;		always @(posedge clk) O23_N2_S0 <=     O23_I4_R0_C0_SM1   +  O23_I5_R0_C0_SM1  ;
 logic signed [31:0] O23_N4_S0;		always @(posedge clk) O23_N4_S0 <=     O23_I8_R0_C0_SM1   +  O23_I11_R0_C0_SM1  ;
 logic signed [31:0] O23_N6_S0;		always @(posedge clk) O23_N6_S0 <=     O23_I12_R0_C0_SM1   +  O23_I13_R0_C0_SM1  ;
 logic signed [31:0] O23_N8_S0;		always @(posedge clk) O23_N8_S0 <=     O23_I14_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O23_N0_S1;		always @(posedge clk) O23_N0_S1 <=     O23_N0_S0  +  O23_N2_S0 ;
 logic signed [31:0] O23_N2_S1;		always @(posedge clk) O23_N2_S1 <=     O23_N4_S0  +  O23_N6_S0 ;
 logic signed [31:0] O23_N4_S1;		always @(posedge clk) O23_N4_S1 <=     O23_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O23_N0_S2;		always @(posedge clk) O23_N0_S2 <=     O23_N0_S1  +  O23_N2_S1 ;
 logic signed [31:0] O23_N2_S2;		always @(posedge clk) O23_N2_S2 <=     O23_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O23_N0_S3;		always @(posedge clk) O23_N0_S3 <=     O23_N0_S2  +  O23_N2_S2 ;
 assign conv_mac_23 = O23_N0_S3;

logic signed [31:0] conv_mac_24;
logic signed [31:0] O24_N0_S0;		always @(posedge clk) O24_N0_S0 <=     O24_I0_R0_C0_SM1   +  O24_I1_R0_C0_SM1  ;
 logic signed [31:0] O24_N2_S0;		always @(posedge clk) O24_N2_S0 <=     O24_I2_R0_C0_SM1   +  O24_I3_R0_C0_SM1  ;
 logic signed [31:0] O24_N4_S0;		always @(posedge clk) O24_N4_S0 <=     O24_I4_R0_C0_SM1   +  O24_I5_R0_C0_SM1  ;
 logic signed [31:0] O24_N6_S0;		always @(posedge clk) O24_N6_S0 <=     O24_I6_R0_C0_SM1   +  O24_I7_R0_C0_SM1  ;
 logic signed [31:0] O24_N8_S0;		always @(posedge clk) O24_N8_S0 <=     O24_I8_R0_C0_SM1   +  O24_I9_R0_C0_SM1  ;
 logic signed [31:0] O24_N10_S0;		always @(posedge clk) O24_N10_S0 <=     O24_I10_R0_C0_SM1   +  O24_I11_R0_C0_SM1  ;
 logic signed [31:0] O24_N12_S0;		always @(posedge clk) O24_N12_S0 <=     O24_I13_R0_C0_SM1   +  O24_I14_R0_C0_SM1  ;
 logic signed [31:0] O24_N14_S0;		always @(posedge clk) O24_N14_S0 <=     O24_I15_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O24_N0_S1;		always @(posedge clk) O24_N0_S1 <=     O24_N0_S0  +  O24_N2_S0 ;
 logic signed [31:0] O24_N2_S1;		always @(posedge clk) O24_N2_S1 <=     O24_N4_S0  +  O24_N6_S0 ;
 logic signed [31:0] O24_N4_S1;		always @(posedge clk) O24_N4_S1 <=     O24_N8_S0  +  O24_N10_S0 ;
 logic signed [31:0] O24_N6_S1;		always @(posedge clk) O24_N6_S1 <=     O24_N12_S0  +  O24_N14_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O24_N0_S2;		always @(posedge clk) O24_N0_S2 <=     O24_N0_S1  +  O24_N2_S1 ;
 logic signed [31:0] O24_N2_S2;		always @(posedge clk) O24_N2_S2 <=     O24_N4_S1  +  O24_N6_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O24_N0_S3;		always @(posedge clk) O24_N0_S3 <=     O24_N0_S2  +  O24_N2_S2 ;
 assign conv_mac_24 = O24_N0_S3;

logic signed [31:0] conv_mac_25;
logic signed [31:0] O25_N0_S0;		always @(posedge clk) O25_N0_S0 <=     O25_I1_R0_C0_SM1   +  O25_I3_R0_C0_SM1  ;
 logic signed [31:0] O25_N2_S0;		always @(posedge clk) O25_N2_S0 <=     O25_I5_R0_C0_SM1   +  O25_I6_R0_C0_SM1  ;
 logic signed [31:0] O25_N4_S0;		always @(posedge clk) O25_N4_S0 <=     O25_I7_R0_C0_SM1   +  O25_I8_R0_C0_SM1  ;
 logic signed [31:0] O25_N6_S0;		always @(posedge clk) O25_N6_S0 <=     O25_I9_R0_C0_SM1   +  O25_I10_R0_C0_SM1  ;
 logic signed [31:0] O25_N8_S0;		always @(posedge clk) O25_N8_S0 <=     O25_I11_R0_C0_SM1   +  O25_I12_R0_C0_SM1  ;
 logic signed [31:0] O25_N10_S0;		always @(posedge clk) O25_N10_S0 <=     O25_I14_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O25_N0_S1;		always @(posedge clk) O25_N0_S1 <=     O25_N0_S0  +  O25_N2_S0 ;
 logic signed [31:0] O25_N2_S1;		always @(posedge clk) O25_N2_S1 <=     O25_N4_S0  +  O25_N6_S0 ;
 logic signed [31:0] O25_N4_S1;		always @(posedge clk) O25_N4_S1 <=     O25_N8_S0  +  O25_N10_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O25_N0_S2;		always @(posedge clk) O25_N0_S2 <=     O25_N0_S1  +  O25_N2_S1 ;
 logic signed [31:0] O25_N2_S2;		always @(posedge clk) O25_N2_S2 <=     O25_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O25_N0_S3;		always @(posedge clk) O25_N0_S3 <=     O25_N0_S2  +  O25_N2_S2 ;
 assign conv_mac_25 = O25_N0_S3;

logic signed [31:0] conv_mac_26;
logic signed [31:0] O26_N0_S0;		always @(posedge clk) O26_N0_S0 <=     O26_I1_R0_C0_SM1   +  O26_I2_R0_C0_SM1  ;
 logic signed [31:0] O26_N2_S0;		always @(posedge clk) O26_N2_S0 <=     O26_I3_R0_C0_SM1   +  O26_I4_R0_C0_SM1  ;
 logic signed [31:0] O26_N4_S0;		always @(posedge clk) O26_N4_S0 <=     O26_I6_R0_C0_SM1   +  O26_I8_R0_C0_SM1  ;
 logic signed [31:0] O26_N6_S0;		always @(posedge clk) O26_N6_S0 <=     O26_I11_R0_C0_SM1   +  O26_I14_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O26_N0_S1;		always @(posedge clk) O26_N0_S1 <=     O26_N0_S0  +  O26_N2_S0 ;
 logic signed [31:0] O26_N2_S1;		always @(posedge clk) O26_N2_S1 <=     O26_N4_S0  +  O26_N6_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O26_N0_S2;		always @(posedge clk) O26_N0_S2 <=     O26_N0_S1  +  O26_N2_S1 ;
 assign conv_mac_26 = O26_N0_S2;

logic signed [31:0] conv_mac_27;
logic signed [31:0] O27_N0_S0;		always @(posedge clk) O27_N0_S0 <=     O27_I0_R0_C0_SM1   +  O27_I5_R0_C0_SM1  ;
 logic signed [31:0] O27_N2_S0;		always @(posedge clk) O27_N2_S0 <=     O27_I12_R0_C0_SM1   +  O27_I15_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O27_N0_S1;		always @(posedge clk) O27_N0_S1 <=     O27_N0_S0  +  O27_N2_S0 ;
 assign conv_mac_27 = O27_N0_S1;

logic signed [31:0] conv_mac_28;
logic signed [31:0] O28_N0_S0;		always @(posedge clk) O28_N0_S0 <=     O28_I0_R0_C0_SM1   +  O28_I1_R0_C0_SM1  ;
 logic signed [31:0] O28_N2_S0;		always @(posedge clk) O28_N2_S0 <=     O28_I3_R0_C0_SM1   +  O28_I4_R0_C0_SM1  ;
 logic signed [31:0] O28_N4_S0;		always @(posedge clk) O28_N4_S0 <=     O28_I5_R0_C0_SM1   +  O28_I6_R0_C0_SM1  ;
 logic signed [31:0] O28_N6_S0;		always @(posedge clk) O28_N6_S0 <=     O28_I7_R0_C0_SM1   +  O28_I8_R0_C0_SM1  ;
 logic signed [31:0] O28_N8_S0;		always @(posedge clk) O28_N8_S0 <=     O28_I9_R0_C0_SM1   +  O28_I10_R0_C0_SM1  ;
 logic signed [31:0] O28_N10_S0;		always @(posedge clk) O28_N10_S0 <=     O28_I12_R0_C0_SM1   +  O28_I14_R0_C0_SM1  ;
 logic signed [31:0] O28_N12_S0;		always @(posedge clk) O28_N12_S0 <=     O28_I15_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O28_N0_S1;		always @(posedge clk) O28_N0_S1 <=     O28_N0_S0  +  O28_N2_S0 ;
 logic signed [31:0] O28_N2_S1;		always @(posedge clk) O28_N2_S1 <=     O28_N4_S0  +  O28_N6_S0 ;
 logic signed [31:0] O28_N4_S1;		always @(posedge clk) O28_N4_S1 <=     O28_N8_S0  +  O28_N10_S0 ;
 logic signed [31:0] O28_N6_S1;		always @(posedge clk) O28_N6_S1 <=     O28_N12_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O28_N0_S2;		always @(posedge clk) O28_N0_S2 <=     O28_N0_S1  +  O28_N2_S1 ;
 logic signed [31:0] O28_N2_S2;		always @(posedge clk) O28_N2_S2 <=     O28_N4_S1  +  O28_N6_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O28_N0_S3;		always @(posedge clk) O28_N0_S3 <=     O28_N0_S2  +  O28_N2_S2 ;
 assign conv_mac_28 = O28_N0_S3;

logic signed [31:0] conv_mac_29;
logic signed [31:0] O29_N0_S0;		always @(posedge clk) O29_N0_S0 <=     O29_I0_R0_C0_SM1   +  O29_I1_R0_C0_SM1  ;
 logic signed [31:0] O29_N2_S0;		always @(posedge clk) O29_N2_S0 <=     O29_I5_R0_C0_SM1   +  O29_I7_R0_C0_SM1  ;
 logic signed [31:0] O29_N4_S0;		always @(posedge clk) O29_N4_S0 <=     O29_I9_R0_C0_SM1   +  O29_I10_R0_C0_SM1  ;
 logic signed [31:0] O29_N6_S0;		always @(posedge clk) O29_N6_S0 <=     O29_I12_R0_C0_SM1   +  O29_I14_R0_C0_SM1  ;
 logic signed [31:0] O29_N8_S0;		always @(posedge clk) O29_N8_S0 <=     O29_I15_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O29_N0_S1;		always @(posedge clk) O29_N0_S1 <=     O29_N0_S0  +  O29_N2_S0 ;
 logic signed [31:0] O29_N2_S1;		always @(posedge clk) O29_N2_S1 <=     O29_N4_S0  +  O29_N6_S0 ;
 logic signed [31:0] O29_N4_S1;		always @(posedge clk) O29_N4_S1 <=     O29_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O29_N0_S2;		always @(posedge clk) O29_N0_S2 <=     O29_N0_S1  +  O29_N2_S1 ;
 logic signed [31:0] O29_N2_S2;		always @(posedge clk) O29_N2_S2 <=     O29_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O29_N0_S3;		always @(posedge clk) O29_N0_S3 <=     O29_N0_S2  +  O29_N2_S2 ;
 assign conv_mac_29 = O29_N0_S3;

logic signed [31:0] conv_mac_30;
logic signed [31:0] O30_N0_S0;		always @(posedge clk) O30_N0_S0 <=     O30_I0_R0_C0_SM1   +  O30_I1_R0_C0_SM1  ;
 logic signed [31:0] O30_N2_S0;		always @(posedge clk) O30_N2_S0 <=     O30_I2_R0_C0_SM1   +  O30_I3_R0_C0_SM1  ;
 logic signed [31:0] O30_N4_S0;		always @(posedge clk) O30_N4_S0 <=     O30_I6_R0_C0_SM1   +  O30_I8_R0_C0_SM1  ;
 logic signed [31:0] O30_N6_S0;		always @(posedge clk) O30_N6_S0 <=     O30_I11_R0_C0_SM1   +  O30_I12_R0_C0_SM1  ;
 logic signed [31:0] O30_N8_S0;		always @(posedge clk) O30_N8_S0 <=     O30_I13_R0_C0_SM1   +  O30_I14_R0_C0_SM1  ;
 logic signed [31:0] O30_N10_S0;		always @(posedge clk) O30_N10_S0 <=     O30_I15_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O30_N0_S1;		always @(posedge clk) O30_N0_S1 <=     O30_N0_S0  +  O30_N2_S0 ;
 logic signed [31:0] O30_N2_S1;		always @(posedge clk) O30_N2_S1 <=     O30_N4_S0  +  O30_N6_S0 ;
 logic signed [31:0] O30_N4_S1;		always @(posedge clk) O30_N4_S1 <=     O30_N8_S0  +  O30_N10_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O30_N0_S2;		always @(posedge clk) O30_N0_S2 <=     O30_N0_S1  +  O30_N2_S1 ;
 logic signed [31:0] O30_N2_S2;		always @(posedge clk) O30_N2_S2 <=     O30_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O30_N0_S3;		always @(posedge clk) O30_N0_S3 <=     O30_N0_S2  +  O30_N2_S2 ;
 assign conv_mac_30 = O30_N0_S3;

logic signed [31:0] conv_mac_31;
logic signed [31:0] O31_N0_S0;		always @(posedge clk) O31_N0_S0 <=     O31_I0_R0_C0_SM1   +  O31_I1_R0_C0_SM1  ;
 logic signed [31:0] O31_N2_S0;		always @(posedge clk) O31_N2_S0 <=     O31_I2_R0_C0_SM1   +  O31_I3_R0_C0_SM1  ;
 logic signed [31:0] O31_N4_S0;		always @(posedge clk) O31_N4_S0 <=     O31_I4_R0_C0_SM1   +  O31_I8_R0_C0_SM1  ;
 logic signed [31:0] O31_N6_S0;		always @(posedge clk) O31_N6_S0 <=     O31_I11_R0_C0_SM1   +  O31_I12_R0_C0_SM1  ;
 logic signed [31:0] O31_N8_S0;		always @(posedge clk) O31_N8_S0 <=     O31_I13_R0_C0_SM1   +  O31_I15_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O31_N0_S1;		always @(posedge clk) O31_N0_S1 <=     O31_N0_S0  +  O31_N2_S0 ;
 logic signed [31:0] O31_N2_S1;		always @(posedge clk) O31_N2_S1 <=     O31_N4_S0  +  O31_N6_S0 ;
 logic signed [31:0] O31_N4_S1;		always @(posedge clk) O31_N4_S1 <=     O31_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O31_N0_S2;		always @(posedge clk) O31_N0_S2 <=     O31_N0_S1  +  O31_N2_S1 ;
 logic signed [31:0] O31_N2_S2;		always @(posedge clk) O31_N2_S2 <=     O31_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O31_N0_S3;		always @(posedge clk) O31_N0_S3 <=     O31_N0_S2  +  O31_N2_S2 ;
 assign conv_mac_31 = O31_N0_S3;

logic valid_D1;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D1<= 0 ;
	else valid_D1<=valid;
end
logic valid_D2;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D2<= 0 ;
	else valid_D2<=valid_D1;
end
logic valid_D3;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D3<= 0 ;
	else valid_D3<=valid_D2;
end
logic valid_D4;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D4<= 0 ;
	else valid_D4<=valid_D3;
end
logic valid_D5;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D5<= 0 ;
	else valid_D5<=valid_D4;
end
always_ff @(posedge clk) begin
	if (rstn == 0) ready <= 0 ;
	else ready <=valid_D5;
end
logic [31:0] bias_add_0;
assign bias_add_0 = conv_mac_0 + 6'd20;
logic [31:0] bias_add_1;
assign bias_add_1 = conv_mac_1 + 6'd29;
logic [31:0] bias_add_2;
assign bias_add_2 = conv_mac_2 + 6'd31;
logic [31:0] bias_add_3;
assign bias_add_3 = conv_mac_3 + 6'd17;
logic [31:0] bias_add_4;
assign bias_add_4 = conv_mac_4;
logic [31:0] bias_add_5;
assign bias_add_5 = conv_mac_5 + 5'd12;
logic [31:0] bias_add_6;
assign bias_add_6 = conv_mac_6 + 7'd36;
logic [31:0] bias_add_7;
assign bias_add_7 = conv_mac_7 + 6'd31;
logic [31:0] bias_add_8;
assign bias_add_8 = conv_mac_8 + 5'd13;
logic [31:0] bias_add_9;
assign bias_add_9 = conv_mac_9 + 6'd22;
logic [31:0] bias_add_10;
assign bias_add_10 = conv_mac_10 - 5'd8;
logic [31:0] bias_add_11;
assign bias_add_11 = conv_mac_11 + 4'd7;
logic [31:0] bias_add_12;
assign bias_add_12 = conv_mac_12 + 3'd3;
logic [31:0] bias_add_13;
assign bias_add_13 = conv_mac_13 + 6'd24;
logic [31:0] bias_add_14;
assign bias_add_14 = conv_mac_14 + 5'd15;
logic [31:0] bias_add_15;
assign bias_add_15 = conv_mac_15 + 6'd17;
logic [31:0] bias_add_16;
assign bias_add_16 = conv_mac_16 + 6'd28;
logic [31:0] bias_add_17;
assign bias_add_17 = conv_mac_17 + 6'd19;
logic [31:0] bias_add_18;
assign bias_add_18 = conv_mac_18 + 6'd23;
logic [31:0] bias_add_19;
assign bias_add_19 = conv_mac_19 + 6'd21;
logic [31:0] bias_add_20;
assign bias_add_20 = conv_mac_20 + 6'd24;
logic [31:0] bias_add_21;
assign bias_add_21 = conv_mac_21 + 4'd7;
logic [31:0] bias_add_22;
assign bias_add_22 = conv_mac_22 + 5'd10;
logic [31:0] bias_add_23;
assign bias_add_23 = conv_mac_23 - 4'd4;
logic [31:0] bias_add_24;
assign bias_add_24 = conv_mac_24 - 6'd24;
logic [31:0] bias_add_25;
assign bias_add_25 = conv_mac_25 + 6'd16;
logic [31:0] bias_add_26;
assign bias_add_26 = conv_mac_26 + 6'd20;
logic [31:0] bias_add_27;
assign bias_add_27 = conv_mac_27 + 5'd11;
logic [31:0] bias_add_28;
assign bias_add_28 = conv_mac_28 + 7'd52;
logic [31:0] bias_add_29;
assign bias_add_29 = conv_mac_29 + 5'd11;
logic [31:0] bias_add_30;
assign bias_add_30 = conv_mac_30 + 6'd23;
logic [31:0] bias_add_31;
assign bias_add_31 = conv_mac_31 + 6'd19;

logic [7:0] relu_0;
assign relu_0[7:0] = (bias_add_0[31]==0) ? ((bias_add_0<3'd6) ? {{bias_add_0[31],bias_add_0[10:4]}} :'d6) : '0;
logic [7:0] relu_1;
assign relu_1[7:0] = (bias_add_1[31]==0) ? ((bias_add_1<3'd6) ? {{bias_add_1[31],bias_add_1[10:4]}} :'d6) : '0;
logic [7:0] relu_2;
assign relu_2[7:0] = (bias_add_2[31]==0) ? ((bias_add_2<3'd6) ? {{bias_add_2[31],bias_add_2[10:4]}} :'d6) : '0;
logic [7:0] relu_3;
assign relu_3[7:0] = (bias_add_3[31]==0) ? ((bias_add_3<3'd6) ? {{bias_add_3[31],bias_add_3[10:4]}} :'d6) : '0;
logic [7:0] relu_4;
assign relu_4[7:0] = (bias_add_4[31]==0) ? ((bias_add_4<3'd6) ? {{bias_add_4[31],bias_add_4[10:4]}} :'d6) : '0;
logic [7:0] relu_5;
assign relu_5[7:0] = (bias_add_5[31]==0) ? ((bias_add_5<3'd6) ? {{bias_add_5[31],bias_add_5[10:4]}} :'d6) : '0;
logic [7:0] relu_6;
assign relu_6[7:0] = (bias_add_6[31]==0) ? ((bias_add_6<3'd6) ? {{bias_add_6[31],bias_add_6[10:4]}} :'d6) : '0;
logic [7:0] relu_7;
assign relu_7[7:0] = (bias_add_7[31]==0) ? ((bias_add_7<3'd6) ? {{bias_add_7[31],bias_add_7[10:4]}} :'d6) : '0;
logic [7:0] relu_8;
assign relu_8[7:0] = (bias_add_8[31]==0) ? ((bias_add_8<3'd6) ? {{bias_add_8[31],bias_add_8[10:4]}} :'d6) : '0;
logic [7:0] relu_9;
assign relu_9[7:0] = (bias_add_9[31]==0) ? ((bias_add_9<3'd6) ? {{bias_add_9[31],bias_add_9[10:4]}} :'d6) : '0;
logic [7:0] relu_10;
assign relu_10[7:0] = (bias_add_10[31]==0) ? ((bias_add_10<3'd6) ? {{bias_add_10[31],bias_add_10[10:4]}} :'d6) : '0;
logic [7:0] relu_11;
assign relu_11[7:0] = (bias_add_11[31]==0) ? ((bias_add_11<3'd6) ? {{bias_add_11[31],bias_add_11[10:4]}} :'d6) : '0;
logic [7:0] relu_12;
assign relu_12[7:0] = (bias_add_12[31]==0) ? ((bias_add_12<3'd6) ? {{bias_add_12[31],bias_add_12[10:4]}} :'d6) : '0;
logic [7:0] relu_13;
assign relu_13[7:0] = (bias_add_13[31]==0) ? ((bias_add_13<3'd6) ? {{bias_add_13[31],bias_add_13[10:4]}} :'d6) : '0;
logic [7:0] relu_14;
assign relu_14[7:0] = (bias_add_14[31]==0) ? ((bias_add_14<3'd6) ? {{bias_add_14[31],bias_add_14[10:4]}} :'d6) : '0;
logic [7:0] relu_15;
assign relu_15[7:0] = (bias_add_15[31]==0) ? ((bias_add_15<3'd6) ? {{bias_add_15[31],bias_add_15[10:4]}} :'d6) : '0;
logic [7:0] relu_16;
assign relu_16[7:0] = (bias_add_16[31]==0) ? ((bias_add_16<3'd6) ? {{bias_add_16[31],bias_add_16[10:4]}} :'d6) : '0;
logic [7:0] relu_17;
assign relu_17[7:0] = (bias_add_17[31]==0) ? ((bias_add_17<3'd6) ? {{bias_add_17[31],bias_add_17[10:4]}} :'d6) : '0;
logic [7:0] relu_18;
assign relu_18[7:0] = (bias_add_18[31]==0) ? ((bias_add_18<3'd6) ? {{bias_add_18[31],bias_add_18[10:4]}} :'d6) : '0;
logic [7:0] relu_19;
assign relu_19[7:0] = (bias_add_19[31]==0) ? ((bias_add_19<3'd6) ? {{bias_add_19[31],bias_add_19[10:4]}} :'d6) : '0;
logic [7:0] relu_20;
assign relu_20[7:0] = (bias_add_20[31]==0) ? ((bias_add_20<3'd6) ? {{bias_add_20[31],bias_add_20[10:4]}} :'d6) : '0;
logic [7:0] relu_21;
assign relu_21[7:0] = (bias_add_21[31]==0) ? ((bias_add_21<3'd6) ? {{bias_add_21[31],bias_add_21[10:4]}} :'d6) : '0;
logic [7:0] relu_22;
assign relu_22[7:0] = (bias_add_22[31]==0) ? ((bias_add_22<3'd6) ? {{bias_add_22[31],bias_add_22[10:4]}} :'d6) : '0;
logic [7:0] relu_23;
assign relu_23[7:0] = (bias_add_23[31]==0) ? ((bias_add_23<3'd6) ? {{bias_add_23[31],bias_add_23[10:4]}} :'d6) : '0;
logic [7:0] relu_24;
assign relu_24[7:0] = (bias_add_24[31]==0) ? ((bias_add_24<3'd6) ? {{bias_add_24[31],bias_add_24[10:4]}} :'d6) : '0;
logic [7:0] relu_25;
assign relu_25[7:0] = (bias_add_25[31]==0) ? ((bias_add_25<3'd6) ? {{bias_add_25[31],bias_add_25[10:4]}} :'d6) : '0;
logic [7:0] relu_26;
assign relu_26[7:0] = (bias_add_26[31]==0) ? ((bias_add_26<3'd6) ? {{bias_add_26[31],bias_add_26[10:4]}} :'d6) : '0;
logic [7:0] relu_27;
assign relu_27[7:0] = (bias_add_27[31]==0) ? ((bias_add_27<3'd6) ? {{bias_add_27[31],bias_add_27[10:4]}} :'d6) : '0;
logic [7:0] relu_28;
assign relu_28[7:0] = (bias_add_28[31]==0) ? ((bias_add_28<3'd6) ? {{bias_add_28[31],bias_add_28[10:4]}} :'d6) : '0;
logic [7:0] relu_29;
assign relu_29[7:0] = (bias_add_29[31]==0) ? ((bias_add_29<3'd6) ? {{bias_add_29[31],bias_add_29[10:4]}} :'d6) : '0;
logic [7:0] relu_30;
assign relu_30[7:0] = (bias_add_30[31]==0) ? ((bias_add_30<3'd6) ? {{bias_add_30[31],bias_add_30[10:4]}} :'d6) : '0;
logic [7:0] relu_31;
assign relu_31[7:0] = (bias_add_31[31]==0) ? ((bias_add_31<3'd6) ? {{bias_add_31[31],bias_add_31[10:4]}} :'d6) : '0;

assign output_act = {
	relu_31,
	relu_30,
	relu_29,
	relu_28,
	relu_27,
	relu_26,
	relu_25,
	relu_24,
	relu_23,
	relu_22,
	relu_21,
	relu_20,
	relu_19,
	relu_18,
	relu_17,
	relu_16,
	relu_15,
	relu_14,
	relu_13,
	relu_12,
	relu_11,
	relu_10,
	relu_9,
	relu_8,
	relu_7,
	relu_6,
	relu_5,
	relu_4,
	relu_3,
	relu_2,
	relu_1,
	relu_0
};

endmodule
module conv5_pw (
    input logic clk,
    input logic rstn,
    input logic valid,
    input logic [256-1:0] input_act,
    output logic [256-1:0] output_act,
    output logic ready
);
logic we;
logic [8:0] zero_number; 
assign zero_number = 9'd0; 
//1
logic [256-1:0] input_act_ff ;
always_ff @(posedge clk) begin
    if (rstn == 0) begin
        input_act_ff <= '0;
      //  ready <= '0;
    end
    else begin
        input_act_ff <= input_act;
     //   ready <= valid;
    end
end
logic [7:0] input_fmap_0;
assign input_fmap_0 = input_act_ff[7:0];
logic [7:0] input_fmap_1;
assign input_fmap_1 = input_act_ff[15:8];
logic [7:0] input_fmap_2;
assign input_fmap_2 = input_act_ff[23:16];
logic [7:0] input_fmap_3;
assign input_fmap_3 = input_act_ff[31:24];
logic [7:0] input_fmap_4;
assign input_fmap_4 = input_act_ff[39:32];
logic [7:0] input_fmap_5;
assign input_fmap_5 = input_act_ff[47:40];
logic [7:0] input_fmap_6;
assign input_fmap_6 = input_act_ff[55:48];
logic [7:0] input_fmap_7;
assign input_fmap_7 = input_act_ff[63:56];
logic [7:0] input_fmap_8;
assign input_fmap_8 = input_act_ff[71:64];
logic [7:0] input_fmap_9;
assign input_fmap_9 = input_act_ff[79:72];
logic [7:0] input_fmap_10;
assign input_fmap_10 = input_act_ff[87:80];
logic [7:0] input_fmap_11;
assign input_fmap_11 = input_act_ff[95:88];
logic [7:0] input_fmap_12;
assign input_fmap_12 = input_act_ff[103:96];
logic [7:0] input_fmap_13;
assign input_fmap_13 = input_act_ff[111:104];
logic [7:0] input_fmap_14;
assign input_fmap_14 = input_act_ff[119:112];
logic [7:0] input_fmap_15;
assign input_fmap_15 = input_act_ff[127:120];
logic [7:0] input_fmap_16;
assign input_fmap_16 = input_act_ff[135:128];
logic [7:0] input_fmap_17;
assign input_fmap_17 = input_act_ff[143:136];
logic [7:0] input_fmap_18;
assign input_fmap_18 = input_act_ff[151:144];
logic [7:0] input_fmap_19;
assign input_fmap_19 = input_act_ff[159:152];
logic [7:0] input_fmap_20;
assign input_fmap_20 = input_act_ff[167:160];
logic [7:0] input_fmap_21;
assign input_fmap_21 = input_act_ff[175:168];
logic [7:0] input_fmap_22;
assign input_fmap_22 = input_act_ff[183:176];
logic [7:0] input_fmap_23;
assign input_fmap_23 = input_act_ff[191:184];
logic [7:0] input_fmap_24;
assign input_fmap_24 = input_act_ff[199:192];
logic [7:0] input_fmap_25;
assign input_fmap_25 = input_act_ff[207:200];
logic [7:0] input_fmap_26;
assign input_fmap_26 = input_act_ff[215:208];
logic [7:0] input_fmap_27;
assign input_fmap_27 = input_act_ff[223:216];
logic [7:0] input_fmap_28;
assign input_fmap_28 = input_act_ff[231:224];
logic [7:0] input_fmap_29;
assign input_fmap_29 = input_act_ff[239:232];
logic [7:0] input_fmap_30;
assign input_fmap_30 = input_act_ff[247:240];
logic [7:0] input_fmap_31;
assign input_fmap_31 = input_act_ff[255:248];

logic [10-1:0] O0_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O0_I0_R0_C01_rom_inst (.q(O0_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I0_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O0_I0_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O0_I0_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O0_I0_R0_C01_rom_inst (.q(O0_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [11-1:0] O0_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O0_I2_R0_C02_rom_inst (.q(O0_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I2_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O0_I2_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O0_I2_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O0_I2_R0_C02_rom_inst (.q(O0_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [10-1:0] O0_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O0_I4_R0_C01_rom_inst (.q(O0_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I4_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O0_I4_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O0_I4_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O0_I4_R0_C01_rom_inst (.q(O0_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [10-1:0] O0_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O0_I5_R0_C01_rom_inst (.q(O0_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I5_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O0_I5_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O0_I5_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O0_I5_R0_C01_rom_inst (.q(O0_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [10-1:0] O0_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O0_I6_R0_C01_rom_inst (.q(O0_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I6_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O0_I6_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O0_I6_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O0_I6_R0_C01_rom_inst (.q(O0_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [10-1:0] O0_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O0_I7_R0_C01_rom_inst (.q(O0_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I7_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O0_I7_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O0_I7_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O0_I7_R0_C01_rom_inst (.q(O0_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [10-1:0] O0_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O0_I8_R0_C01_rom_inst (.q(O0_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I8_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O0_I8_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O0_I8_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O0_I8_R0_C01_rom_inst (.q(O0_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [10-1:0] O0_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O0_I9_R0_C01_rom_inst (.q(O0_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I9_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O0_I9_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O0_I9_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O0_I9_R0_C01_rom_inst (.q(O0_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [10-1:0] O0_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O0_I11_R0_C01_rom_inst (.q(O0_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I11_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O0_I11_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O0_I11_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O0_I11_R0_C01_rom_inst (.q(O0_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [10-1:0] O0_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O0_I13_R0_C01_rom_inst (.q(O0_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I13_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O0_I13_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O0_I13_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O0_I13_R0_C01_rom_inst (.q(O0_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [10-1:0] O0_I17_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O0_I17_R0_C01_rom_inst (.q(O0_I17_R0_C0_SM1 ),.address(input_fmap_17[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I17_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O0_I17_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O0_I17_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O0_I17_R0_C01_rom_inst (.q(O0_I17_R0_C0_SM1 ),.address(input_fmap_17[7:0]),.clock  (clk));
logic [10-1:0] O0_I19_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O0_I19_R0_C01_rom_inst (.q(O0_I19_R0_C0_SM1 ),.address(input_fmap_19[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I19_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O0_I19_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O0_I19_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O0_I19_R0_C01_rom_inst (.q(O0_I19_R0_C0_SM1 ),.address(input_fmap_19[7:0]),.clock  (clk));
logic [11-1:0] O0_I20_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O0_I20_R0_C03_rom_inst (.q(O0_I20_R0_C0_SM1 ),.address(input_fmap_20[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I20_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O0_I20_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O0_I20_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O0_I20_R0_C03_rom_inst (.q(O0_I20_R0_C0_SM1 ),.address(input_fmap_20[7:0]),.clock  (clk));
logic [10-1:0] O0_I23_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O0_I23_R0_C01_rom_inst (.q(O0_I23_R0_C0_SM1 ),.address(input_fmap_23[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I23_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O0_I23_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O0_I23_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O0_I23_R0_C01_rom_inst (.q(O0_I23_R0_C0_SM1 ),.address(input_fmap_23[7:0]),.clock  (clk));
logic [10-1:0] O0_I25_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O0_I25_R0_C01_rom_inst (.q(O0_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I25_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O0_I25_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O0_I25_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O0_I25_R0_C01_rom_inst (.q(O0_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clock  (clk));
logic [10-1:0] O0_I29_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O0_I29_R0_C01_rom_inst (.q(O0_I29_R0_C0_SM1 ),.address(input_fmap_29[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I29_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O0_I29_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O0_I29_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O0_I29_R0_C01_rom_inst (.q(O0_I29_R0_C0_SM1 ),.address(input_fmap_29[7:0]),.clock  (clk));
logic [10-1:0] O0_I31_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O0_I31_R0_C01_rom_inst (.q(O0_I31_R0_C0_SM1 ),.address(input_fmap_31[7:0]),.clk(clk),.d(0),.we(0));
//assign O0_I31_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O0_I31_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O0_I31_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O0_I31_R0_C01_rom_inst (.q(O0_I31_R0_C0_SM1 ),.address(input_fmap_31[7:0]),.clock  (clk));
logic [10-1:0] O1_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O1_I9_R0_C01_rom_inst (.q(O1_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I9_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O1_I9_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O1_I9_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O1_I9_R0_C01_rom_inst (.q(O1_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [11-1:0] O1_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O1_I11_R0_C02_rom_inst (.q(O1_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I11_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O1_I11_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O1_I11_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O1_I11_R0_C02_rom_inst (.q(O1_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [10-1:0] O1_I23_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O1_I23_R0_C01_rom_inst (.q(O1_I23_R0_C0_SM1 ),.address(input_fmap_23[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I23_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O1_I23_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O1_I23_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O1_I23_R0_C01_rom_inst (.q(O1_I23_R0_C0_SM1 ),.address(input_fmap_23[7:0]),.clock  (clk));
logic [10-1:0] O1_I26_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O1_I26_R0_C01_rom_inst (.q(O1_I26_R0_C0_SM1 ),.address(input_fmap_26[7:0]),.clk(clk),.d(0),.we(0));
//assign O1_I26_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O1_I26_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O1_I26_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O1_I26_R0_C01_rom_inst (.q(O1_I26_R0_C0_SM1 ),.address(input_fmap_26[7:0]),.clock  (clk));
logic [10-1:0] O2_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O2_I3_R0_C01_rom_inst (.q(O2_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O2_I3_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O2_I3_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O2_I3_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O2_I3_R0_C01_rom_inst (.q(O2_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [10-1:0] O2_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O2_I7_R0_C01_rom_inst (.q(O2_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O2_I7_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O2_I7_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O2_I7_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O2_I7_R0_C01_rom_inst (.q(O2_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [10-1:0] O2_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O2_I9_R0_C01_rom_inst (.q(O2_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O2_I9_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O2_I9_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O2_I9_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O2_I9_R0_C01_rom_inst (.q(O2_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [11-1:0] O2_I10_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O2_I10_R0_C03_rom_inst (.q(O2_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clk(clk),.d(0),.we(0));
//assign O2_I10_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O2_I10_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O2_I10_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O2_I10_R0_C03_rom_inst (.q(O2_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clock  (clk));
logic [10-1:0] O2_I14_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O2_I14_R0_C01_rom_inst (.q(O2_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clk(clk),.d(0),.we(0));
//assign O2_I14_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O2_I14_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O2_I14_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O2_I14_R0_C01_rom_inst (.q(O2_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clock  (clk));
logic [10-1:0] O2_I23_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O2_I23_R0_C01_rom_inst (.q(O2_I23_R0_C0_SM1 ),.address(input_fmap_23[7:0]),.clk(clk),.d(0),.we(0));
//assign O2_I23_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O2_I23_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O2_I23_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O2_I23_R0_C01_rom_inst (.q(O2_I23_R0_C0_SM1 ),.address(input_fmap_23[7:0]),.clock  (clk));
logic [10-1:0] O2_I25_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O2_I25_R0_C01_rom_inst (.q(O2_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clk(clk),.d(0),.we(0));
//assign O2_I25_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O2_I25_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O2_I25_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O2_I25_R0_C01_rom_inst (.q(O2_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clock  (clk));
logic [11-1:0] O2_I28_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O2_I28_R0_C02_rom_inst (.q(O2_I28_R0_C0_SM1 ),.address(input_fmap_28[7:0]),.clk(clk),.d(0),.we(0));
//assign O2_I28_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O2_I28_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O2_I28_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O2_I28_R0_C02_rom_inst (.q(O2_I28_R0_C0_SM1 ),.address(input_fmap_28[7:0]),.clock  (clk));
logic [11-1:0] O2_I29_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O2_I29_R0_C02_rom_inst (.q(O2_I29_R0_C0_SM1 ),.address(input_fmap_29[7:0]),.clk(clk),.d(0),.we(0));
//assign O2_I29_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O2_I29_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O2_I29_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O2_I29_R0_C02_rom_inst (.q(O2_I29_R0_C0_SM1 ),.address(input_fmap_29[7:0]),.clock  (clk));
logic [10-1:0] O3_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O3_I1_R0_C01_rom_inst (.q(O3_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I1_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O3_I1_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O3_I1_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O3_I1_R0_C01_rom_inst (.q(O3_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [10-1:0] O3_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O3_I2_R0_C01_rom_inst (.q(O3_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O3_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O3_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O3_I2_R0_C01_rom_inst (.q(O3_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [11-1:0] O3_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O3_I3_R0_C03_rom_inst (.q(O3_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I3_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O3_I3_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O3_I3_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O3_I3_R0_C03_rom_inst (.q(O3_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [10-1:0] O3_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O3_I5_R0_C01_rom_inst (.q(O3_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I5_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O3_I5_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O3_I5_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O3_I5_R0_C01_rom_inst (.q(O3_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [10-1:0] O3_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O3_I6_R0_C01_rom_inst (.q(O3_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I6_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O3_I6_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O3_I6_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O3_I6_R0_C01_rom_inst (.q(O3_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [10-1:0] O3_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O3_I7_R0_C01_rom_inst (.q(O3_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I7_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O3_I7_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O3_I7_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O3_I7_R0_C01_rom_inst (.q(O3_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [10-1:0] O3_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O3_I8_R0_C01_rom_inst (.q(O3_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I8_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O3_I8_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O3_I8_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O3_I8_R0_C01_rom_inst (.q(O3_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [10-1:0] O3_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O3_I9_R0_C01_rom_inst (.q(O3_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I9_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O3_I9_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O3_I9_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O3_I9_R0_C01_rom_inst (.q(O3_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [12-1:0] O3_I10_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_pw_O3_I10_R0_C04_rom_inst (.q(O3_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I10_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O3_I10_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O3_I10_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_pw_O3_I10_R0_C04_rom_inst (.q(O3_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clock  (clk));
logic [10-1:0] O3_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O3_I12_R0_C01_rom_inst (.q(O3_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I12_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O3_I12_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O3_I12_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O3_I12_R0_C01_rom_inst (.q(O3_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [10-1:0] O3_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O3_I13_R0_C01_rom_inst (.q(O3_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I13_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O3_I13_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O3_I13_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O3_I13_R0_C01_rom_inst (.q(O3_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [12-1:0] O3_I14_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_pw_O3_I14_R0_C07_rom_inst (.q(O3_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I14_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O3_I14_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O3_I14_R0_C07_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_pw_O3_I14_R0_C07_rom_inst (.q(O3_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clock  (clk));
logic [10-1:0] O3_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O3_I15_R0_C01_rom_inst (.q(O3_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I15_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O3_I15_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O3_I15_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O3_I15_R0_C01_rom_inst (.q(O3_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [10-1:0] O3_I16_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O3_I16_R0_C01_rom_inst (.q(O3_I16_R0_C0_SM1 ),.address(input_fmap_16[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I16_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O3_I16_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O3_I16_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O3_I16_R0_C01_rom_inst (.q(O3_I16_R0_C0_SM1 ),.address(input_fmap_16[7:0]),.clock  (clk));
logic [12-1:0] O3_I18_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_pw_O3_I18_R0_C04_rom_inst (.q(O3_I18_R0_C0_SM1 ),.address(input_fmap_18[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I18_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O3_I18_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O3_I18_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_pw_O3_I18_R0_C04_rom_inst (.q(O3_I18_R0_C0_SM1 ),.address(input_fmap_18[7:0]),.clock  (clk));
logic [10-1:0] O3_I21_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O3_I21_R0_C01_rom_inst (.q(O3_I21_R0_C0_SM1 ),.address(input_fmap_21[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I21_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O3_I21_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O3_I21_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O3_I21_R0_C01_rom_inst (.q(O3_I21_R0_C0_SM1 ),.address(input_fmap_21[7:0]),.clock  (clk));
logic [11-1:0] O3_I22_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O3_I22_R0_C02_rom_inst (.q(O3_I22_R0_C0_SM1 ),.address(input_fmap_22[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I22_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O3_I22_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O3_I22_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O3_I22_R0_C02_rom_inst (.q(O3_I22_R0_C0_SM1 ),.address(input_fmap_22[7:0]),.clock  (clk));
logic [10-1:0] O3_I23_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O3_I23_R0_C01_rom_inst (.q(O3_I23_R0_C0_SM1 ),.address(input_fmap_23[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I23_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O3_I23_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O3_I23_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O3_I23_R0_C01_rom_inst (.q(O3_I23_R0_C0_SM1 ),.address(input_fmap_23[7:0]),.clock  (clk));
logic [10-1:0] O3_I24_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O3_I24_R0_C01_rom_inst (.q(O3_I24_R0_C0_SM1 ),.address(input_fmap_24[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I24_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O3_I24_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O3_I24_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O3_I24_R0_C01_rom_inst (.q(O3_I24_R0_C0_SM1 ),.address(input_fmap_24[7:0]),.clock  (clk));
logic [10-1:0] O3_I25_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O3_I25_R0_C01_rom_inst (.q(O3_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I25_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O3_I25_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O3_I25_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O3_I25_R0_C01_rom_inst (.q(O3_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clock  (clk));
logic [11-1:0] O3_I29_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O3_I29_R0_C03_rom_inst (.q(O3_I29_R0_C0_SM1 ),.address(input_fmap_29[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I29_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O3_I29_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O3_I29_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O3_I29_R0_C03_rom_inst (.q(O3_I29_R0_C0_SM1 ),.address(input_fmap_29[7:0]),.clock  (clk));
logic [10-1:0] O3_I30_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O3_I30_R0_C01_rom_inst (.q(O3_I30_R0_C0_SM1 ),.address(input_fmap_30[7:0]),.clk(clk),.d(0),.we(0));
//assign O3_I30_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O3_I30_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O3_I30_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O3_I30_R0_C01_rom_inst (.q(O3_I30_R0_C0_SM1 ),.address(input_fmap_30[7:0]),.clock  (clk));
logic [10-1:0] O4_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O4_I0_R0_C01_rom_inst (.q(O4_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I0_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I0_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O4_I0_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O4_I0_R0_C01_rom_inst (.q(O4_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [10-1:0] O4_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O4_I3_R0_C01_rom_inst (.q(O4_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I3_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I3_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O4_I3_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O4_I3_R0_C01_rom_inst (.q(O4_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [10-1:0] O4_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O4_I4_R0_C01_rom_inst (.q(O4_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I4_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I4_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O4_I4_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O4_I4_R0_C01_rom_inst (.q(O4_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [10-1:0] O4_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O4_I5_R0_C01_rom_inst (.q(O4_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I5_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I5_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O4_I5_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O4_I5_R0_C01_rom_inst (.q(O4_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [10-1:0] O4_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O4_I8_R0_C01_rom_inst (.q(O4_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I8_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I8_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O4_I8_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O4_I8_R0_C01_rom_inst (.q(O4_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [10-1:0] O4_I10_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O4_I10_R0_C01_rom_inst (.q(O4_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I10_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I10_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O4_I10_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O4_I10_R0_C01_rom_inst (.q(O4_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clock  (clk));
logic [10-1:0] O4_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O4_I11_R0_C01_rom_inst (.q(O4_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I11_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I11_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O4_I11_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O4_I11_R0_C01_rom_inst (.q(O4_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [10-1:0] O4_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O4_I12_R0_C01_rom_inst (.q(O4_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I12_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I12_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O4_I12_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O4_I12_R0_C01_rom_inst (.q(O4_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [10-1:0] O4_I14_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O4_I14_R0_C01_rom_inst (.q(O4_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I14_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I14_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O4_I14_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O4_I14_R0_C01_rom_inst (.q(O4_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clock  (clk));
logic [10-1:0] O4_I16_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O4_I16_R0_C01_rom_inst (.q(O4_I16_R0_C0_SM1 ),.address(input_fmap_16[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I16_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I16_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O4_I16_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O4_I16_R0_C01_rom_inst (.q(O4_I16_R0_C0_SM1 ),.address(input_fmap_16[7:0]),.clock  (clk));
logic [10-1:0] O4_I17_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O4_I17_R0_C01_rom_inst (.q(O4_I17_R0_C0_SM1 ),.address(input_fmap_17[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I17_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I17_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O4_I17_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O4_I17_R0_C01_rom_inst (.q(O4_I17_R0_C0_SM1 ),.address(input_fmap_17[7:0]),.clock  (clk));
logic [10-1:0] O4_I18_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O4_I18_R0_C01_rom_inst (.q(O4_I18_R0_C0_SM1 ),.address(input_fmap_18[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I18_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I18_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O4_I18_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O4_I18_R0_C01_rom_inst (.q(O4_I18_R0_C0_SM1 ),.address(input_fmap_18[7:0]),.clock  (clk));
logic [11-1:0] O4_I19_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O4_I19_R0_C02_rom_inst (.q(O4_I19_R0_C0_SM1 ),.address(input_fmap_19[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I19_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O4_I19_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O4_I19_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O4_I19_R0_C02_rom_inst (.q(O4_I19_R0_C0_SM1 ),.address(input_fmap_19[7:0]),.clock  (clk));
logic [10-1:0] O4_I20_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O4_I20_R0_C01_rom_inst (.q(O4_I20_R0_C0_SM1 ),.address(input_fmap_20[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I20_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I20_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O4_I20_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O4_I20_R0_C01_rom_inst (.q(O4_I20_R0_C0_SM1 ),.address(input_fmap_20[7:0]),.clock  (clk));
logic [10-1:0] O4_I21_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O4_I21_R0_C01_rom_inst (.q(O4_I21_R0_C0_SM1 ),.address(input_fmap_21[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I21_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I21_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O4_I21_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O4_I21_R0_C01_rom_inst (.q(O4_I21_R0_C0_SM1 ),.address(input_fmap_21[7:0]),.clock  (clk));
logic [12-1:0] O4_I25_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_pw_O4_I25_R0_C04_rom_inst (.q(O4_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I25_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O4_I25_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O4_I25_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_pw_O4_I25_R0_C04_rom_inst (.q(O4_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clock  (clk));
logic [11-1:0] O4_I26_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O4_I26_R0_C02_rom_inst (.q(O4_I26_R0_C0_SM1 ),.address(input_fmap_26[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I26_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O4_I26_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O4_I26_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O4_I26_R0_C02_rom_inst (.q(O4_I26_R0_C0_SM1 ),.address(input_fmap_26[7:0]),.clock  (clk));
logic [10-1:0] O4_I27_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O4_I27_R0_C01_rom_inst (.q(O4_I27_R0_C0_SM1 ),.address(input_fmap_27[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I27_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I27_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O4_I27_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O4_I27_R0_C01_rom_inst (.q(O4_I27_R0_C0_SM1 ),.address(input_fmap_27[7:0]),.clock  (clk));
logic [11-1:0] O4_I29_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O4_I29_R0_C02_rom_inst (.q(O4_I29_R0_C0_SM1 ),.address(input_fmap_29[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I29_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O4_I29_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O4_I29_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O4_I29_R0_C02_rom_inst (.q(O4_I29_R0_C0_SM1 ),.address(input_fmap_29[7:0]),.clock  (clk));
logic [10-1:0] O4_I30_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O4_I30_R0_C01_rom_inst (.q(O4_I30_R0_C0_SM1 ),.address(input_fmap_30[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I30_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I30_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O4_I30_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O4_I30_R0_C01_rom_inst (.q(O4_I30_R0_C0_SM1 ),.address(input_fmap_30[7:0]),.clock  (clk));
logic [10-1:0] O4_I31_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O4_I31_R0_C01_rom_inst (.q(O4_I31_R0_C0_SM1 ),.address(input_fmap_31[7:0]),.clk(clk),.d(0),.we(0));
//assign O4_I31_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O4_I31_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O4_I31_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O4_I31_R0_C01_rom_inst (.q(O4_I31_R0_C0_SM1 ),.address(input_fmap_31[7:0]),.clock  (clk));
logic [10-1:0] O5_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O5_I0_R0_C01_rom_inst (.q(O5_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I0_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I0_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O5_I0_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O5_I0_R0_C01_rom_inst (.q(O5_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [10-1:0] O5_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O5_I1_R0_C01_rom_inst (.q(O5_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I1_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I1_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O5_I1_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O5_I1_R0_C01_rom_inst (.q(O5_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [12-1:0] O5_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_pw_O5_I2_R0_C04_rom_inst (.q(O5_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I2_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O5_I2_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O5_I2_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_pw_O5_I2_R0_C04_rom_inst (.q(O5_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [11-1:0] O5_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O5_I5_R0_C03_rom_inst (.q(O5_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I5_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O5_I5_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O5_I5_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O5_I5_R0_C03_rom_inst (.q(O5_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [10-1:0] O5_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O5_I9_R0_C01_rom_inst (.q(O5_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I9_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I9_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O5_I9_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O5_I9_R0_C01_rom_inst (.q(O5_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [11-1:0] O5_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O5_I12_R0_C03_rom_inst (.q(O5_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I12_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O5_I12_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O5_I12_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O5_I12_R0_C03_rom_inst (.q(O5_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [10-1:0] O5_I19_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O5_I19_R0_C01_rom_inst (.q(O5_I19_R0_C0_SM1 ),.address(input_fmap_19[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I19_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I19_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O5_I19_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O5_I19_R0_C01_rom_inst (.q(O5_I19_R0_C0_SM1 ),.address(input_fmap_19[7:0]),.clock  (clk));
logic [10-1:0] O5_I20_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O5_I20_R0_C01_rom_inst (.q(O5_I20_R0_C0_SM1 ),.address(input_fmap_20[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I20_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I20_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O5_I20_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O5_I20_R0_C01_rom_inst (.q(O5_I20_R0_C0_SM1 ),.address(input_fmap_20[7:0]),.clock  (clk));
logic [10-1:0] O5_I23_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O5_I23_R0_C01_rom_inst (.q(O5_I23_R0_C0_SM1 ),.address(input_fmap_23[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I23_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I23_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O5_I23_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O5_I23_R0_C01_rom_inst (.q(O5_I23_R0_C0_SM1 ),.address(input_fmap_23[7:0]),.clock  (clk));
logic [10-1:0] O5_I24_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O5_I24_R0_C01_rom_inst (.q(O5_I24_R0_C0_SM1 ),.address(input_fmap_24[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I24_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I24_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O5_I24_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O5_I24_R0_C01_rom_inst (.q(O5_I24_R0_C0_SM1 ),.address(input_fmap_24[7:0]),.clock  (clk));
logic [10-1:0] O5_I25_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O5_I25_R0_C01_rom_inst (.q(O5_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I25_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I25_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O5_I25_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O5_I25_R0_C01_rom_inst (.q(O5_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clock  (clk));
logic [11-1:0] O5_I28_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O5_I28_R0_C02_rom_inst (.q(O5_I28_R0_C0_SM1 ),.address(input_fmap_28[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I28_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O5_I28_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O5_I28_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O5_I28_R0_C02_rom_inst (.q(O5_I28_R0_C0_SM1 ),.address(input_fmap_28[7:0]),.clock  (clk));
logic [10-1:0] O5_I30_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O5_I30_R0_C01_rom_inst (.q(O5_I30_R0_C0_SM1 ),.address(input_fmap_30[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I30_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O5_I30_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O5_I30_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O5_I30_R0_C01_rom_inst (.q(O5_I30_R0_C0_SM1 ),.address(input_fmap_30[7:0]),.clock  (clk));
logic [11-1:0] O5_I31_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O5_I31_R0_C02_rom_inst (.q(O5_I31_R0_C0_SM1 ),.address(input_fmap_31[7:0]),.clk(clk),.d(0),.we(0));
//assign O5_I31_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O5_I31_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O5_I31_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O5_I31_R0_C02_rom_inst (.q(O5_I31_R0_C0_SM1 ),.address(input_fmap_31[7:0]),.clock  (clk));
logic [10-1:0] O6_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O6_I0_R0_C01_rom_inst (.q(O6_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I0_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O6_I0_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O6_I0_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O6_I0_R0_C01_rom_inst (.q(O6_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [10-1:0] O6_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O6_I1_R0_C01_rom_inst (.q(O6_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I1_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O6_I1_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O6_I1_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O6_I1_R0_C01_rom_inst (.q(O6_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [11-1:0] O6_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O6_I2_R0_C03_rom_inst (.q(O6_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I2_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O6_I2_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O6_I2_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O6_I2_R0_C03_rom_inst (.q(O6_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [11-1:0] O6_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O6_I4_R0_C02_rom_inst (.q(O6_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I4_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O6_I4_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O6_I4_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O6_I4_R0_C02_rom_inst (.q(O6_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [10-1:0] O6_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O6_I6_R0_C01_rom_inst (.q(O6_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I6_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O6_I6_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O6_I6_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O6_I6_R0_C01_rom_inst (.q(O6_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [12-1:0] O6_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_pw_O6_I7_R0_C04_rom_inst (.q(O6_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I7_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O6_I7_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O6_I7_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_pw_O6_I7_R0_C04_rom_inst (.q(O6_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [11-1:0] O6_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O6_I8_R0_C02_rom_inst (.q(O6_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I8_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O6_I8_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O6_I8_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O6_I8_R0_C02_rom_inst (.q(O6_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [11-1:0] O6_I10_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O6_I10_R0_C02_rom_inst (.q(O6_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I10_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O6_I10_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O6_I10_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O6_I10_R0_C02_rom_inst (.q(O6_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clock  (clk));
logic [10-1:0] O6_I14_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O6_I14_R0_C01_rom_inst (.q(O6_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I14_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O6_I14_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O6_I14_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O6_I14_R0_C01_rom_inst (.q(O6_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clock  (clk));
logic [11-1:0] O6_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O6_I15_R0_C02_rom_inst (.q(O6_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I15_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O6_I15_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O6_I15_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O6_I15_R0_C02_rom_inst (.q(O6_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [10-1:0] O6_I16_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O6_I16_R0_C01_rom_inst (.q(O6_I16_R0_C0_SM1 ),.address(input_fmap_16[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I16_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O6_I16_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O6_I16_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O6_I16_R0_C01_rom_inst (.q(O6_I16_R0_C0_SM1 ),.address(input_fmap_16[7:0]),.clock  (clk));
logic [12-1:0] O6_I17_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_pw_O6_I17_R0_C05_rom_inst (.q(O6_I17_R0_C0_SM1 ),.address(input_fmap_17[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I17_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O6_I17_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O6_I17_R0_C05_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_pw_O6_I17_R0_C05_rom_inst (.q(O6_I17_R0_C0_SM1 ),.address(input_fmap_17[7:0]),.clock  (clk));
logic [11-1:0] O6_I19_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O6_I19_R0_C03_rom_inst (.q(O6_I19_R0_C0_SM1 ),.address(input_fmap_19[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I19_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O6_I19_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O6_I19_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O6_I19_R0_C03_rom_inst (.q(O6_I19_R0_C0_SM1 ),.address(input_fmap_19[7:0]),.clock  (clk));
logic [11-1:0] O6_I20_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O6_I20_R0_C03_rom_inst (.q(O6_I20_R0_C0_SM1 ),.address(input_fmap_20[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I20_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O6_I20_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O6_I20_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O6_I20_R0_C03_rom_inst (.q(O6_I20_R0_C0_SM1 ),.address(input_fmap_20[7:0]),.clock  (clk));
logic [12-1:0] O6_I21_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_pw_O6_I21_R0_C05_rom_inst (.q(O6_I21_R0_C0_SM1 ),.address(input_fmap_21[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I21_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O6_I21_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O6_I21_R0_C05_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_pw_O6_I21_R0_C05_rom_inst (.q(O6_I21_R0_C0_SM1 ),.address(input_fmap_21[7:0]),.clock  (clk));
logic [10-1:0] O6_I22_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O6_I22_R0_C01_rom_inst (.q(O6_I22_R0_C0_SM1 ),.address(input_fmap_22[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I22_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O6_I22_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O6_I22_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O6_I22_R0_C01_rom_inst (.q(O6_I22_R0_C0_SM1 ),.address(input_fmap_22[7:0]),.clock  (clk));
logic [10-1:0] O6_I23_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O6_I23_R0_C01_rom_inst (.q(O6_I23_R0_C0_SM1 ),.address(input_fmap_23[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I23_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O6_I23_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O6_I23_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O6_I23_R0_C01_rom_inst (.q(O6_I23_R0_C0_SM1 ),.address(input_fmap_23[7:0]),.clock  (clk));
logic [10-1:0] O6_I24_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O6_I24_R0_C01_rom_inst (.q(O6_I24_R0_C0_SM1 ),.address(input_fmap_24[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I24_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O6_I24_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O6_I24_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O6_I24_R0_C01_rom_inst (.q(O6_I24_R0_C0_SM1 ),.address(input_fmap_24[7:0]),.clock  (clk));
logic [11-1:0] O6_I25_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O6_I25_R0_C03_rom_inst (.q(O6_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I25_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O6_I25_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O6_I25_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O6_I25_R0_C03_rom_inst (.q(O6_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clock  (clk));
logic [11-1:0] O6_I26_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O6_I26_R0_C03_rom_inst (.q(O6_I26_R0_C0_SM1 ),.address(input_fmap_26[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I26_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O6_I26_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O6_I26_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O6_I26_R0_C03_rom_inst (.q(O6_I26_R0_C0_SM1 ),.address(input_fmap_26[7:0]),.clock  (clk));
logic [13-1:0] O6_I27_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(13),.INIT_FILE("deepfreeze_rom/deepfreeze_8_13.txt"))
    conv5_pw_O6_I27_R0_C010_rom_inst (.q(O6_I27_R0_C0_SM1 ),.address(input_fmap_27[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I27_R0_C0_SM1  = 13'h1234;
//always@(posedge clk) begin 
//O6_I27_R0_C0_SM1  <= 13'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O6_I27_R0_C010_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(13))
//    conv5_pw_O6_I27_R0_C010_rom_inst (.q(O6_I27_R0_C0_SM1 ),.address(input_fmap_27[7:0]),.clock  (clk));
logic [12-1:0] O6_I28_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_pw_O6_I28_R0_C04_rom_inst (.q(O6_I28_R0_C0_SM1 ),.address(input_fmap_28[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I28_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O6_I28_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O6_I28_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_pw_O6_I28_R0_C04_rom_inst (.q(O6_I28_R0_C0_SM1 ),.address(input_fmap_28[7:0]),.clock  (clk));
logic [11-1:0] O6_I29_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O6_I29_R0_C02_rom_inst (.q(O6_I29_R0_C0_SM1 ),.address(input_fmap_29[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I29_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O6_I29_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O6_I29_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O6_I29_R0_C02_rom_inst (.q(O6_I29_R0_C0_SM1 ),.address(input_fmap_29[7:0]),.clock  (clk));
logic [11-1:0] O6_I31_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O6_I31_R0_C02_rom_inst (.q(O6_I31_R0_C0_SM1 ),.address(input_fmap_31[7:0]),.clk(clk),.d(0),.we(0));
//assign O6_I31_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O6_I31_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O6_I31_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O6_I31_R0_C02_rom_inst (.q(O6_I31_R0_C0_SM1 ),.address(input_fmap_31[7:0]),.clock  (clk));
logic [10-1:0] O7_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O7_I3_R0_C01_rom_inst (.q(O7_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I3_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O7_I3_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O7_I3_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O7_I3_R0_C01_rom_inst (.q(O7_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [10-1:0] O7_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O7_I9_R0_C01_rom_inst (.q(O7_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I9_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O7_I9_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O7_I9_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O7_I9_R0_C01_rom_inst (.q(O7_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [11-1:0] O7_I14_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O7_I14_R0_C03_rom_inst (.q(O7_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I14_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O7_I14_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O7_I14_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O7_I14_R0_C03_rom_inst (.q(O7_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clock  (clk));
logic [11-1:0] O7_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O7_I15_R0_C02_rom_inst (.q(O7_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I15_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O7_I15_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O7_I15_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O7_I15_R0_C02_rom_inst (.q(O7_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [11-1:0] O7_I18_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O7_I18_R0_C02_rom_inst (.q(O7_I18_R0_C0_SM1 ),.address(input_fmap_18[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I18_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O7_I18_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O7_I18_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O7_I18_R0_C02_rom_inst (.q(O7_I18_R0_C0_SM1 ),.address(input_fmap_18[7:0]),.clock  (clk));
logic [10-1:0] O7_I23_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O7_I23_R0_C01_rom_inst (.q(O7_I23_R0_C0_SM1 ),.address(input_fmap_23[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I23_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O7_I23_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O7_I23_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O7_I23_R0_C01_rom_inst (.q(O7_I23_R0_C0_SM1 ),.address(input_fmap_23[7:0]),.clock  (clk));
logic [10-1:0] O7_I27_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O7_I27_R0_C01_rom_inst (.q(O7_I27_R0_C0_SM1 ),.address(input_fmap_27[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I27_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O7_I27_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O7_I27_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O7_I27_R0_C01_rom_inst (.q(O7_I27_R0_C0_SM1 ),.address(input_fmap_27[7:0]),.clock  (clk));
logic [10-1:0] O7_I28_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O7_I28_R0_C01_rom_inst (.q(O7_I28_R0_C0_SM1 ),.address(input_fmap_28[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I28_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O7_I28_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O7_I28_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O7_I28_R0_C01_rom_inst (.q(O7_I28_R0_C0_SM1 ),.address(input_fmap_28[7:0]),.clock  (clk));
logic [11-1:0] O7_I29_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O7_I29_R0_C02_rom_inst (.q(O7_I29_R0_C0_SM1 ),.address(input_fmap_29[7:0]),.clk(clk),.d(0),.we(0));
//assign O7_I29_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O7_I29_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O7_I29_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O7_I29_R0_C02_rom_inst (.q(O7_I29_R0_C0_SM1 ),.address(input_fmap_29[7:0]),.clock  (clk));
logic [10-1:0] O8_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O8_I2_R0_C01_rom_inst (.q(O8_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O8_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O8_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O8_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O8_I2_R0_C01_rom_inst (.q(O8_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [10-1:0] O8_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O8_I4_R0_C01_rom_inst (.q(O8_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O8_I4_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O8_I4_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O8_I4_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O8_I4_R0_C01_rom_inst (.q(O8_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [10-1:0] O8_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O8_I5_R0_C01_rom_inst (.q(O8_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O8_I5_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O8_I5_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O8_I5_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O8_I5_R0_C01_rom_inst (.q(O8_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [10-1:0] O8_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O8_I6_R0_C01_rom_inst (.q(O8_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O8_I6_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O8_I6_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O8_I6_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O8_I6_R0_C01_rom_inst (.q(O8_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [10-1:0] O8_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O8_I7_R0_C01_rom_inst (.q(O8_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O8_I7_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O8_I7_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O8_I7_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O8_I7_R0_C01_rom_inst (.q(O8_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [10-1:0] O8_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O8_I9_R0_C01_rom_inst (.q(O8_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O8_I9_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O8_I9_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O8_I9_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O8_I9_R0_C01_rom_inst (.q(O8_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [10-1:0] O8_I10_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O8_I10_R0_C01_rom_inst (.q(O8_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clk(clk),.d(0),.we(0));
//assign O8_I10_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O8_I10_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O8_I10_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O8_I10_R0_C01_rom_inst (.q(O8_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clock  (clk));
logic [10-1:0] O8_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O8_I13_R0_C01_rom_inst (.q(O8_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O8_I13_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O8_I13_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O8_I13_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O8_I13_R0_C01_rom_inst (.q(O8_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [10-1:0] O8_I14_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O8_I14_R0_C01_rom_inst (.q(O8_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clk(clk),.d(0),.we(0));
//assign O8_I14_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O8_I14_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O8_I14_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O8_I14_R0_C01_rom_inst (.q(O8_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clock  (clk));
logic [10-1:0] O8_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O8_I15_R0_C01_rom_inst (.q(O8_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O8_I15_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O8_I15_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O8_I15_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O8_I15_R0_C01_rom_inst (.q(O8_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [11-1:0] O8_I16_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O8_I16_R0_C02_rom_inst (.q(O8_I16_R0_C0_SM1 ),.address(input_fmap_16[7:0]),.clk(clk),.d(0),.we(0));
//assign O8_I16_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O8_I16_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O8_I16_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O8_I16_R0_C02_rom_inst (.q(O8_I16_R0_C0_SM1 ),.address(input_fmap_16[7:0]),.clock  (clk));
logic [10-1:0] O8_I17_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O8_I17_R0_C01_rom_inst (.q(O8_I17_R0_C0_SM1 ),.address(input_fmap_17[7:0]),.clk(clk),.d(0),.we(0));
//assign O8_I17_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O8_I17_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O8_I17_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O8_I17_R0_C01_rom_inst (.q(O8_I17_R0_C0_SM1 ),.address(input_fmap_17[7:0]),.clock  (clk));
logic [12-1:0] O8_I18_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_pw_O8_I18_R0_C04_rom_inst (.q(O8_I18_R0_C0_SM1 ),.address(input_fmap_18[7:0]),.clk(clk),.d(0),.we(0));
//assign O8_I18_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O8_I18_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O8_I18_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_pw_O8_I18_R0_C04_rom_inst (.q(O8_I18_R0_C0_SM1 ),.address(input_fmap_18[7:0]),.clock  (clk));
logic [10-1:0] O8_I20_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O8_I20_R0_C01_rom_inst (.q(O8_I20_R0_C0_SM1 ),.address(input_fmap_20[7:0]),.clk(clk),.d(0),.we(0));
//assign O8_I20_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O8_I20_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O8_I20_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O8_I20_R0_C01_rom_inst (.q(O8_I20_R0_C0_SM1 ),.address(input_fmap_20[7:0]),.clock  (clk));
logic [10-1:0] O8_I21_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O8_I21_R0_C01_rom_inst (.q(O8_I21_R0_C0_SM1 ),.address(input_fmap_21[7:0]),.clk(clk),.d(0),.we(0));
//assign O8_I21_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O8_I21_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O8_I21_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O8_I21_R0_C01_rom_inst (.q(O8_I21_R0_C0_SM1 ),.address(input_fmap_21[7:0]),.clock  (clk));
logic [10-1:0] O8_I24_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O8_I24_R0_C01_rom_inst (.q(O8_I24_R0_C0_SM1 ),.address(input_fmap_24[7:0]),.clk(clk),.d(0),.we(0));
//assign O8_I24_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O8_I24_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O8_I24_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O8_I24_R0_C01_rom_inst (.q(O8_I24_R0_C0_SM1 ),.address(input_fmap_24[7:0]),.clock  (clk));
logic [11-1:0] O8_I25_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O8_I25_R0_C03_rom_inst (.q(O8_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clk(clk),.d(0),.we(0));
//assign O8_I25_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O8_I25_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O8_I25_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O8_I25_R0_C03_rom_inst (.q(O8_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clock  (clk));
logic [11-1:0] O8_I26_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O8_I26_R0_C02_rom_inst (.q(O8_I26_R0_C0_SM1 ),.address(input_fmap_26[7:0]),.clk(clk),.d(0),.we(0));
//assign O8_I26_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O8_I26_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O8_I26_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O8_I26_R0_C02_rom_inst (.q(O8_I26_R0_C0_SM1 ),.address(input_fmap_26[7:0]),.clock  (clk));
logic [11-1:0] O8_I27_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O8_I27_R0_C03_rom_inst (.q(O8_I27_R0_C0_SM1 ),.address(input_fmap_27[7:0]),.clk(clk),.d(0),.we(0));
//assign O8_I27_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O8_I27_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O8_I27_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O8_I27_R0_C03_rom_inst (.q(O8_I27_R0_C0_SM1 ),.address(input_fmap_27[7:0]),.clock  (clk));
logic [10-1:0] O8_I29_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O8_I29_R0_C01_rom_inst (.q(O8_I29_R0_C0_SM1 ),.address(input_fmap_29[7:0]),.clk(clk),.d(0),.we(0));
//assign O8_I29_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O8_I29_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O8_I29_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O8_I29_R0_C01_rom_inst (.q(O8_I29_R0_C0_SM1 ),.address(input_fmap_29[7:0]),.clock  (clk));
logic [10-1:0] O8_I31_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O8_I31_R0_C01_rom_inst (.q(O8_I31_R0_C0_SM1 ),.address(input_fmap_31[7:0]),.clk(clk),.d(0),.we(0));
//assign O8_I31_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O8_I31_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O8_I31_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O8_I31_R0_C01_rom_inst (.q(O8_I31_R0_C0_SM1 ),.address(input_fmap_31[7:0]),.clock  (clk));
logic [12-1:0] O9_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_pw_O9_I0_R0_C04_rom_inst (.q(O9_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O9_I0_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O9_I0_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O9_I0_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_pw_O9_I0_R0_C04_rom_inst (.q(O9_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [10-1:0] O9_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O9_I1_R0_C01_rom_inst (.q(O9_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O9_I1_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O9_I1_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O9_I1_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O9_I1_R0_C01_rom_inst (.q(O9_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [10-1:0] O9_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O9_I2_R0_C01_rom_inst (.q(O9_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O9_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O9_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O9_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O9_I2_R0_C01_rom_inst (.q(O9_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [10-1:0] O9_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O9_I5_R0_C01_rom_inst (.q(O9_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O9_I5_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O9_I5_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O9_I5_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O9_I5_R0_C01_rom_inst (.q(O9_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [10-1:0] O9_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O9_I6_R0_C01_rom_inst (.q(O9_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O9_I6_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O9_I6_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O9_I6_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O9_I6_R0_C01_rom_inst (.q(O9_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [10-1:0] O9_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O9_I9_R0_C01_rom_inst (.q(O9_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O9_I9_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O9_I9_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O9_I9_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O9_I9_R0_C01_rom_inst (.q(O9_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [10-1:0] O9_I10_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O9_I10_R0_C01_rom_inst (.q(O9_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clk(clk),.d(0),.we(0));
//assign O9_I10_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O9_I10_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O9_I10_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O9_I10_R0_C01_rom_inst (.q(O9_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clock  (clk));
logic [10-1:0] O9_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O9_I11_R0_C01_rom_inst (.q(O9_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O9_I11_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O9_I11_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O9_I11_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O9_I11_R0_C01_rom_inst (.q(O9_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [11-1:0] O9_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O9_I13_R0_C03_rom_inst (.q(O9_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O9_I13_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O9_I13_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O9_I13_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O9_I13_R0_C03_rom_inst (.q(O9_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [10-1:0] O9_I14_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O9_I14_R0_C01_rom_inst (.q(O9_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clk(clk),.d(0),.we(0));
//assign O9_I14_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O9_I14_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O9_I14_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O9_I14_R0_C01_rom_inst (.q(O9_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clock  (clk));
logic [11-1:0] O9_I16_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O9_I16_R0_C02_rom_inst (.q(O9_I16_R0_C0_SM1 ),.address(input_fmap_16[7:0]),.clk(clk),.d(0),.we(0));
//assign O9_I16_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O9_I16_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O9_I16_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O9_I16_R0_C02_rom_inst (.q(O9_I16_R0_C0_SM1 ),.address(input_fmap_16[7:0]),.clock  (clk));
logic [10-1:0] O9_I17_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O9_I17_R0_C01_rom_inst (.q(O9_I17_R0_C0_SM1 ),.address(input_fmap_17[7:0]),.clk(clk),.d(0),.we(0));
//assign O9_I17_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O9_I17_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O9_I17_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O9_I17_R0_C01_rom_inst (.q(O9_I17_R0_C0_SM1 ),.address(input_fmap_17[7:0]),.clock  (clk));
logic [10-1:0] O9_I19_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O9_I19_R0_C01_rom_inst (.q(O9_I19_R0_C0_SM1 ),.address(input_fmap_19[7:0]),.clk(clk),.d(0),.we(0));
//assign O9_I19_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O9_I19_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O9_I19_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O9_I19_R0_C01_rom_inst (.q(O9_I19_R0_C0_SM1 ),.address(input_fmap_19[7:0]),.clock  (clk));
logic [10-1:0] O9_I24_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O9_I24_R0_C01_rom_inst (.q(O9_I24_R0_C0_SM1 ),.address(input_fmap_24[7:0]),.clk(clk),.d(0),.we(0));
//assign O9_I24_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O9_I24_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O9_I24_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O9_I24_R0_C01_rom_inst (.q(O9_I24_R0_C0_SM1 ),.address(input_fmap_24[7:0]),.clock  (clk));
logic [10-1:0] O9_I25_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O9_I25_R0_C01_rom_inst (.q(O9_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clk(clk),.d(0),.we(0));
//assign O9_I25_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O9_I25_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O9_I25_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O9_I25_R0_C01_rom_inst (.q(O9_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clock  (clk));
logic [10-1:0] O9_I26_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O9_I26_R0_C01_rom_inst (.q(O9_I26_R0_C0_SM1 ),.address(input_fmap_26[7:0]),.clk(clk),.d(0),.we(0));
//assign O9_I26_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O9_I26_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O9_I26_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O9_I26_R0_C01_rom_inst (.q(O9_I26_R0_C0_SM1 ),.address(input_fmap_26[7:0]),.clock  (clk));
logic [10-1:0] O9_I28_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O9_I28_R0_C01_rom_inst (.q(O9_I28_R0_C0_SM1 ),.address(input_fmap_28[7:0]),.clk(clk),.d(0),.we(0));
//assign O9_I28_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O9_I28_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O9_I28_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O9_I28_R0_C01_rom_inst (.q(O9_I28_R0_C0_SM1 ),.address(input_fmap_28[7:0]),.clock  (clk));
logic [10-1:0] O9_I31_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O9_I31_R0_C01_rom_inst (.q(O9_I31_R0_C0_SM1 ),.address(input_fmap_31[7:0]),.clk(clk),.d(0),.we(0));
//assign O9_I31_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O9_I31_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O9_I31_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O9_I31_R0_C01_rom_inst (.q(O9_I31_R0_C0_SM1 ),.address(input_fmap_31[7:0]),.clock  (clk));
logic [10-1:0] O10_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O10_I1_R0_C01_rom_inst (.q(O10_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O10_I1_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O10_I1_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O10_I1_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O10_I1_R0_C01_rom_inst (.q(O10_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [11-1:0] O10_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O10_I2_R0_C02_rom_inst (.q(O10_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O10_I2_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O10_I2_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O10_I2_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O10_I2_R0_C02_rom_inst (.q(O10_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [10-1:0] O10_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O10_I4_R0_C01_rom_inst (.q(O10_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O10_I4_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O10_I4_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O10_I4_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O10_I4_R0_C01_rom_inst (.q(O10_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [10-1:0] O10_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O10_I8_R0_C01_rom_inst (.q(O10_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O10_I8_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O10_I8_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O10_I8_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O10_I8_R0_C01_rom_inst (.q(O10_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [11-1:0] O10_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O10_I9_R0_C02_rom_inst (.q(O10_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O10_I9_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O10_I9_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O10_I9_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O10_I9_R0_C02_rom_inst (.q(O10_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [10-1:0] O10_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O10_I11_R0_C01_rom_inst (.q(O10_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O10_I11_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O10_I11_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O10_I11_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O10_I11_R0_C01_rom_inst (.q(O10_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [10-1:0] O10_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O10_I12_R0_C01_rom_inst (.q(O10_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O10_I12_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O10_I12_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O10_I12_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O10_I12_R0_C01_rom_inst (.q(O10_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [11-1:0] O10_I16_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O10_I16_R0_C03_rom_inst (.q(O10_I16_R0_C0_SM1 ),.address(input_fmap_16[7:0]),.clk(clk),.d(0),.we(0));
//assign O10_I16_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O10_I16_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O10_I16_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O10_I16_R0_C03_rom_inst (.q(O10_I16_R0_C0_SM1 ),.address(input_fmap_16[7:0]),.clock  (clk));
logic [11-1:0] O10_I19_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O10_I19_R0_C03_rom_inst (.q(O10_I19_R0_C0_SM1 ),.address(input_fmap_19[7:0]),.clk(clk),.d(0),.we(0));
//assign O10_I19_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O10_I19_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O10_I19_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O10_I19_R0_C03_rom_inst (.q(O10_I19_R0_C0_SM1 ),.address(input_fmap_19[7:0]),.clock  (clk));
logic [11-1:0] O10_I20_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O10_I20_R0_C02_rom_inst (.q(O10_I20_R0_C0_SM1 ),.address(input_fmap_20[7:0]),.clk(clk),.d(0),.we(0));
//assign O10_I20_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O10_I20_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O10_I20_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O10_I20_R0_C02_rom_inst (.q(O10_I20_R0_C0_SM1 ),.address(input_fmap_20[7:0]),.clock  (clk));
logic [10-1:0] O10_I23_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O10_I23_R0_C01_rom_inst (.q(O10_I23_R0_C0_SM1 ),.address(input_fmap_23[7:0]),.clk(clk),.d(0),.we(0));
//assign O10_I23_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O10_I23_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O10_I23_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O10_I23_R0_C01_rom_inst (.q(O10_I23_R0_C0_SM1 ),.address(input_fmap_23[7:0]),.clock  (clk));
logic [10-1:0] O10_I25_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O10_I25_R0_C01_rom_inst (.q(O10_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clk(clk),.d(0),.we(0));
//assign O10_I25_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O10_I25_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O10_I25_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O10_I25_R0_C01_rom_inst (.q(O10_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clock  (clk));
logic [11-1:0] O10_I26_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O10_I26_R0_C02_rom_inst (.q(O10_I26_R0_C0_SM1 ),.address(input_fmap_26[7:0]),.clk(clk),.d(0),.we(0));
//assign O10_I26_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O10_I26_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O10_I26_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O10_I26_R0_C02_rom_inst (.q(O10_I26_R0_C0_SM1 ),.address(input_fmap_26[7:0]),.clock  (clk));
logic [10-1:0] O10_I28_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O10_I28_R0_C01_rom_inst (.q(O10_I28_R0_C0_SM1 ),.address(input_fmap_28[7:0]),.clk(clk),.d(0),.we(0));
//assign O10_I28_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O10_I28_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O10_I28_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O10_I28_R0_C01_rom_inst (.q(O10_I28_R0_C0_SM1 ),.address(input_fmap_28[7:0]),.clock  (clk));
logic [10-1:0] O10_I30_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O10_I30_R0_C01_rom_inst (.q(O10_I30_R0_C0_SM1 ),.address(input_fmap_30[7:0]),.clk(clk),.d(0),.we(0));
//assign O10_I30_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O10_I30_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O10_I30_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O10_I30_R0_C01_rom_inst (.q(O10_I30_R0_C0_SM1 ),.address(input_fmap_30[7:0]),.clock  (clk));
logic [10-1:0] O10_I31_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O10_I31_R0_C01_rom_inst (.q(O10_I31_R0_C0_SM1 ),.address(input_fmap_31[7:0]),.clk(clk),.d(0),.we(0));
//assign O10_I31_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O10_I31_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O10_I31_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O10_I31_R0_C01_rom_inst (.q(O10_I31_R0_C0_SM1 ),.address(input_fmap_31[7:0]),.clock  (clk));
logic [11-1:0] O11_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O11_I0_R0_C02_rom_inst (.q(O11_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I0_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O11_I0_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O11_I0_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O11_I0_R0_C02_rom_inst (.q(O11_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [10-1:0] O11_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O11_I1_R0_C01_rom_inst (.q(O11_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I1_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O11_I1_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O11_I1_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O11_I1_R0_C01_rom_inst (.q(O11_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [10-1:0] O11_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O11_I5_R0_C01_rom_inst (.q(O11_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I5_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O11_I5_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O11_I5_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O11_I5_R0_C01_rom_inst (.q(O11_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [10-1:0] O11_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O11_I7_R0_C01_rom_inst (.q(O11_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I7_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O11_I7_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O11_I7_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O11_I7_R0_C01_rom_inst (.q(O11_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [11-1:0] O11_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O11_I8_R0_C02_rom_inst (.q(O11_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I8_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O11_I8_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O11_I8_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O11_I8_R0_C02_rom_inst (.q(O11_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [10-1:0] O11_I10_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O11_I10_R0_C01_rom_inst (.q(O11_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I10_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O11_I10_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O11_I10_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O11_I10_R0_C01_rom_inst (.q(O11_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clock  (clk));
logic [10-1:0] O11_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O11_I11_R0_C01_rom_inst (.q(O11_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I11_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O11_I11_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O11_I11_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O11_I11_R0_C01_rom_inst (.q(O11_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [11-1:0] O11_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O11_I12_R0_C02_rom_inst (.q(O11_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I12_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O11_I12_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O11_I12_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O11_I12_R0_C02_rom_inst (.q(O11_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [11-1:0] O11_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O11_I13_R0_C02_rom_inst (.q(O11_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I13_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O11_I13_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O11_I13_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O11_I13_R0_C02_rom_inst (.q(O11_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [10-1:0] O11_I16_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O11_I16_R0_C01_rom_inst (.q(O11_I16_R0_C0_SM1 ),.address(input_fmap_16[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I16_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O11_I16_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O11_I16_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O11_I16_R0_C01_rom_inst (.q(O11_I16_R0_C0_SM1 ),.address(input_fmap_16[7:0]),.clock  (clk));
logic [10-1:0] O11_I19_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O11_I19_R0_C01_rom_inst (.q(O11_I19_R0_C0_SM1 ),.address(input_fmap_19[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I19_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O11_I19_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O11_I19_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O11_I19_R0_C01_rom_inst (.q(O11_I19_R0_C0_SM1 ),.address(input_fmap_19[7:0]),.clock  (clk));
logic [10-1:0] O11_I20_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O11_I20_R0_C01_rom_inst (.q(O11_I20_R0_C0_SM1 ),.address(input_fmap_20[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I20_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O11_I20_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O11_I20_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O11_I20_R0_C01_rom_inst (.q(O11_I20_R0_C0_SM1 ),.address(input_fmap_20[7:0]),.clock  (clk));
logic [10-1:0] O11_I22_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O11_I22_R0_C01_rom_inst (.q(O11_I22_R0_C0_SM1 ),.address(input_fmap_22[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I22_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O11_I22_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O11_I22_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O11_I22_R0_C01_rom_inst (.q(O11_I22_R0_C0_SM1 ),.address(input_fmap_22[7:0]),.clock  (clk));
logic [10-1:0] O11_I24_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O11_I24_R0_C01_rom_inst (.q(O11_I24_R0_C0_SM1 ),.address(input_fmap_24[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I24_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O11_I24_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O11_I24_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O11_I24_R0_C01_rom_inst (.q(O11_I24_R0_C0_SM1 ),.address(input_fmap_24[7:0]),.clock  (clk));
logic [11-1:0] O11_I25_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O11_I25_R0_C02_rom_inst (.q(O11_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I25_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O11_I25_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O11_I25_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O11_I25_R0_C02_rom_inst (.q(O11_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clock  (clk));
logic [10-1:0] O11_I26_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O11_I26_R0_C01_rom_inst (.q(O11_I26_R0_C0_SM1 ),.address(input_fmap_26[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I26_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O11_I26_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O11_I26_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O11_I26_R0_C01_rom_inst (.q(O11_I26_R0_C0_SM1 ),.address(input_fmap_26[7:0]),.clock  (clk));
logic [10-1:0] O11_I27_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O11_I27_R0_C01_rom_inst (.q(O11_I27_R0_C0_SM1 ),.address(input_fmap_27[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I27_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O11_I27_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O11_I27_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O11_I27_R0_C01_rom_inst (.q(O11_I27_R0_C0_SM1 ),.address(input_fmap_27[7:0]),.clock  (clk));
logic [11-1:0] O11_I30_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O11_I30_R0_C03_rom_inst (.q(O11_I30_R0_C0_SM1 ),.address(input_fmap_30[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I30_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O11_I30_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O11_I30_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O11_I30_R0_C03_rom_inst (.q(O11_I30_R0_C0_SM1 ),.address(input_fmap_30[7:0]),.clock  (clk));
logic [10-1:0] O11_I31_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O11_I31_R0_C01_rom_inst (.q(O11_I31_R0_C0_SM1 ),.address(input_fmap_31[7:0]),.clk(clk),.d(0),.we(0));
//assign O11_I31_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O11_I31_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O11_I31_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O11_I31_R0_C01_rom_inst (.q(O11_I31_R0_C0_SM1 ),.address(input_fmap_31[7:0]),.clock  (clk));
logic [11-1:0] O12_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O12_I0_R0_C02_rom_inst (.q(O12_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I0_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O12_I0_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O12_I0_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O12_I0_R0_C02_rom_inst (.q(O12_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [12-1:0] O12_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_pw_O12_I1_R0_C05_rom_inst (.q(O12_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I1_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O12_I1_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O12_I1_R0_C05_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_pw_O12_I1_R0_C05_rom_inst (.q(O12_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [10-1:0] O12_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O12_I2_R0_C01_rom_inst (.q(O12_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O12_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O12_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O12_I2_R0_C01_rom_inst (.q(O12_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [11-1:0] O12_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O12_I3_R0_C02_rom_inst (.q(O12_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I3_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O12_I3_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O12_I3_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O12_I3_R0_C02_rom_inst (.q(O12_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [11-1:0] O12_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O12_I5_R0_C03_rom_inst (.q(O12_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I5_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O12_I5_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O12_I5_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O12_I5_R0_C03_rom_inst (.q(O12_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [10-1:0] O12_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O12_I6_R0_C01_rom_inst (.q(O12_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I6_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O12_I6_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O12_I6_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O12_I6_R0_C01_rom_inst (.q(O12_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [10-1:0] O12_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O12_I7_R0_C01_rom_inst (.q(O12_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I7_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O12_I7_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O12_I7_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O12_I7_R0_C01_rom_inst (.q(O12_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [11-1:0] O12_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O12_I9_R0_C02_rom_inst (.q(O12_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I9_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O12_I9_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O12_I9_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O12_I9_R0_C02_rom_inst (.q(O12_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [10-1:0] O12_I10_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O12_I10_R0_C01_rom_inst (.q(O12_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I10_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O12_I10_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O12_I10_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O12_I10_R0_C01_rom_inst (.q(O12_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clock  (clk));
logic [10-1:0] O12_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O12_I11_R0_C01_rom_inst (.q(O12_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I11_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O12_I11_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O12_I11_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O12_I11_R0_C01_rom_inst (.q(O12_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [10-1:0] O12_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O12_I12_R0_C01_rom_inst (.q(O12_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I12_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O12_I12_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O12_I12_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O12_I12_R0_C01_rom_inst (.q(O12_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [11-1:0] O12_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O12_I13_R0_C03_rom_inst (.q(O12_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I13_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O12_I13_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O12_I13_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O12_I13_R0_C03_rom_inst (.q(O12_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [10-1:0] O12_I14_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O12_I14_R0_C01_rom_inst (.q(O12_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I14_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O12_I14_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O12_I14_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O12_I14_R0_C01_rom_inst (.q(O12_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clock  (clk));
logic [10-1:0] O12_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O12_I15_R0_C01_rom_inst (.q(O12_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I15_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O12_I15_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O12_I15_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O12_I15_R0_C01_rom_inst (.q(O12_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [12-1:0] O12_I17_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_pw_O12_I17_R0_C04_rom_inst (.q(O12_I17_R0_C0_SM1 ),.address(input_fmap_17[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I17_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O12_I17_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O12_I17_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_pw_O12_I17_R0_C04_rom_inst (.q(O12_I17_R0_C0_SM1 ),.address(input_fmap_17[7:0]),.clock  (clk));
logic [10-1:0] O12_I18_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O12_I18_R0_C01_rom_inst (.q(O12_I18_R0_C0_SM1 ),.address(input_fmap_18[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I18_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O12_I18_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O12_I18_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O12_I18_R0_C01_rom_inst (.q(O12_I18_R0_C0_SM1 ),.address(input_fmap_18[7:0]),.clock  (clk));
logic [11-1:0] O12_I20_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O12_I20_R0_C02_rom_inst (.q(O12_I20_R0_C0_SM1 ),.address(input_fmap_20[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I20_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O12_I20_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O12_I20_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O12_I20_R0_C02_rom_inst (.q(O12_I20_R0_C0_SM1 ),.address(input_fmap_20[7:0]),.clock  (clk));
logic [10-1:0] O12_I24_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O12_I24_R0_C01_rom_inst (.q(O12_I24_R0_C0_SM1 ),.address(input_fmap_24[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I24_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O12_I24_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O12_I24_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O12_I24_R0_C01_rom_inst (.q(O12_I24_R0_C0_SM1 ),.address(input_fmap_24[7:0]),.clock  (clk));
logic [11-1:0] O12_I25_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O12_I25_R0_C02_rom_inst (.q(O12_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I25_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O12_I25_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O12_I25_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O12_I25_R0_C02_rom_inst (.q(O12_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clock  (clk));
logic [11-1:0] O12_I27_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O12_I27_R0_C03_rom_inst (.q(O12_I27_R0_C0_SM1 ),.address(input_fmap_27[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I27_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O12_I27_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O12_I27_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O12_I27_R0_C03_rom_inst (.q(O12_I27_R0_C0_SM1 ),.address(input_fmap_27[7:0]),.clock  (clk));
logic [10-1:0] O12_I29_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O12_I29_R0_C01_rom_inst (.q(O12_I29_R0_C0_SM1 ),.address(input_fmap_29[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I29_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O12_I29_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O12_I29_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O12_I29_R0_C01_rom_inst (.q(O12_I29_R0_C0_SM1 ),.address(input_fmap_29[7:0]),.clock  (clk));
logic [10-1:0] O12_I30_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O12_I30_R0_C01_rom_inst (.q(O12_I30_R0_C0_SM1 ),.address(input_fmap_30[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I30_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O12_I30_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O12_I30_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O12_I30_R0_C01_rom_inst (.q(O12_I30_R0_C0_SM1 ),.address(input_fmap_30[7:0]),.clock  (clk));
logic [10-1:0] O12_I31_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O12_I31_R0_C01_rom_inst (.q(O12_I31_R0_C0_SM1 ),.address(input_fmap_31[7:0]),.clk(clk),.d(0),.we(0));
//assign O12_I31_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O12_I31_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O12_I31_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O12_I31_R0_C01_rom_inst (.q(O12_I31_R0_C0_SM1 ),.address(input_fmap_31[7:0]),.clock  (clk));
logic [11-1:0] O13_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O13_I1_R0_C02_rom_inst (.q(O13_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O13_I1_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O13_I1_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O13_I1_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O13_I1_R0_C02_rom_inst (.q(O13_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [10-1:0] O13_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O13_I2_R0_C01_rom_inst (.q(O13_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O13_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O13_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O13_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O13_I2_R0_C01_rom_inst (.q(O13_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [10-1:0] O13_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O13_I4_R0_C01_rom_inst (.q(O13_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O13_I4_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O13_I4_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O13_I4_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O13_I4_R0_C01_rom_inst (.q(O13_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [10-1:0] O13_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O13_I5_R0_C01_rom_inst (.q(O13_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O13_I5_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O13_I5_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O13_I5_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O13_I5_R0_C01_rom_inst (.q(O13_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [10-1:0] O13_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O13_I9_R0_C01_rom_inst (.q(O13_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O13_I9_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O13_I9_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O13_I9_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O13_I9_R0_C01_rom_inst (.q(O13_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [10-1:0] O13_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O13_I11_R0_C01_rom_inst (.q(O13_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O13_I11_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O13_I11_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O13_I11_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O13_I11_R0_C01_rom_inst (.q(O13_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [10-1:0] O13_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O13_I15_R0_C01_rom_inst (.q(O13_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O13_I15_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O13_I15_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O13_I15_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O13_I15_R0_C01_rom_inst (.q(O13_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [10-1:0] O13_I16_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O13_I16_R0_C01_rom_inst (.q(O13_I16_R0_C0_SM1 ),.address(input_fmap_16[7:0]),.clk(clk),.d(0),.we(0));
//assign O13_I16_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O13_I16_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O13_I16_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O13_I16_R0_C01_rom_inst (.q(O13_I16_R0_C0_SM1 ),.address(input_fmap_16[7:0]),.clock  (clk));
logic [10-1:0] O13_I20_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O13_I20_R0_C01_rom_inst (.q(O13_I20_R0_C0_SM1 ),.address(input_fmap_20[7:0]),.clk(clk),.d(0),.we(0));
//assign O13_I20_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O13_I20_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O13_I20_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O13_I20_R0_C01_rom_inst (.q(O13_I20_R0_C0_SM1 ),.address(input_fmap_20[7:0]),.clock  (clk));
logic [10-1:0] O13_I21_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O13_I21_R0_C01_rom_inst (.q(O13_I21_R0_C0_SM1 ),.address(input_fmap_21[7:0]),.clk(clk),.d(0),.we(0));
//assign O13_I21_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O13_I21_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O13_I21_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O13_I21_R0_C01_rom_inst (.q(O13_I21_R0_C0_SM1 ),.address(input_fmap_21[7:0]),.clock  (clk));
logic [12-1:0] O13_I22_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_pw_O13_I22_R0_C05_rom_inst (.q(O13_I22_R0_C0_SM1 ),.address(input_fmap_22[7:0]),.clk(clk),.d(0),.we(0));
//assign O13_I22_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O13_I22_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O13_I22_R0_C05_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_pw_O13_I22_R0_C05_rom_inst (.q(O13_I22_R0_C0_SM1 ),.address(input_fmap_22[7:0]),.clock  (clk));
logic [11-1:0] O13_I25_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O13_I25_R0_C02_rom_inst (.q(O13_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clk(clk),.d(0),.we(0));
//assign O13_I25_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O13_I25_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O13_I25_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O13_I25_R0_C02_rom_inst (.q(O13_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clock  (clk));
logic [10-1:0] O13_I27_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O13_I27_R0_C01_rom_inst (.q(O13_I27_R0_C0_SM1 ),.address(input_fmap_27[7:0]),.clk(clk),.d(0),.we(0));
//assign O13_I27_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O13_I27_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O13_I27_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O13_I27_R0_C01_rom_inst (.q(O13_I27_R0_C0_SM1 ),.address(input_fmap_27[7:0]),.clock  (clk));
logic [10-1:0] O13_I28_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O13_I28_R0_C01_rom_inst (.q(O13_I28_R0_C0_SM1 ),.address(input_fmap_28[7:0]),.clk(clk),.d(0),.we(0));
//assign O13_I28_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O13_I28_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O13_I28_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O13_I28_R0_C01_rom_inst (.q(O13_I28_R0_C0_SM1 ),.address(input_fmap_28[7:0]),.clock  (clk));
logic [10-1:0] O13_I30_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O13_I30_R0_C01_rom_inst (.q(O13_I30_R0_C0_SM1 ),.address(input_fmap_30[7:0]),.clk(clk),.d(0),.we(0));
//assign O13_I30_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O13_I30_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O13_I30_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O13_I30_R0_C01_rom_inst (.q(O13_I30_R0_C0_SM1 ),.address(input_fmap_30[7:0]),.clock  (clk));
logic [11-1:0] O14_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O14_I2_R0_C02_rom_inst (.q(O14_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I2_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O14_I2_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O14_I2_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O14_I2_R0_C02_rom_inst (.q(O14_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [10-1:0] O14_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O14_I3_R0_C01_rom_inst (.q(O14_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I3_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O14_I3_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O14_I3_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O14_I3_R0_C01_rom_inst (.q(O14_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [10-1:0] O14_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O14_I5_R0_C01_rom_inst (.q(O14_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I5_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O14_I5_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O14_I5_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O14_I5_R0_C01_rom_inst (.q(O14_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [10-1:0] O14_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O14_I6_R0_C01_rom_inst (.q(O14_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I6_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O14_I6_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O14_I6_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O14_I6_R0_C01_rom_inst (.q(O14_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [11-1:0] O14_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O14_I9_R0_C02_rom_inst (.q(O14_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I9_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O14_I9_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O14_I9_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O14_I9_R0_C02_rom_inst (.q(O14_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [10-1:0] O14_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O14_I11_R0_C01_rom_inst (.q(O14_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I11_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O14_I11_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O14_I11_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O14_I11_R0_C01_rom_inst (.q(O14_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [10-1:0] O14_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O14_I13_R0_C01_rom_inst (.q(O14_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I13_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O14_I13_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O14_I13_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O14_I13_R0_C01_rom_inst (.q(O14_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [11-1:0] O14_I16_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O14_I16_R0_C02_rom_inst (.q(O14_I16_R0_C0_SM1 ),.address(input_fmap_16[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I16_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O14_I16_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O14_I16_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O14_I16_R0_C02_rom_inst (.q(O14_I16_R0_C0_SM1 ),.address(input_fmap_16[7:0]),.clock  (clk));
logic [10-1:0] O14_I17_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O14_I17_R0_C01_rom_inst (.q(O14_I17_R0_C0_SM1 ),.address(input_fmap_17[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I17_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O14_I17_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O14_I17_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O14_I17_R0_C01_rom_inst (.q(O14_I17_R0_C0_SM1 ),.address(input_fmap_17[7:0]),.clock  (clk));
logic [10-1:0] O14_I18_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O14_I18_R0_C01_rom_inst (.q(O14_I18_R0_C0_SM1 ),.address(input_fmap_18[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I18_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O14_I18_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O14_I18_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O14_I18_R0_C01_rom_inst (.q(O14_I18_R0_C0_SM1 ),.address(input_fmap_18[7:0]),.clock  (clk));
logic [11-1:0] O14_I19_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O14_I19_R0_C03_rom_inst (.q(O14_I19_R0_C0_SM1 ),.address(input_fmap_19[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I19_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O14_I19_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O14_I19_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O14_I19_R0_C03_rom_inst (.q(O14_I19_R0_C0_SM1 ),.address(input_fmap_19[7:0]),.clock  (clk));
logic [11-1:0] O14_I20_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O14_I20_R0_C03_rom_inst (.q(O14_I20_R0_C0_SM1 ),.address(input_fmap_20[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I20_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O14_I20_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O14_I20_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O14_I20_R0_C03_rom_inst (.q(O14_I20_R0_C0_SM1 ),.address(input_fmap_20[7:0]),.clock  (clk));
logic [10-1:0] O14_I24_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O14_I24_R0_C01_rom_inst (.q(O14_I24_R0_C0_SM1 ),.address(input_fmap_24[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I24_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O14_I24_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O14_I24_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O14_I24_R0_C01_rom_inst (.q(O14_I24_R0_C0_SM1 ),.address(input_fmap_24[7:0]),.clock  (clk));
logic [11-1:0] O14_I25_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O14_I25_R0_C03_rom_inst (.q(O14_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I25_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O14_I25_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O14_I25_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O14_I25_R0_C03_rom_inst (.q(O14_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clock  (clk));
logic [10-1:0] O14_I26_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O14_I26_R0_C01_rom_inst (.q(O14_I26_R0_C0_SM1 ),.address(input_fmap_26[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I26_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O14_I26_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O14_I26_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O14_I26_R0_C01_rom_inst (.q(O14_I26_R0_C0_SM1 ),.address(input_fmap_26[7:0]),.clock  (clk));
logic [10-1:0] O14_I27_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O14_I27_R0_C01_rom_inst (.q(O14_I27_R0_C0_SM1 ),.address(input_fmap_27[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I27_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O14_I27_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O14_I27_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O14_I27_R0_C01_rom_inst (.q(O14_I27_R0_C0_SM1 ),.address(input_fmap_27[7:0]),.clock  (clk));
logic [10-1:0] O14_I28_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O14_I28_R0_C01_rom_inst (.q(O14_I28_R0_C0_SM1 ),.address(input_fmap_28[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I28_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O14_I28_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O14_I28_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O14_I28_R0_C01_rom_inst (.q(O14_I28_R0_C0_SM1 ),.address(input_fmap_28[7:0]),.clock  (clk));
logic [10-1:0] O14_I29_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O14_I29_R0_C01_rom_inst (.q(O14_I29_R0_C0_SM1 ),.address(input_fmap_29[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I29_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O14_I29_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O14_I29_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O14_I29_R0_C01_rom_inst (.q(O14_I29_R0_C0_SM1 ),.address(input_fmap_29[7:0]),.clock  (clk));
logic [10-1:0] O14_I30_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O14_I30_R0_C01_rom_inst (.q(O14_I30_R0_C0_SM1 ),.address(input_fmap_30[7:0]),.clk(clk),.d(0),.we(0));
//assign O14_I30_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O14_I30_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O14_I30_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O14_I30_R0_C01_rom_inst (.q(O14_I30_R0_C0_SM1 ),.address(input_fmap_30[7:0]),.clock  (clk));
logic [11-1:0] O15_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O15_I0_R0_C02_rom_inst (.q(O15_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I0_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O15_I0_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O15_I0_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O15_I0_R0_C02_rom_inst (.q(O15_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [10-1:0] O15_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O15_I2_R0_C01_rom_inst (.q(O15_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O15_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O15_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O15_I2_R0_C01_rom_inst (.q(O15_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [11-1:0] O15_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O15_I4_R0_C03_rom_inst (.q(O15_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I4_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O15_I4_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O15_I4_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O15_I4_R0_C03_rom_inst (.q(O15_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [10-1:0] O15_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O15_I5_R0_C01_rom_inst (.q(O15_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I5_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O15_I5_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O15_I5_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O15_I5_R0_C01_rom_inst (.q(O15_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [10-1:0] O15_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O15_I6_R0_C01_rom_inst (.q(O15_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I6_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O15_I6_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O15_I6_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O15_I6_R0_C01_rom_inst (.q(O15_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [11-1:0] O15_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O15_I7_R0_C02_rom_inst (.q(O15_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I7_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O15_I7_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O15_I7_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O15_I7_R0_C02_rom_inst (.q(O15_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [11-1:0] O15_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O15_I8_R0_C02_rom_inst (.q(O15_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I8_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O15_I8_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O15_I8_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O15_I8_R0_C02_rom_inst (.q(O15_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [10-1:0] O15_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O15_I9_R0_C01_rom_inst (.q(O15_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I9_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O15_I9_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O15_I9_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O15_I9_R0_C01_rom_inst (.q(O15_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [10-1:0] O15_I10_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O15_I10_R0_C01_rom_inst (.q(O15_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I10_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O15_I10_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O15_I10_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O15_I10_R0_C01_rom_inst (.q(O15_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clock  (clk));
logic [11-1:0] O15_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O15_I11_R0_C02_rom_inst (.q(O15_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I11_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O15_I11_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O15_I11_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O15_I11_R0_C02_rom_inst (.q(O15_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [10-1:0] O15_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O15_I12_R0_C01_rom_inst (.q(O15_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I12_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O15_I12_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O15_I12_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O15_I12_R0_C01_rom_inst (.q(O15_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [10-1:0] O15_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O15_I13_R0_C01_rom_inst (.q(O15_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I13_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O15_I13_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O15_I13_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O15_I13_R0_C01_rom_inst (.q(O15_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [10-1:0] O15_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O15_I15_R0_C01_rom_inst (.q(O15_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I15_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O15_I15_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O15_I15_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O15_I15_R0_C01_rom_inst (.q(O15_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [12-1:0] O15_I16_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_pw_O15_I16_R0_C04_rom_inst (.q(O15_I16_R0_C0_SM1 ),.address(input_fmap_16[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I16_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O15_I16_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O15_I16_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_pw_O15_I16_R0_C04_rom_inst (.q(O15_I16_R0_C0_SM1 ),.address(input_fmap_16[7:0]),.clock  (clk));
logic [10-1:0] O15_I18_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O15_I18_R0_C01_rom_inst (.q(O15_I18_R0_C0_SM1 ),.address(input_fmap_18[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I18_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O15_I18_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O15_I18_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O15_I18_R0_C01_rom_inst (.q(O15_I18_R0_C0_SM1 ),.address(input_fmap_18[7:0]),.clock  (clk));
logic [10-1:0] O15_I19_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O15_I19_R0_C01_rom_inst (.q(O15_I19_R0_C0_SM1 ),.address(input_fmap_19[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I19_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O15_I19_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O15_I19_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O15_I19_R0_C01_rom_inst (.q(O15_I19_R0_C0_SM1 ),.address(input_fmap_19[7:0]),.clock  (clk));
logic [10-1:0] O15_I20_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O15_I20_R0_C01_rom_inst (.q(O15_I20_R0_C0_SM1 ),.address(input_fmap_20[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I20_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O15_I20_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O15_I20_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O15_I20_R0_C01_rom_inst (.q(O15_I20_R0_C0_SM1 ),.address(input_fmap_20[7:0]),.clock  (clk));
logic [10-1:0] O15_I21_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O15_I21_R0_C01_rom_inst (.q(O15_I21_R0_C0_SM1 ),.address(input_fmap_21[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I21_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O15_I21_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O15_I21_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O15_I21_R0_C01_rom_inst (.q(O15_I21_R0_C0_SM1 ),.address(input_fmap_21[7:0]),.clock  (clk));
logic [10-1:0] O15_I22_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O15_I22_R0_C01_rom_inst (.q(O15_I22_R0_C0_SM1 ),.address(input_fmap_22[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I22_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O15_I22_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O15_I22_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O15_I22_R0_C01_rom_inst (.q(O15_I22_R0_C0_SM1 ),.address(input_fmap_22[7:0]),.clock  (clk));
logic [10-1:0] O15_I23_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O15_I23_R0_C01_rom_inst (.q(O15_I23_R0_C0_SM1 ),.address(input_fmap_23[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I23_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O15_I23_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O15_I23_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O15_I23_R0_C01_rom_inst (.q(O15_I23_R0_C0_SM1 ),.address(input_fmap_23[7:0]),.clock  (clk));
logic [11-1:0] O15_I24_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O15_I24_R0_C03_rom_inst (.q(O15_I24_R0_C0_SM1 ),.address(input_fmap_24[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I24_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O15_I24_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O15_I24_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O15_I24_R0_C03_rom_inst (.q(O15_I24_R0_C0_SM1 ),.address(input_fmap_24[7:0]),.clock  (clk));
logic [10-1:0] O15_I25_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O15_I25_R0_C01_rom_inst (.q(O15_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I25_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O15_I25_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O15_I25_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O15_I25_R0_C01_rom_inst (.q(O15_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clock  (clk));
logic [11-1:0] O15_I26_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O15_I26_R0_C02_rom_inst (.q(O15_I26_R0_C0_SM1 ),.address(input_fmap_26[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I26_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O15_I26_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O15_I26_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O15_I26_R0_C02_rom_inst (.q(O15_I26_R0_C0_SM1 ),.address(input_fmap_26[7:0]),.clock  (clk));
logic [10-1:0] O15_I28_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O15_I28_R0_C01_rom_inst (.q(O15_I28_R0_C0_SM1 ),.address(input_fmap_28[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I28_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O15_I28_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O15_I28_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O15_I28_R0_C01_rom_inst (.q(O15_I28_R0_C0_SM1 ),.address(input_fmap_28[7:0]),.clock  (clk));
logic [11-1:0] O15_I30_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O15_I30_R0_C02_rom_inst (.q(O15_I30_R0_C0_SM1 ),.address(input_fmap_30[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I30_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O15_I30_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O15_I30_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O15_I30_R0_C02_rom_inst (.q(O15_I30_R0_C0_SM1 ),.address(input_fmap_30[7:0]),.clock  (clk));
logic [11-1:0] O15_I31_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O15_I31_R0_C02_rom_inst (.q(O15_I31_R0_C0_SM1 ),.address(input_fmap_31[7:0]),.clk(clk),.d(0),.we(0));
//assign O15_I31_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O15_I31_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O15_I31_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O15_I31_R0_C02_rom_inst (.q(O15_I31_R0_C0_SM1 ),.address(input_fmap_31[7:0]),.clock  (clk));
logic [10-1:0] O16_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O16_I1_R0_C01_rom_inst (.q(O16_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O16_I1_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O16_I1_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O16_I1_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O16_I1_R0_C01_rom_inst (.q(O16_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [10-1:0] O16_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O16_I4_R0_C01_rom_inst (.q(O16_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O16_I4_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O16_I4_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O16_I4_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O16_I4_R0_C01_rom_inst (.q(O16_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [10-1:0] O16_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O16_I5_R0_C01_rom_inst (.q(O16_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O16_I5_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O16_I5_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O16_I5_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O16_I5_R0_C01_rom_inst (.q(O16_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [10-1:0] O16_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O16_I7_R0_C01_rom_inst (.q(O16_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O16_I7_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O16_I7_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O16_I7_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O16_I7_R0_C01_rom_inst (.q(O16_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [10-1:0] O16_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O16_I8_R0_C01_rom_inst (.q(O16_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O16_I8_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O16_I8_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O16_I8_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O16_I8_R0_C01_rom_inst (.q(O16_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [11-1:0] O16_I10_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O16_I10_R0_C03_rom_inst (.q(O16_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clk(clk),.d(0),.we(0));
//assign O16_I10_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O16_I10_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O16_I10_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O16_I10_R0_C03_rom_inst (.q(O16_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clock  (clk));
logic [10-1:0] O16_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O16_I11_R0_C01_rom_inst (.q(O16_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O16_I11_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O16_I11_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O16_I11_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O16_I11_R0_C01_rom_inst (.q(O16_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [10-1:0] O16_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O16_I12_R0_C01_rom_inst (.q(O16_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O16_I12_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O16_I12_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O16_I12_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O16_I12_R0_C01_rom_inst (.q(O16_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [10-1:0] O16_I14_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O16_I14_R0_C01_rom_inst (.q(O16_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clk(clk),.d(0),.we(0));
//assign O16_I14_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O16_I14_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O16_I14_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O16_I14_R0_C01_rom_inst (.q(O16_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clock  (clk));
logic [10-1:0] O16_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O16_I15_R0_C01_rom_inst (.q(O16_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O16_I15_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O16_I15_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O16_I15_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O16_I15_R0_C01_rom_inst (.q(O16_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [11-1:0] O16_I17_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O16_I17_R0_C02_rom_inst (.q(O16_I17_R0_C0_SM1 ),.address(input_fmap_17[7:0]),.clk(clk),.d(0),.we(0));
//assign O16_I17_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O16_I17_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O16_I17_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O16_I17_R0_C02_rom_inst (.q(O16_I17_R0_C0_SM1 ),.address(input_fmap_17[7:0]),.clock  (clk));
logic [12-1:0] O16_I18_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_pw_O16_I18_R0_C06_rom_inst (.q(O16_I18_R0_C0_SM1 ),.address(input_fmap_18[7:0]),.clk(clk),.d(0),.we(0));
//assign O16_I18_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O16_I18_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O16_I18_R0_C06_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_pw_O16_I18_R0_C06_rom_inst (.q(O16_I18_R0_C0_SM1 ),.address(input_fmap_18[7:0]),.clock  (clk));
logic [10-1:0] O16_I19_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O16_I19_R0_C01_rom_inst (.q(O16_I19_R0_C0_SM1 ),.address(input_fmap_19[7:0]),.clk(clk),.d(0),.we(0));
//assign O16_I19_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O16_I19_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O16_I19_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O16_I19_R0_C01_rom_inst (.q(O16_I19_R0_C0_SM1 ),.address(input_fmap_19[7:0]),.clock  (clk));
logic [10-1:0] O16_I20_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O16_I20_R0_C01_rom_inst (.q(O16_I20_R0_C0_SM1 ),.address(input_fmap_20[7:0]),.clk(clk),.d(0),.we(0));
//assign O16_I20_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O16_I20_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O16_I20_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O16_I20_R0_C01_rom_inst (.q(O16_I20_R0_C0_SM1 ),.address(input_fmap_20[7:0]),.clock  (clk));
logic [10-1:0] O16_I23_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O16_I23_R0_C01_rom_inst (.q(O16_I23_R0_C0_SM1 ),.address(input_fmap_23[7:0]),.clk(clk),.d(0),.we(0));
//assign O16_I23_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O16_I23_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O16_I23_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O16_I23_R0_C01_rom_inst (.q(O16_I23_R0_C0_SM1 ),.address(input_fmap_23[7:0]),.clock  (clk));
logic [10-1:0] O16_I25_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O16_I25_R0_C01_rom_inst (.q(O16_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clk(clk),.d(0),.we(0));
//assign O16_I25_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O16_I25_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O16_I25_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O16_I25_R0_C01_rom_inst (.q(O16_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clock  (clk));
logic [10-1:0] O16_I26_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O16_I26_R0_C01_rom_inst (.q(O16_I26_R0_C0_SM1 ),.address(input_fmap_26[7:0]),.clk(clk),.d(0),.we(0));
//assign O16_I26_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O16_I26_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O16_I26_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O16_I26_R0_C01_rom_inst (.q(O16_I26_R0_C0_SM1 ),.address(input_fmap_26[7:0]),.clock  (clk));
logic [11-1:0] O16_I27_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O16_I27_R0_C02_rom_inst (.q(O16_I27_R0_C0_SM1 ),.address(input_fmap_27[7:0]),.clk(clk),.d(0),.we(0));
//assign O16_I27_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O16_I27_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O16_I27_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O16_I27_R0_C02_rom_inst (.q(O16_I27_R0_C0_SM1 ),.address(input_fmap_27[7:0]),.clock  (clk));
logic [10-1:0] O16_I28_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O16_I28_R0_C01_rom_inst (.q(O16_I28_R0_C0_SM1 ),.address(input_fmap_28[7:0]),.clk(clk),.d(0),.we(0));
//assign O16_I28_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O16_I28_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O16_I28_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O16_I28_R0_C01_rom_inst (.q(O16_I28_R0_C0_SM1 ),.address(input_fmap_28[7:0]),.clock  (clk));
logic [10-1:0] O16_I29_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O16_I29_R0_C01_rom_inst (.q(O16_I29_R0_C0_SM1 ),.address(input_fmap_29[7:0]),.clk(clk),.d(0),.we(0));
//assign O16_I29_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O16_I29_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O16_I29_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O16_I29_R0_C01_rom_inst (.q(O16_I29_R0_C0_SM1 ),.address(input_fmap_29[7:0]),.clock  (clk));
logic [10-1:0] O16_I30_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O16_I30_R0_C01_rom_inst (.q(O16_I30_R0_C0_SM1 ),.address(input_fmap_30[7:0]),.clk(clk),.d(0),.we(0));
//assign O16_I30_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O16_I30_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O16_I30_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O16_I30_R0_C01_rom_inst (.q(O16_I30_R0_C0_SM1 ),.address(input_fmap_30[7:0]),.clock  (clk));
logic [10-1:0] O16_I31_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O16_I31_R0_C01_rom_inst (.q(O16_I31_R0_C0_SM1 ),.address(input_fmap_31[7:0]),.clk(clk),.d(0),.we(0));
//assign O16_I31_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O16_I31_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O16_I31_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O16_I31_R0_C01_rom_inst (.q(O16_I31_R0_C0_SM1 ),.address(input_fmap_31[7:0]),.clock  (clk));
logic [10-1:0] O17_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O17_I0_R0_C01_rom_inst (.q(O17_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O17_I0_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O17_I0_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O17_I0_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O17_I0_R0_C01_rom_inst (.q(O17_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [11-1:0] O17_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O17_I2_R0_C02_rom_inst (.q(O17_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O17_I2_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O17_I2_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O17_I2_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O17_I2_R0_C02_rom_inst (.q(O17_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [11-1:0] O17_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O17_I5_R0_C02_rom_inst (.q(O17_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O17_I5_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O17_I5_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O17_I5_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O17_I5_R0_C02_rom_inst (.q(O17_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [11-1:0] O17_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O17_I7_R0_C02_rom_inst (.q(O17_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O17_I7_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O17_I7_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O17_I7_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O17_I7_R0_C02_rom_inst (.q(O17_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [10-1:0] O17_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O17_I9_R0_C01_rom_inst (.q(O17_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O17_I9_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O17_I9_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O17_I9_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O17_I9_R0_C01_rom_inst (.q(O17_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [10-1:0] O17_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O17_I11_R0_C01_rom_inst (.q(O17_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O17_I11_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O17_I11_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O17_I11_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O17_I11_R0_C01_rom_inst (.q(O17_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [11-1:0] O17_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O17_I12_R0_C02_rom_inst (.q(O17_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O17_I12_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O17_I12_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O17_I12_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O17_I12_R0_C02_rom_inst (.q(O17_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [10-1:0] O17_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O17_I13_R0_C01_rom_inst (.q(O17_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O17_I13_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O17_I13_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O17_I13_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O17_I13_R0_C01_rom_inst (.q(O17_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [11-1:0] O17_I14_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O17_I14_R0_C02_rom_inst (.q(O17_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clk(clk),.d(0),.we(0));
//assign O17_I14_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O17_I14_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O17_I14_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O17_I14_R0_C02_rom_inst (.q(O17_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clock  (clk));
logic [10-1:0] O17_I16_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O17_I16_R0_C01_rom_inst (.q(O17_I16_R0_C0_SM1 ),.address(input_fmap_16[7:0]),.clk(clk),.d(0),.we(0));
//assign O17_I16_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O17_I16_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O17_I16_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O17_I16_R0_C01_rom_inst (.q(O17_I16_R0_C0_SM1 ),.address(input_fmap_16[7:0]),.clock  (clk));
logic [10-1:0] O17_I17_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O17_I17_R0_C01_rom_inst (.q(O17_I17_R0_C0_SM1 ),.address(input_fmap_17[7:0]),.clk(clk),.d(0),.we(0));
//assign O17_I17_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O17_I17_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O17_I17_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O17_I17_R0_C01_rom_inst (.q(O17_I17_R0_C0_SM1 ),.address(input_fmap_17[7:0]),.clock  (clk));
logic [10-1:0] O17_I19_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O17_I19_R0_C01_rom_inst (.q(O17_I19_R0_C0_SM1 ),.address(input_fmap_19[7:0]),.clk(clk),.d(0),.we(0));
//assign O17_I19_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O17_I19_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O17_I19_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O17_I19_R0_C01_rom_inst (.q(O17_I19_R0_C0_SM1 ),.address(input_fmap_19[7:0]),.clock  (clk));
logic [10-1:0] O17_I20_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O17_I20_R0_C01_rom_inst (.q(O17_I20_R0_C0_SM1 ),.address(input_fmap_20[7:0]),.clk(clk),.d(0),.we(0));
//assign O17_I20_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O17_I20_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O17_I20_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O17_I20_R0_C01_rom_inst (.q(O17_I20_R0_C0_SM1 ),.address(input_fmap_20[7:0]),.clock  (clk));
logic [10-1:0] O17_I21_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O17_I21_R0_C01_rom_inst (.q(O17_I21_R0_C0_SM1 ),.address(input_fmap_21[7:0]),.clk(clk),.d(0),.we(0));
//assign O17_I21_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O17_I21_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O17_I21_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O17_I21_R0_C01_rom_inst (.q(O17_I21_R0_C0_SM1 ),.address(input_fmap_21[7:0]),.clock  (clk));
logic [10-1:0] O17_I24_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O17_I24_R0_C01_rom_inst (.q(O17_I24_R0_C0_SM1 ),.address(input_fmap_24[7:0]),.clk(clk),.d(0),.we(0));
//assign O17_I24_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O17_I24_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O17_I24_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O17_I24_R0_C01_rom_inst (.q(O17_I24_R0_C0_SM1 ),.address(input_fmap_24[7:0]),.clock  (clk));
logic [12-1:0] O17_I25_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_pw_O17_I25_R0_C04_rom_inst (.q(O17_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clk(clk),.d(0),.we(0));
//assign O17_I25_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O17_I25_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O17_I25_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_pw_O17_I25_R0_C04_rom_inst (.q(O17_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clock  (clk));
logic [11-1:0] O17_I26_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O17_I26_R0_C02_rom_inst (.q(O17_I26_R0_C0_SM1 ),.address(input_fmap_26[7:0]),.clk(clk),.d(0),.we(0));
//assign O17_I26_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O17_I26_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O17_I26_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O17_I26_R0_C02_rom_inst (.q(O17_I26_R0_C0_SM1 ),.address(input_fmap_26[7:0]),.clock  (clk));
logic [10-1:0] O17_I27_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O17_I27_R0_C01_rom_inst (.q(O17_I27_R0_C0_SM1 ),.address(input_fmap_27[7:0]),.clk(clk),.d(0),.we(0));
//assign O17_I27_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O17_I27_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O17_I27_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O17_I27_R0_C01_rom_inst (.q(O17_I27_R0_C0_SM1 ),.address(input_fmap_27[7:0]),.clock  (clk));
logic [10-1:0] O17_I28_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O17_I28_R0_C01_rom_inst (.q(O17_I28_R0_C0_SM1 ),.address(input_fmap_28[7:0]),.clk(clk),.d(0),.we(0));
//assign O17_I28_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O17_I28_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O17_I28_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O17_I28_R0_C01_rom_inst (.q(O17_I28_R0_C0_SM1 ),.address(input_fmap_28[7:0]),.clock  (clk));
logic [10-1:0] O17_I29_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O17_I29_R0_C01_rom_inst (.q(O17_I29_R0_C0_SM1 ),.address(input_fmap_29[7:0]),.clk(clk),.d(0),.we(0));
//assign O17_I29_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O17_I29_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O17_I29_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O17_I29_R0_C01_rom_inst (.q(O17_I29_R0_C0_SM1 ),.address(input_fmap_29[7:0]),.clock  (clk));
logic [11-1:0] O17_I31_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O17_I31_R0_C02_rom_inst (.q(O17_I31_R0_C0_SM1 ),.address(input_fmap_31[7:0]),.clk(clk),.d(0),.we(0));
//assign O17_I31_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O17_I31_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O17_I31_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O17_I31_R0_C02_rom_inst (.q(O17_I31_R0_C0_SM1 ),.address(input_fmap_31[7:0]),.clock  (clk));
logic [10-1:0] O18_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O18_I2_R0_C01_rom_inst (.q(O18_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O18_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O18_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O18_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O18_I2_R0_C01_rom_inst (.q(O18_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [10-1:0] O18_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O18_I4_R0_C01_rom_inst (.q(O18_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O18_I4_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O18_I4_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O18_I4_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O18_I4_R0_C01_rom_inst (.q(O18_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [10-1:0] O18_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O18_I5_R0_C01_rom_inst (.q(O18_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O18_I5_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O18_I5_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O18_I5_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O18_I5_R0_C01_rom_inst (.q(O18_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [11-1:0] O18_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O18_I6_R0_C02_rom_inst (.q(O18_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O18_I6_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O18_I6_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O18_I6_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O18_I6_R0_C02_rom_inst (.q(O18_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [10-1:0] O18_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O18_I7_R0_C01_rom_inst (.q(O18_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O18_I7_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O18_I7_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O18_I7_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O18_I7_R0_C01_rom_inst (.q(O18_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [10-1:0] O18_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O18_I9_R0_C01_rom_inst (.q(O18_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O18_I9_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O18_I9_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O18_I9_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O18_I9_R0_C01_rom_inst (.q(O18_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [10-1:0] O18_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O18_I11_R0_C01_rom_inst (.q(O18_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O18_I11_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O18_I11_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O18_I11_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O18_I11_R0_C01_rom_inst (.q(O18_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [10-1:0] O18_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O18_I12_R0_C01_rom_inst (.q(O18_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O18_I12_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O18_I12_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O18_I12_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O18_I12_R0_C01_rom_inst (.q(O18_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [10-1:0] O18_I17_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O18_I17_R0_C01_rom_inst (.q(O18_I17_R0_C0_SM1 ),.address(input_fmap_17[7:0]),.clk(clk),.d(0),.we(0));
//assign O18_I17_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O18_I17_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O18_I17_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O18_I17_R0_C01_rom_inst (.q(O18_I17_R0_C0_SM1 ),.address(input_fmap_17[7:0]),.clock  (clk));
logic [10-1:0] O18_I19_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O18_I19_R0_C01_rom_inst (.q(O18_I19_R0_C0_SM1 ),.address(input_fmap_19[7:0]),.clk(clk),.d(0),.we(0));
//assign O18_I19_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O18_I19_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O18_I19_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O18_I19_R0_C01_rom_inst (.q(O18_I19_R0_C0_SM1 ),.address(input_fmap_19[7:0]),.clock  (clk));
logic [10-1:0] O18_I21_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O18_I21_R0_C01_rom_inst (.q(O18_I21_R0_C0_SM1 ),.address(input_fmap_21[7:0]),.clk(clk),.d(0),.we(0));
//assign O18_I21_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O18_I21_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O18_I21_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O18_I21_R0_C01_rom_inst (.q(O18_I21_R0_C0_SM1 ),.address(input_fmap_21[7:0]),.clock  (clk));
logic [10-1:0] O18_I22_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O18_I22_R0_C01_rom_inst (.q(O18_I22_R0_C0_SM1 ),.address(input_fmap_22[7:0]),.clk(clk),.d(0),.we(0));
//assign O18_I22_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O18_I22_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O18_I22_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O18_I22_R0_C01_rom_inst (.q(O18_I22_R0_C0_SM1 ),.address(input_fmap_22[7:0]),.clock  (clk));
logic [10-1:0] O18_I23_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O18_I23_R0_C01_rom_inst (.q(O18_I23_R0_C0_SM1 ),.address(input_fmap_23[7:0]),.clk(clk),.d(0),.we(0));
//assign O18_I23_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O18_I23_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O18_I23_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O18_I23_R0_C01_rom_inst (.q(O18_I23_R0_C0_SM1 ),.address(input_fmap_23[7:0]),.clock  (clk));
logic [10-1:0] O18_I26_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O18_I26_R0_C01_rom_inst (.q(O18_I26_R0_C0_SM1 ),.address(input_fmap_26[7:0]),.clk(clk),.d(0),.we(0));
//assign O18_I26_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O18_I26_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O18_I26_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O18_I26_R0_C01_rom_inst (.q(O18_I26_R0_C0_SM1 ),.address(input_fmap_26[7:0]),.clock  (clk));
logic [10-1:0] O18_I28_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O18_I28_R0_C01_rom_inst (.q(O18_I28_R0_C0_SM1 ),.address(input_fmap_28[7:0]),.clk(clk),.d(0),.we(0));
//assign O18_I28_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O18_I28_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O18_I28_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O18_I28_R0_C01_rom_inst (.q(O18_I28_R0_C0_SM1 ),.address(input_fmap_28[7:0]),.clock  (clk));
logic [10-1:0] O19_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O19_I4_R0_C01_rom_inst (.q(O19_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O19_I4_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O19_I4_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O19_I4_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O19_I4_R0_C01_rom_inst (.q(O19_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [10-1:0] O19_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O19_I7_R0_C01_rom_inst (.q(O19_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O19_I7_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O19_I7_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O19_I7_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O19_I7_R0_C01_rom_inst (.q(O19_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [10-1:0] O19_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O19_I9_R0_C01_rom_inst (.q(O19_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O19_I9_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O19_I9_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O19_I9_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O19_I9_R0_C01_rom_inst (.q(O19_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [10-1:0] O19_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O19_I11_R0_C01_rom_inst (.q(O19_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O19_I11_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O19_I11_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O19_I11_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O19_I11_R0_C01_rom_inst (.q(O19_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [10-1:0] O19_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O19_I12_R0_C01_rom_inst (.q(O19_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O19_I12_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O19_I12_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O19_I12_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O19_I12_R0_C01_rom_inst (.q(O19_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [10-1:0] O19_I20_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O19_I20_R0_C01_rom_inst (.q(O19_I20_R0_C0_SM1 ),.address(input_fmap_20[7:0]),.clk(clk),.d(0),.we(0));
//assign O19_I20_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O19_I20_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O19_I20_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O19_I20_R0_C01_rom_inst (.q(O19_I20_R0_C0_SM1 ),.address(input_fmap_20[7:0]),.clock  (clk));
logic [10-1:0] O19_I23_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O19_I23_R0_C01_rom_inst (.q(O19_I23_R0_C0_SM1 ),.address(input_fmap_23[7:0]),.clk(clk),.d(0),.we(0));
//assign O19_I23_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O19_I23_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O19_I23_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O19_I23_R0_C01_rom_inst (.q(O19_I23_R0_C0_SM1 ),.address(input_fmap_23[7:0]),.clock  (clk));
logic [10-1:0] O19_I24_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O19_I24_R0_C01_rom_inst (.q(O19_I24_R0_C0_SM1 ),.address(input_fmap_24[7:0]),.clk(clk),.d(0),.we(0));
//assign O19_I24_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O19_I24_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O19_I24_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O19_I24_R0_C01_rom_inst (.q(O19_I24_R0_C0_SM1 ),.address(input_fmap_24[7:0]),.clock  (clk));
logic [10-1:0] O19_I26_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O19_I26_R0_C01_rom_inst (.q(O19_I26_R0_C0_SM1 ),.address(input_fmap_26[7:0]),.clk(clk),.d(0),.we(0));
//assign O19_I26_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O19_I26_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O19_I26_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O19_I26_R0_C01_rom_inst (.q(O19_I26_R0_C0_SM1 ),.address(input_fmap_26[7:0]),.clock  (clk));
logic [10-1:0] O19_I31_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O19_I31_R0_C01_rom_inst (.q(O19_I31_R0_C0_SM1 ),.address(input_fmap_31[7:0]),.clk(clk),.d(0),.we(0));
//assign O19_I31_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O19_I31_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O19_I31_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O19_I31_R0_C01_rom_inst (.q(O19_I31_R0_C0_SM1 ),.address(input_fmap_31[7:0]),.clock  (clk));
logic [10-1:0] O20_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O20_I3_R0_C01_rom_inst (.q(O20_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O20_I3_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O20_I3_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O20_I3_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O20_I3_R0_C01_rom_inst (.q(O20_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [10-1:0] O20_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O20_I6_R0_C01_rom_inst (.q(O20_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O20_I6_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O20_I6_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O20_I6_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O20_I6_R0_C01_rom_inst (.q(O20_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [10-1:0] O20_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O20_I7_R0_C01_rom_inst (.q(O20_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O20_I7_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O20_I7_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O20_I7_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O20_I7_R0_C01_rom_inst (.q(O20_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [10-1:0] O20_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O20_I8_R0_C01_rom_inst (.q(O20_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O20_I8_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O20_I8_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O20_I8_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O20_I8_R0_C01_rom_inst (.q(O20_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [10-1:0] O20_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O20_I9_R0_C01_rom_inst (.q(O20_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O20_I9_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O20_I9_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O20_I9_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O20_I9_R0_C01_rom_inst (.q(O20_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [10-1:0] O20_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O20_I13_R0_C01_rom_inst (.q(O20_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O20_I13_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O20_I13_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O20_I13_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O20_I13_R0_C01_rom_inst (.q(O20_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [10-1:0] O20_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O20_I15_R0_C01_rom_inst (.q(O20_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O20_I15_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O20_I15_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O20_I15_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O20_I15_R0_C01_rom_inst (.q(O20_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [11-1:0] O20_I17_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O20_I17_R0_C02_rom_inst (.q(O20_I17_R0_C0_SM1 ),.address(input_fmap_17[7:0]),.clk(clk),.d(0),.we(0));
//assign O20_I17_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O20_I17_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O20_I17_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O20_I17_R0_C02_rom_inst (.q(O20_I17_R0_C0_SM1 ),.address(input_fmap_17[7:0]),.clock  (clk));
logic [10-1:0] O20_I18_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O20_I18_R0_C01_rom_inst (.q(O20_I18_R0_C0_SM1 ),.address(input_fmap_18[7:0]),.clk(clk),.d(0),.we(0));
//assign O20_I18_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O20_I18_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O20_I18_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O20_I18_R0_C01_rom_inst (.q(O20_I18_R0_C0_SM1 ),.address(input_fmap_18[7:0]),.clock  (clk));
logic [10-1:0] O20_I21_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O20_I21_R0_C01_rom_inst (.q(O20_I21_R0_C0_SM1 ),.address(input_fmap_21[7:0]),.clk(clk),.d(0),.we(0));
//assign O20_I21_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O20_I21_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O20_I21_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O20_I21_R0_C01_rom_inst (.q(O20_I21_R0_C0_SM1 ),.address(input_fmap_21[7:0]),.clock  (clk));
logic [10-1:0] O20_I22_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O20_I22_R0_C01_rom_inst (.q(O20_I22_R0_C0_SM1 ),.address(input_fmap_22[7:0]),.clk(clk),.d(0),.we(0));
//assign O20_I22_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O20_I22_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O20_I22_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O20_I22_R0_C01_rom_inst (.q(O20_I22_R0_C0_SM1 ),.address(input_fmap_22[7:0]),.clock  (clk));
logic [10-1:0] O20_I23_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O20_I23_R0_C01_rom_inst (.q(O20_I23_R0_C0_SM1 ),.address(input_fmap_23[7:0]),.clk(clk),.d(0),.we(0));
//assign O20_I23_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O20_I23_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O20_I23_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O20_I23_R0_C01_rom_inst (.q(O20_I23_R0_C0_SM1 ),.address(input_fmap_23[7:0]),.clock  (clk));
logic [11-1:0] O20_I24_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O20_I24_R0_C02_rom_inst (.q(O20_I24_R0_C0_SM1 ),.address(input_fmap_24[7:0]),.clk(clk),.d(0),.we(0));
//assign O20_I24_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O20_I24_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O20_I24_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O20_I24_R0_C02_rom_inst (.q(O20_I24_R0_C0_SM1 ),.address(input_fmap_24[7:0]),.clock  (clk));
logic [11-1:0] O20_I25_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O20_I25_R0_C03_rom_inst (.q(O20_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clk(clk),.d(0),.we(0));
//assign O20_I25_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O20_I25_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O20_I25_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O20_I25_R0_C03_rom_inst (.q(O20_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clock  (clk));
logic [10-1:0] O20_I28_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O20_I28_R0_C01_rom_inst (.q(O20_I28_R0_C0_SM1 ),.address(input_fmap_28[7:0]),.clk(clk),.d(0),.we(0));
//assign O20_I28_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O20_I28_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O20_I28_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O20_I28_R0_C01_rom_inst (.q(O20_I28_R0_C0_SM1 ),.address(input_fmap_28[7:0]),.clock  (clk));
logic [10-1:0] O20_I30_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O20_I30_R0_C01_rom_inst (.q(O20_I30_R0_C0_SM1 ),.address(input_fmap_30[7:0]),.clk(clk),.d(0),.we(0));
//assign O20_I30_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O20_I30_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O20_I30_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O20_I30_R0_C01_rom_inst (.q(O20_I30_R0_C0_SM1 ),.address(input_fmap_30[7:0]),.clock  (clk));
logic [10-1:0] O20_I31_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O20_I31_R0_C01_rom_inst (.q(O20_I31_R0_C0_SM1 ),.address(input_fmap_31[7:0]),.clk(clk),.d(0),.we(0));
//assign O20_I31_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O20_I31_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O20_I31_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O20_I31_R0_C01_rom_inst (.q(O20_I31_R0_C0_SM1 ),.address(input_fmap_31[7:0]),.clock  (clk));
logic [10-1:0] O21_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O21_I0_R0_C01_rom_inst (.q(O21_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O21_I0_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O21_I0_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O21_I0_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O21_I0_R0_C01_rom_inst (.q(O21_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [12-1:0] O21_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_pw_O21_I1_R0_C06_rom_inst (.q(O21_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O21_I1_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O21_I1_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O21_I1_R0_C06_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_pw_O21_I1_R0_C06_rom_inst (.q(O21_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [11-1:0] O21_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O21_I2_R0_C02_rom_inst (.q(O21_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O21_I2_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O21_I2_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O21_I2_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O21_I2_R0_C02_rom_inst (.q(O21_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [10-1:0] O21_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O21_I3_R0_C01_rom_inst (.q(O21_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O21_I3_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O21_I3_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O21_I3_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O21_I3_R0_C01_rom_inst (.q(O21_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [10-1:0] O21_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O21_I4_R0_C01_rom_inst (.q(O21_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O21_I4_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O21_I4_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O21_I4_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O21_I4_R0_C01_rom_inst (.q(O21_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [11-1:0] O21_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O21_I5_R0_C03_rom_inst (.q(O21_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O21_I5_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O21_I5_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O21_I5_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O21_I5_R0_C03_rom_inst (.q(O21_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [11-1:0] O21_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O21_I6_R0_C02_rom_inst (.q(O21_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O21_I6_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O21_I6_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O21_I6_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O21_I6_R0_C02_rom_inst (.q(O21_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [10-1:0] O21_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O21_I7_R0_C01_rom_inst (.q(O21_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O21_I7_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O21_I7_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O21_I7_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O21_I7_R0_C01_rom_inst (.q(O21_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [12-1:0] O21_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_pw_O21_I8_R0_C04_rom_inst (.q(O21_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O21_I8_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O21_I8_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O21_I8_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_pw_O21_I8_R0_C04_rom_inst (.q(O21_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [11-1:0] O21_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O21_I9_R0_C02_rom_inst (.q(O21_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O21_I9_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O21_I9_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O21_I9_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O21_I9_R0_C02_rom_inst (.q(O21_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [10-1:0] O21_I10_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O21_I10_R0_C01_rom_inst (.q(O21_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clk(clk),.d(0),.we(0));
//assign O21_I10_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O21_I10_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O21_I10_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O21_I10_R0_C01_rom_inst (.q(O21_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clock  (clk));
logic [10-1:0] O21_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O21_I13_R0_C01_rom_inst (.q(O21_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O21_I13_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O21_I13_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O21_I13_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O21_I13_R0_C01_rom_inst (.q(O21_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [10-1:0] O21_I16_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O21_I16_R0_C01_rom_inst (.q(O21_I16_R0_C0_SM1 ),.address(input_fmap_16[7:0]),.clk(clk),.d(0),.we(0));
//assign O21_I16_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O21_I16_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O21_I16_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O21_I16_R0_C01_rom_inst (.q(O21_I16_R0_C0_SM1 ),.address(input_fmap_16[7:0]),.clock  (clk));
logic [11-1:0] O21_I17_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O21_I17_R0_C03_rom_inst (.q(O21_I17_R0_C0_SM1 ),.address(input_fmap_17[7:0]),.clk(clk),.d(0),.we(0));
//assign O21_I17_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O21_I17_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O21_I17_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O21_I17_R0_C03_rom_inst (.q(O21_I17_R0_C0_SM1 ),.address(input_fmap_17[7:0]),.clock  (clk));
logic [10-1:0] O21_I18_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O21_I18_R0_C01_rom_inst (.q(O21_I18_R0_C0_SM1 ),.address(input_fmap_18[7:0]),.clk(clk),.d(0),.we(0));
//assign O21_I18_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O21_I18_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O21_I18_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O21_I18_R0_C01_rom_inst (.q(O21_I18_R0_C0_SM1 ),.address(input_fmap_18[7:0]),.clock  (clk));
logic [11-1:0] O21_I19_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O21_I19_R0_C02_rom_inst (.q(O21_I19_R0_C0_SM1 ),.address(input_fmap_19[7:0]),.clk(clk),.d(0),.we(0));
//assign O21_I19_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O21_I19_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O21_I19_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O21_I19_R0_C02_rom_inst (.q(O21_I19_R0_C0_SM1 ),.address(input_fmap_19[7:0]),.clock  (clk));
logic [11-1:0] O21_I21_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O21_I21_R0_C03_rom_inst (.q(O21_I21_R0_C0_SM1 ),.address(input_fmap_21[7:0]),.clk(clk),.d(0),.we(0));
//assign O21_I21_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O21_I21_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O21_I21_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O21_I21_R0_C03_rom_inst (.q(O21_I21_R0_C0_SM1 ),.address(input_fmap_21[7:0]),.clock  (clk));
logic [12-1:0] O21_I22_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_pw_O21_I22_R0_C04_rom_inst (.q(O21_I22_R0_C0_SM1 ),.address(input_fmap_22[7:0]),.clk(clk),.d(0),.we(0));
//assign O21_I22_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O21_I22_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O21_I22_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_pw_O21_I22_R0_C04_rom_inst (.q(O21_I22_R0_C0_SM1 ),.address(input_fmap_22[7:0]),.clock  (clk));
logic [11-1:0] O21_I24_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O21_I24_R0_C03_rom_inst (.q(O21_I24_R0_C0_SM1 ),.address(input_fmap_24[7:0]),.clk(clk),.d(0),.we(0));
//assign O21_I24_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O21_I24_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O21_I24_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O21_I24_R0_C03_rom_inst (.q(O21_I24_R0_C0_SM1 ),.address(input_fmap_24[7:0]),.clock  (clk));
logic [11-1:0] O21_I25_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O21_I25_R0_C03_rom_inst (.q(O21_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clk(clk),.d(0),.we(0));
//assign O21_I25_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O21_I25_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O21_I25_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O21_I25_R0_C03_rom_inst (.q(O21_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clock  (clk));
logic [11-1:0] O21_I27_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O21_I27_R0_C02_rom_inst (.q(O21_I27_R0_C0_SM1 ),.address(input_fmap_27[7:0]),.clk(clk),.d(0),.we(0));
//assign O21_I27_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O21_I27_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O21_I27_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O21_I27_R0_C02_rom_inst (.q(O21_I27_R0_C0_SM1 ),.address(input_fmap_27[7:0]),.clock  (clk));
logic [11-1:0] O21_I28_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O21_I28_R0_C02_rom_inst (.q(O21_I28_R0_C0_SM1 ),.address(input_fmap_28[7:0]),.clk(clk),.d(0),.we(0));
//assign O21_I28_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O21_I28_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O21_I28_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O21_I28_R0_C02_rom_inst (.q(O21_I28_R0_C0_SM1 ),.address(input_fmap_28[7:0]),.clock  (clk));
logic [11-1:0] O21_I29_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O21_I29_R0_C03_rom_inst (.q(O21_I29_R0_C0_SM1 ),.address(input_fmap_29[7:0]),.clk(clk),.d(0),.we(0));
//assign O21_I29_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O21_I29_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O21_I29_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O21_I29_R0_C03_rom_inst (.q(O21_I29_R0_C0_SM1 ),.address(input_fmap_29[7:0]),.clock  (clk));
logic [11-1:0] O21_I30_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O21_I30_R0_C03_rom_inst (.q(O21_I30_R0_C0_SM1 ),.address(input_fmap_30[7:0]),.clk(clk),.d(0),.we(0));
//assign O21_I30_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O21_I30_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O21_I30_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O21_I30_R0_C03_rom_inst (.q(O21_I30_R0_C0_SM1 ),.address(input_fmap_30[7:0]),.clock  (clk));
logic [10-1:0] O21_I31_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O21_I31_R0_C01_rom_inst (.q(O21_I31_R0_C0_SM1 ),.address(input_fmap_31[7:0]),.clk(clk),.d(0),.we(0));
//assign O21_I31_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O21_I31_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O21_I31_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O21_I31_R0_C01_rom_inst (.q(O21_I31_R0_C0_SM1 ),.address(input_fmap_31[7:0]),.clock  (clk));
logic [10-1:0] O22_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O22_I2_R0_C01_rom_inst (.q(O22_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O22_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O22_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O22_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O22_I2_R0_C01_rom_inst (.q(O22_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [11-1:0] O22_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O22_I3_R0_C02_rom_inst (.q(O22_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O22_I3_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O22_I3_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O22_I3_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O22_I3_R0_C02_rom_inst (.q(O22_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [10-1:0] O22_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O22_I6_R0_C01_rom_inst (.q(O22_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O22_I6_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O22_I6_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O22_I6_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O22_I6_R0_C01_rom_inst (.q(O22_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [11-1:0] O22_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O22_I7_R0_C02_rom_inst (.q(O22_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O22_I7_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O22_I7_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O22_I7_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O22_I7_R0_C02_rom_inst (.q(O22_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [11-1:0] O22_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O22_I8_R0_C02_rom_inst (.q(O22_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O22_I8_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O22_I8_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O22_I8_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O22_I8_R0_C02_rom_inst (.q(O22_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [11-1:0] O22_I10_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O22_I10_R0_C02_rom_inst (.q(O22_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clk(clk),.d(0),.we(0));
//assign O22_I10_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O22_I10_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O22_I10_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O22_I10_R0_C02_rom_inst (.q(O22_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clock  (clk));
logic [10-1:0] O22_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O22_I12_R0_C01_rom_inst (.q(O22_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O22_I12_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O22_I12_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O22_I12_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O22_I12_R0_C01_rom_inst (.q(O22_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [11-1:0] O22_I14_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O22_I14_R0_C03_rom_inst (.q(O22_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clk(clk),.d(0),.we(0));
//assign O22_I14_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O22_I14_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O22_I14_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O22_I14_R0_C03_rom_inst (.q(O22_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clock  (clk));
logic [10-1:0] O22_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O22_I15_R0_C01_rom_inst (.q(O22_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O22_I15_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O22_I15_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O22_I15_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O22_I15_R0_C01_rom_inst (.q(O22_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [10-1:0] O22_I17_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O22_I17_R0_C01_rom_inst (.q(O22_I17_R0_C0_SM1 ),.address(input_fmap_17[7:0]),.clk(clk),.d(0),.we(0));
//assign O22_I17_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O22_I17_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O22_I17_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O22_I17_R0_C01_rom_inst (.q(O22_I17_R0_C0_SM1 ),.address(input_fmap_17[7:0]),.clock  (clk));
logic [12-1:0] O22_I18_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_pw_O22_I18_R0_C06_rom_inst (.q(O22_I18_R0_C0_SM1 ),.address(input_fmap_18[7:0]),.clk(clk),.d(0),.we(0));
//assign O22_I18_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O22_I18_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O22_I18_R0_C06_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_pw_O22_I18_R0_C06_rom_inst (.q(O22_I18_R0_C0_SM1 ),.address(input_fmap_18[7:0]),.clock  (clk));
logic [10-1:0] O22_I20_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O22_I20_R0_C01_rom_inst (.q(O22_I20_R0_C0_SM1 ),.address(input_fmap_20[7:0]),.clk(clk),.d(0),.we(0));
//assign O22_I20_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O22_I20_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O22_I20_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O22_I20_R0_C01_rom_inst (.q(O22_I20_R0_C0_SM1 ),.address(input_fmap_20[7:0]),.clock  (clk));
logic [11-1:0] O22_I22_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O22_I22_R0_C03_rom_inst (.q(O22_I22_R0_C0_SM1 ),.address(input_fmap_22[7:0]),.clk(clk),.d(0),.we(0));
//assign O22_I22_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O22_I22_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O22_I22_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O22_I22_R0_C03_rom_inst (.q(O22_I22_R0_C0_SM1 ),.address(input_fmap_22[7:0]),.clock  (clk));
logic [10-1:0] O22_I23_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O22_I23_R0_C01_rom_inst (.q(O22_I23_R0_C0_SM1 ),.address(input_fmap_23[7:0]),.clk(clk),.d(0),.we(0));
//assign O22_I23_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O22_I23_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O22_I23_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O22_I23_R0_C01_rom_inst (.q(O22_I23_R0_C0_SM1 ),.address(input_fmap_23[7:0]),.clock  (clk));
logic [10-1:0] O22_I25_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O22_I25_R0_C01_rom_inst (.q(O22_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clk(clk),.d(0),.we(0));
//assign O22_I25_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O22_I25_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O22_I25_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O22_I25_R0_C01_rom_inst (.q(O22_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clock  (clk));
logic [11-1:0] O22_I27_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O22_I27_R0_C03_rom_inst (.q(O22_I27_R0_C0_SM1 ),.address(input_fmap_27[7:0]),.clk(clk),.d(0),.we(0));
//assign O22_I27_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O22_I27_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O22_I27_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O22_I27_R0_C03_rom_inst (.q(O22_I27_R0_C0_SM1 ),.address(input_fmap_27[7:0]),.clock  (clk));
logic [10-1:0] O22_I28_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O22_I28_R0_C01_rom_inst (.q(O22_I28_R0_C0_SM1 ),.address(input_fmap_28[7:0]),.clk(clk),.d(0),.we(0));
//assign O22_I28_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O22_I28_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O22_I28_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O22_I28_R0_C01_rom_inst (.q(O22_I28_R0_C0_SM1 ),.address(input_fmap_28[7:0]),.clock  (clk));
logic [12-1:0] O22_I29_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_pw_O22_I29_R0_C04_rom_inst (.q(O22_I29_R0_C0_SM1 ),.address(input_fmap_29[7:0]),.clk(clk),.d(0),.we(0));
//assign O22_I29_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O22_I29_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O22_I29_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_pw_O22_I29_R0_C04_rom_inst (.q(O22_I29_R0_C0_SM1 ),.address(input_fmap_29[7:0]),.clock  (clk));
logic [10-1:0] O22_I30_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O22_I30_R0_C01_rom_inst (.q(O22_I30_R0_C0_SM1 ),.address(input_fmap_30[7:0]),.clk(clk),.d(0),.we(0));
//assign O22_I30_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O22_I30_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O22_I30_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O22_I30_R0_C01_rom_inst (.q(O22_I30_R0_C0_SM1 ),.address(input_fmap_30[7:0]),.clock  (clk));
logic [10-1:0] O23_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O23_I3_R0_C01_rom_inst (.q(O23_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O23_I3_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O23_I3_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O23_I3_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O23_I3_R0_C01_rom_inst (.q(O23_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [10-1:0] O23_I10_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O23_I10_R0_C01_rom_inst (.q(O23_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clk(clk),.d(0),.we(0));
//assign O23_I10_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O23_I10_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O23_I10_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O23_I10_R0_C01_rom_inst (.q(O23_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clock  (clk));
logic [11-1:0] O23_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O23_I15_R0_C02_rom_inst (.q(O23_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O23_I15_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O23_I15_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O23_I15_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O23_I15_R0_C02_rom_inst (.q(O23_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [10-1:0] O23_I17_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O23_I17_R0_C01_rom_inst (.q(O23_I17_R0_C0_SM1 ),.address(input_fmap_17[7:0]),.clk(clk),.d(0),.we(0));
//assign O23_I17_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O23_I17_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O23_I17_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O23_I17_R0_C01_rom_inst (.q(O23_I17_R0_C0_SM1 ),.address(input_fmap_17[7:0]),.clock  (clk));
logic [12-1:0] O23_I18_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_pw_O23_I18_R0_C05_rom_inst (.q(O23_I18_R0_C0_SM1 ),.address(input_fmap_18[7:0]),.clk(clk),.d(0),.we(0));
//assign O23_I18_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O23_I18_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O23_I18_R0_C05_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_pw_O23_I18_R0_C05_rom_inst (.q(O23_I18_R0_C0_SM1 ),.address(input_fmap_18[7:0]),.clock  (clk));
logic [10-1:0] O23_I22_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O23_I22_R0_C01_rom_inst (.q(O23_I22_R0_C0_SM1 ),.address(input_fmap_22[7:0]),.clk(clk),.d(0),.we(0));
//assign O23_I22_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O23_I22_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O23_I22_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O23_I22_R0_C01_rom_inst (.q(O23_I22_R0_C0_SM1 ),.address(input_fmap_22[7:0]),.clock  (clk));
logic [10-1:0] O23_I25_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O23_I25_R0_C01_rom_inst (.q(O23_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clk(clk),.d(0),.we(0));
//assign O23_I25_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O23_I25_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O23_I25_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O23_I25_R0_C01_rom_inst (.q(O23_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clock  (clk));
logic [12-1:0] O24_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_pw_O24_I0_R0_C04_rom_inst (.q(O24_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O24_I0_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O24_I0_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O24_I0_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_pw_O24_I0_R0_C04_rom_inst (.q(O24_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [10-1:0] O24_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O24_I1_R0_C01_rom_inst (.q(O24_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O24_I1_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O24_I1_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O24_I1_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O24_I1_R0_C01_rom_inst (.q(O24_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [10-1:0] O24_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O24_I2_R0_C01_rom_inst (.q(O24_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O24_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O24_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O24_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O24_I2_R0_C01_rom_inst (.q(O24_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [10-1:0] O24_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O24_I8_R0_C01_rom_inst (.q(O24_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O24_I8_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O24_I8_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O24_I8_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O24_I8_R0_C01_rom_inst (.q(O24_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [10-1:0] O24_I10_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O24_I10_R0_C01_rom_inst (.q(O24_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clk(clk),.d(0),.we(0));
//assign O24_I10_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O24_I10_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O24_I10_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O24_I10_R0_C01_rom_inst (.q(O24_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clock  (clk));
logic [12-1:0] O24_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_pw_O24_I13_R0_C04_rom_inst (.q(O24_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O24_I13_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O24_I13_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O24_I13_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_pw_O24_I13_R0_C04_rom_inst (.q(O24_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [10-1:0] O24_I14_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O24_I14_R0_C01_rom_inst (.q(O24_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clk(clk),.d(0),.we(0));
//assign O24_I14_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O24_I14_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O24_I14_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O24_I14_R0_C01_rom_inst (.q(O24_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clock  (clk));
logic [10-1:0] O24_I17_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O24_I17_R0_C01_rom_inst (.q(O24_I17_R0_C0_SM1 ),.address(input_fmap_17[7:0]),.clk(clk),.d(0),.we(0));
//assign O24_I17_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O24_I17_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O24_I17_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O24_I17_R0_C01_rom_inst (.q(O24_I17_R0_C0_SM1 ),.address(input_fmap_17[7:0]),.clock  (clk));
logic [10-1:0] O24_I23_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O24_I23_R0_C01_rom_inst (.q(O24_I23_R0_C0_SM1 ),.address(input_fmap_23[7:0]),.clk(clk),.d(0),.we(0));
//assign O24_I23_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O24_I23_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O24_I23_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O24_I23_R0_C01_rom_inst (.q(O24_I23_R0_C0_SM1 ),.address(input_fmap_23[7:0]),.clock  (clk));
logic [10-1:0] O24_I25_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O24_I25_R0_C01_rom_inst (.q(O24_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clk(clk),.d(0),.we(0));
//assign O24_I25_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O24_I25_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O24_I25_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O24_I25_R0_C01_rom_inst (.q(O24_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clock  (clk));
logic [10-1:0] O24_I27_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O24_I27_R0_C01_rom_inst (.q(O24_I27_R0_C0_SM1 ),.address(input_fmap_27[7:0]),.clk(clk),.d(0),.we(0));
//assign O24_I27_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O24_I27_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O24_I27_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O24_I27_R0_C01_rom_inst (.q(O24_I27_R0_C0_SM1 ),.address(input_fmap_27[7:0]),.clock  (clk));
logic [10-1:0] O24_I30_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O24_I30_R0_C01_rom_inst (.q(O24_I30_R0_C0_SM1 ),.address(input_fmap_30[7:0]),.clk(clk),.d(0),.we(0));
//assign O24_I30_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O24_I30_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O24_I30_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O24_I30_R0_C01_rom_inst (.q(O24_I30_R0_C0_SM1 ),.address(input_fmap_30[7:0]),.clock  (clk));
logic [11-1:0] O25_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O25_I1_R0_C02_rom_inst (.q(O25_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O25_I1_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O25_I1_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O25_I1_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O25_I1_R0_C02_rom_inst (.q(O25_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [10-1:0] O25_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O25_I2_R0_C01_rom_inst (.q(O25_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O25_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O25_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O25_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O25_I2_R0_C01_rom_inst (.q(O25_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [10-1:0] O25_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O25_I7_R0_C01_rom_inst (.q(O25_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O25_I7_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O25_I7_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O25_I7_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O25_I7_R0_C01_rom_inst (.q(O25_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [10-1:0] O25_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O25_I9_R0_C01_rom_inst (.q(O25_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O25_I9_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O25_I9_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O25_I9_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O25_I9_R0_C01_rom_inst (.q(O25_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [10-1:0] O25_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O25_I12_R0_C01_rom_inst (.q(O25_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O25_I12_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O25_I12_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O25_I12_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O25_I12_R0_C01_rom_inst (.q(O25_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [10-1:0] O25_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O25_I13_R0_C01_rom_inst (.q(O25_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O25_I13_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O25_I13_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O25_I13_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O25_I13_R0_C01_rom_inst (.q(O25_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [10-1:0] O25_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O25_I15_R0_C01_rom_inst (.q(O25_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O25_I15_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O25_I15_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O25_I15_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O25_I15_R0_C01_rom_inst (.q(O25_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [10-1:0] O25_I17_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O25_I17_R0_C01_rom_inst (.q(O25_I17_R0_C0_SM1 ),.address(input_fmap_17[7:0]),.clk(clk),.d(0),.we(0));
//assign O25_I17_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O25_I17_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O25_I17_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O25_I17_R0_C01_rom_inst (.q(O25_I17_R0_C0_SM1 ),.address(input_fmap_17[7:0]),.clock  (clk));
logic [10-1:0] O25_I20_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O25_I20_R0_C01_rom_inst (.q(O25_I20_R0_C0_SM1 ),.address(input_fmap_20[7:0]),.clk(clk),.d(0),.we(0));
//assign O25_I20_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O25_I20_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O25_I20_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O25_I20_R0_C01_rom_inst (.q(O25_I20_R0_C0_SM1 ),.address(input_fmap_20[7:0]),.clock  (clk));
logic [10-1:0] O25_I25_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O25_I25_R0_C01_rom_inst (.q(O25_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clk(clk),.d(0),.we(0));
//assign O25_I25_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O25_I25_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O25_I25_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O25_I25_R0_C01_rom_inst (.q(O25_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clock  (clk));
logic [10-1:0] O25_I27_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O25_I27_R0_C01_rom_inst (.q(O25_I27_R0_C0_SM1 ),.address(input_fmap_27[7:0]),.clk(clk),.d(0),.we(0));
//assign O25_I27_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O25_I27_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O25_I27_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O25_I27_R0_C01_rom_inst (.q(O25_I27_R0_C0_SM1 ),.address(input_fmap_27[7:0]),.clock  (clk));
logic [10-1:0] O25_I28_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O25_I28_R0_C01_rom_inst (.q(O25_I28_R0_C0_SM1 ),.address(input_fmap_28[7:0]),.clk(clk),.d(0),.we(0));
//assign O25_I28_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O25_I28_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O25_I28_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O25_I28_R0_C01_rom_inst (.q(O25_I28_R0_C0_SM1 ),.address(input_fmap_28[7:0]),.clock  (clk));
logic [10-1:0] O26_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O26_I0_R0_C01_rom_inst (.q(O26_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O26_I0_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O26_I0_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O26_I0_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O26_I0_R0_C01_rom_inst (.q(O26_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [10-1:0] O26_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O26_I2_R0_C01_rom_inst (.q(O26_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O26_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O26_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O26_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O26_I2_R0_C01_rom_inst (.q(O26_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [10-1:0] O26_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O26_I3_R0_C01_rom_inst (.q(O26_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O26_I3_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O26_I3_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O26_I3_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O26_I3_R0_C01_rom_inst (.q(O26_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [10-1:0] O26_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O26_I4_R0_C01_rom_inst (.q(O26_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O26_I4_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O26_I4_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O26_I4_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O26_I4_R0_C01_rom_inst (.q(O26_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [10-1:0] O26_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O26_I8_R0_C01_rom_inst (.q(O26_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O26_I8_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O26_I8_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O26_I8_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O26_I8_R0_C01_rom_inst (.q(O26_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [10-1:0] O26_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O26_I9_R0_C01_rom_inst (.q(O26_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O26_I9_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O26_I9_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O26_I9_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O26_I9_R0_C01_rom_inst (.q(O26_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [10-1:0] O26_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O26_I11_R0_C01_rom_inst (.q(O26_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O26_I11_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O26_I11_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O26_I11_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O26_I11_R0_C01_rom_inst (.q(O26_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [10-1:0] O26_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O26_I12_R0_C01_rom_inst (.q(O26_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O26_I12_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O26_I12_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O26_I12_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O26_I12_R0_C01_rom_inst (.q(O26_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [10-1:0] O26_I16_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O26_I16_R0_C01_rom_inst (.q(O26_I16_R0_C0_SM1 ),.address(input_fmap_16[7:0]),.clk(clk),.d(0),.we(0));
//assign O26_I16_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O26_I16_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O26_I16_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O26_I16_R0_C01_rom_inst (.q(O26_I16_R0_C0_SM1 ),.address(input_fmap_16[7:0]),.clock  (clk));
logic [10-1:0] O26_I17_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O26_I17_R0_C01_rom_inst (.q(O26_I17_R0_C0_SM1 ),.address(input_fmap_17[7:0]),.clk(clk),.d(0),.we(0));
//assign O26_I17_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O26_I17_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O26_I17_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O26_I17_R0_C01_rom_inst (.q(O26_I17_R0_C0_SM1 ),.address(input_fmap_17[7:0]),.clock  (clk));
logic [11-1:0] O26_I19_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O26_I19_R0_C02_rom_inst (.q(O26_I19_R0_C0_SM1 ),.address(input_fmap_19[7:0]),.clk(clk),.d(0),.we(0));
//assign O26_I19_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O26_I19_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O26_I19_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O26_I19_R0_C02_rom_inst (.q(O26_I19_R0_C0_SM1 ),.address(input_fmap_19[7:0]),.clock  (clk));
logic [11-1:0] O26_I20_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O26_I20_R0_C02_rom_inst (.q(O26_I20_R0_C0_SM1 ),.address(input_fmap_20[7:0]),.clk(clk),.d(0),.we(0));
//assign O26_I20_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O26_I20_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O26_I20_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O26_I20_R0_C02_rom_inst (.q(O26_I20_R0_C0_SM1 ),.address(input_fmap_20[7:0]),.clock  (clk));
logic [10-1:0] O26_I22_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O26_I22_R0_C01_rom_inst (.q(O26_I22_R0_C0_SM1 ),.address(input_fmap_22[7:0]),.clk(clk),.d(0),.we(0));
//assign O26_I22_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O26_I22_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O26_I22_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O26_I22_R0_C01_rom_inst (.q(O26_I22_R0_C0_SM1 ),.address(input_fmap_22[7:0]),.clock  (clk));
logic [11-1:0] O26_I25_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O26_I25_R0_C02_rom_inst (.q(O26_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clk(clk),.d(0),.we(0));
//assign O26_I25_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O26_I25_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O26_I25_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O26_I25_R0_C02_rom_inst (.q(O26_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clock  (clk));
logic [10-1:0] O26_I26_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O26_I26_R0_C01_rom_inst (.q(O26_I26_R0_C0_SM1 ),.address(input_fmap_26[7:0]),.clk(clk),.d(0),.we(0));
//assign O26_I26_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O26_I26_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O26_I26_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O26_I26_R0_C01_rom_inst (.q(O26_I26_R0_C0_SM1 ),.address(input_fmap_26[7:0]),.clock  (clk));
logic [10-1:0] O26_I29_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O26_I29_R0_C01_rom_inst (.q(O26_I29_R0_C0_SM1 ),.address(input_fmap_29[7:0]),.clk(clk),.d(0),.we(0));
//assign O26_I29_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O26_I29_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O26_I29_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O26_I29_R0_C01_rom_inst (.q(O26_I29_R0_C0_SM1 ),.address(input_fmap_29[7:0]),.clock  (clk));
logic [10-1:0] O27_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O27_I0_R0_C01_rom_inst (.q(O27_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O27_I0_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O27_I0_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O27_I0_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O27_I0_R0_C01_rom_inst (.q(O27_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [10-1:0] O27_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O27_I3_R0_C01_rom_inst (.q(O27_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O27_I3_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O27_I3_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O27_I3_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O27_I3_R0_C01_rom_inst (.q(O27_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [10-1:0] O27_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O27_I4_R0_C01_rom_inst (.q(O27_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O27_I4_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O27_I4_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O27_I4_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O27_I4_R0_C01_rom_inst (.q(O27_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [10-1:0] O27_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O27_I5_R0_C01_rom_inst (.q(O27_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O27_I5_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O27_I5_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O27_I5_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O27_I5_R0_C01_rom_inst (.q(O27_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [10-1:0] O27_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O27_I8_R0_C01_rom_inst (.q(O27_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O27_I8_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O27_I8_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O27_I8_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O27_I8_R0_C01_rom_inst (.q(O27_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [11-1:0] O27_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O27_I9_R0_C02_rom_inst (.q(O27_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O27_I9_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O27_I9_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O27_I9_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O27_I9_R0_C02_rom_inst (.q(O27_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [10-1:0] O27_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O27_I12_R0_C01_rom_inst (.q(O27_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O27_I12_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O27_I12_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O27_I12_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O27_I12_R0_C01_rom_inst (.q(O27_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [10-1:0] O27_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O27_I13_R0_C01_rom_inst (.q(O27_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O27_I13_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O27_I13_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O27_I13_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O27_I13_R0_C01_rom_inst (.q(O27_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [10-1:0] O27_I18_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O27_I18_R0_C01_rom_inst (.q(O27_I18_R0_C0_SM1 ),.address(input_fmap_18[7:0]),.clk(clk),.d(0),.we(0));
//assign O27_I18_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O27_I18_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O27_I18_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O27_I18_R0_C01_rom_inst (.q(O27_I18_R0_C0_SM1 ),.address(input_fmap_18[7:0]),.clock  (clk));
logic [11-1:0] O27_I19_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O27_I19_R0_C02_rom_inst (.q(O27_I19_R0_C0_SM1 ),.address(input_fmap_19[7:0]),.clk(clk),.d(0),.we(0));
//assign O27_I19_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O27_I19_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O27_I19_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O27_I19_R0_C02_rom_inst (.q(O27_I19_R0_C0_SM1 ),.address(input_fmap_19[7:0]),.clock  (clk));
logic [10-1:0] O27_I21_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O27_I21_R0_C01_rom_inst (.q(O27_I21_R0_C0_SM1 ),.address(input_fmap_21[7:0]),.clk(clk),.d(0),.we(0));
//assign O27_I21_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O27_I21_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O27_I21_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O27_I21_R0_C01_rom_inst (.q(O27_I21_R0_C0_SM1 ),.address(input_fmap_21[7:0]),.clock  (clk));
logic [10-1:0] O27_I22_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O27_I22_R0_C01_rom_inst (.q(O27_I22_R0_C0_SM1 ),.address(input_fmap_22[7:0]),.clk(clk),.d(0),.we(0));
//assign O27_I22_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O27_I22_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O27_I22_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O27_I22_R0_C01_rom_inst (.q(O27_I22_R0_C0_SM1 ),.address(input_fmap_22[7:0]),.clock  (clk));
logic [11-1:0] O27_I23_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O27_I23_R0_C02_rom_inst (.q(O27_I23_R0_C0_SM1 ),.address(input_fmap_23[7:0]),.clk(clk),.d(0),.we(0));
//assign O27_I23_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O27_I23_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O27_I23_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O27_I23_R0_C02_rom_inst (.q(O27_I23_R0_C0_SM1 ),.address(input_fmap_23[7:0]),.clock  (clk));
logic [10-1:0] O27_I26_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O27_I26_R0_C01_rom_inst (.q(O27_I26_R0_C0_SM1 ),.address(input_fmap_26[7:0]),.clk(clk),.d(0),.we(0));
//assign O27_I26_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O27_I26_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O27_I26_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O27_I26_R0_C01_rom_inst (.q(O27_I26_R0_C0_SM1 ),.address(input_fmap_26[7:0]),.clock  (clk));
logic [10-1:0] O27_I29_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O27_I29_R0_C01_rom_inst (.q(O27_I29_R0_C0_SM1 ),.address(input_fmap_29[7:0]),.clk(clk),.d(0),.we(0));
//assign O27_I29_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O27_I29_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O27_I29_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O27_I29_R0_C01_rom_inst (.q(O27_I29_R0_C0_SM1 ),.address(input_fmap_29[7:0]),.clock  (clk));
logic [10-1:0] O27_I30_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O27_I30_R0_C01_rom_inst (.q(O27_I30_R0_C0_SM1 ),.address(input_fmap_30[7:0]),.clk(clk),.d(0),.we(0));
//assign O27_I30_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O27_I30_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O27_I30_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O27_I30_R0_C01_rom_inst (.q(O27_I30_R0_C0_SM1 ),.address(input_fmap_30[7:0]),.clock  (clk));
logic [11-1:0] O27_I31_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O27_I31_R0_C03_rom_inst (.q(O27_I31_R0_C0_SM1 ),.address(input_fmap_31[7:0]),.clk(clk),.d(0),.we(0));
//assign O27_I31_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O27_I31_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O27_I31_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O27_I31_R0_C03_rom_inst (.q(O27_I31_R0_C0_SM1 ),.address(input_fmap_31[7:0]),.clock  (clk));
logic [10-1:0] O28_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O28_I0_R0_C01_rom_inst (.q(O28_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O28_I0_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O28_I0_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O28_I0_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O28_I0_R0_C01_rom_inst (.q(O28_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [10-1:0] O28_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O28_I1_R0_C01_rom_inst (.q(O28_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O28_I1_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O28_I1_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O28_I1_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O28_I1_R0_C01_rom_inst (.q(O28_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [10-1:0] O28_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O28_I2_R0_C01_rom_inst (.q(O28_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O28_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O28_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O28_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O28_I2_R0_C01_rom_inst (.q(O28_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [10-1:0] O28_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O28_I6_R0_C01_rom_inst (.q(O28_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O28_I6_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O28_I6_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O28_I6_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O28_I6_R0_C01_rom_inst (.q(O28_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [10-1:0] O28_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O28_I7_R0_C01_rom_inst (.q(O28_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O28_I7_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O28_I7_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O28_I7_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O28_I7_R0_C01_rom_inst (.q(O28_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [10-1:0] O28_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O28_I8_R0_C01_rom_inst (.q(O28_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O28_I8_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O28_I8_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O28_I8_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O28_I8_R0_C01_rom_inst (.q(O28_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [11-1:0] O28_I9_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O28_I9_R0_C03_rom_inst (.q(O28_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clk(clk),.d(0),.we(0));
//assign O28_I9_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O28_I9_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O28_I9_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O28_I9_R0_C03_rom_inst (.q(O28_I9_R0_C0_SM1 ),.address(input_fmap_9[7:0]),.clock  (clk));
logic [11-1:0] O28_I14_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O28_I14_R0_C03_rom_inst (.q(O28_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clk(clk),.d(0),.we(0));
//assign O28_I14_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O28_I14_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O28_I14_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O28_I14_R0_C03_rom_inst (.q(O28_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clock  (clk));
logic [11-1:0] O28_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O28_I15_R0_C02_rom_inst (.q(O28_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O28_I15_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O28_I15_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O28_I15_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O28_I15_R0_C02_rom_inst (.q(O28_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [10-1:0] O28_I16_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O28_I16_R0_C01_rom_inst (.q(O28_I16_R0_C0_SM1 ),.address(input_fmap_16[7:0]),.clk(clk),.d(0),.we(0));
//assign O28_I16_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O28_I16_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O28_I16_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O28_I16_R0_C01_rom_inst (.q(O28_I16_R0_C0_SM1 ),.address(input_fmap_16[7:0]),.clock  (clk));
logic [10-1:0] O28_I18_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O28_I18_R0_C01_rom_inst (.q(O28_I18_R0_C0_SM1 ),.address(input_fmap_18[7:0]),.clk(clk),.d(0),.we(0));
//assign O28_I18_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O28_I18_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O28_I18_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O28_I18_R0_C01_rom_inst (.q(O28_I18_R0_C0_SM1 ),.address(input_fmap_18[7:0]),.clock  (clk));
logic [11-1:0] O28_I21_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O28_I21_R0_C02_rom_inst (.q(O28_I21_R0_C0_SM1 ),.address(input_fmap_21[7:0]),.clk(clk),.d(0),.we(0));
//assign O28_I21_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O28_I21_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O28_I21_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O28_I21_R0_C02_rom_inst (.q(O28_I21_R0_C0_SM1 ),.address(input_fmap_21[7:0]),.clock  (clk));
logic [10-1:0] O28_I22_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O28_I22_R0_C01_rom_inst (.q(O28_I22_R0_C0_SM1 ),.address(input_fmap_22[7:0]),.clk(clk),.d(0),.we(0));
//assign O28_I22_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O28_I22_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O28_I22_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O28_I22_R0_C01_rom_inst (.q(O28_I22_R0_C0_SM1 ),.address(input_fmap_22[7:0]),.clock  (clk));
logic [10-1:0] O28_I23_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O28_I23_R0_C01_rom_inst (.q(O28_I23_R0_C0_SM1 ),.address(input_fmap_23[7:0]),.clk(clk),.d(0),.we(0));
//assign O28_I23_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O28_I23_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O28_I23_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O28_I23_R0_C01_rom_inst (.q(O28_I23_R0_C0_SM1 ),.address(input_fmap_23[7:0]),.clock  (clk));
logic [10-1:0] O28_I24_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O28_I24_R0_C01_rom_inst (.q(O28_I24_R0_C0_SM1 ),.address(input_fmap_24[7:0]),.clk(clk),.d(0),.we(0));
//assign O28_I24_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O28_I24_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O28_I24_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O28_I24_R0_C01_rom_inst (.q(O28_I24_R0_C0_SM1 ),.address(input_fmap_24[7:0]),.clock  (clk));
logic [12-1:0] O28_I25_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(12),.INIT_FILE("deepfreeze_rom/deepfreeze_8_12.txt"))
    conv5_pw_O28_I25_R0_C04_rom_inst (.q(O28_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clk(clk),.d(0),.we(0));
//assign O28_I25_R0_C0_SM1  = 12'h1234;
//always@(posedge clk) begin 
//O28_I25_R0_C0_SM1  <= 12'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O28_I25_R0_C04_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(12))
//    conv5_pw_O28_I25_R0_C04_rom_inst (.q(O28_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clock  (clk));
logic [10-1:0] O28_I27_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O28_I27_R0_C01_rom_inst (.q(O28_I27_R0_C0_SM1 ),.address(input_fmap_27[7:0]),.clk(clk),.d(0),.we(0));
//assign O28_I27_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O28_I27_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O28_I27_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O28_I27_R0_C01_rom_inst (.q(O28_I27_R0_C0_SM1 ),.address(input_fmap_27[7:0]),.clock  (clk));
logic [10-1:0] O28_I28_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O28_I28_R0_C01_rom_inst (.q(O28_I28_R0_C0_SM1 ),.address(input_fmap_28[7:0]),.clk(clk),.d(0),.we(0));
//assign O28_I28_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O28_I28_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O28_I28_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O28_I28_R0_C01_rom_inst (.q(O28_I28_R0_C0_SM1 ),.address(input_fmap_28[7:0]),.clock  (clk));
logic [11-1:0] O28_I30_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O28_I30_R0_C02_rom_inst (.q(O28_I30_R0_C0_SM1 ),.address(input_fmap_30[7:0]),.clk(clk),.d(0),.we(0));
//assign O28_I30_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O28_I30_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O28_I30_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O28_I30_R0_C02_rom_inst (.q(O28_I30_R0_C0_SM1 ),.address(input_fmap_30[7:0]),.clock  (clk));
logic [11-1:0] O29_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O29_I0_R0_C02_rom_inst (.q(O29_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O29_I0_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O29_I0_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O29_I0_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O29_I0_R0_C02_rom_inst (.q(O29_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [10-1:0] O29_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O29_I1_R0_C01_rom_inst (.q(O29_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O29_I1_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O29_I1_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O29_I1_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O29_I1_R0_C01_rom_inst (.q(O29_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [10-1:0] O29_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O29_I2_R0_C01_rom_inst (.q(O29_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O29_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O29_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O29_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O29_I2_R0_C01_rom_inst (.q(O29_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [10-1:0] O29_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O29_I3_R0_C01_rom_inst (.q(O29_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O29_I3_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O29_I3_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O29_I3_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O29_I3_R0_C01_rom_inst (.q(O29_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [10-1:0] O29_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O29_I4_R0_C01_rom_inst (.q(O29_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O29_I4_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O29_I4_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O29_I4_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O29_I4_R0_C01_rom_inst (.q(O29_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [11-1:0] O29_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O29_I5_R0_C02_rom_inst (.q(O29_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O29_I5_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O29_I5_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O29_I5_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O29_I5_R0_C02_rom_inst (.q(O29_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [10-1:0] O29_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O29_I6_R0_C01_rom_inst (.q(O29_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O29_I6_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O29_I6_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O29_I6_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O29_I6_R0_C01_rom_inst (.q(O29_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [10-1:0] O29_I8_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O29_I8_R0_C01_rom_inst (.q(O29_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clk(clk),.d(0),.we(0));
//assign O29_I8_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O29_I8_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O29_I8_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O29_I8_R0_C01_rom_inst (.q(O29_I8_R0_C0_SM1 ),.address(input_fmap_8[7:0]),.clock  (clk));
logic [10-1:0] O29_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O29_I11_R0_C01_rom_inst (.q(O29_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O29_I11_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O29_I11_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O29_I11_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O29_I11_R0_C01_rom_inst (.q(O29_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [11-1:0] O29_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O29_I12_R0_C03_rom_inst (.q(O29_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O29_I12_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O29_I12_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O29_I12_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O29_I12_R0_C03_rom_inst (.q(O29_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [11-1:0] O29_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O29_I13_R0_C02_rom_inst (.q(O29_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O29_I13_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O29_I13_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O29_I13_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O29_I13_R0_C02_rom_inst (.q(O29_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [10-1:0] O29_I16_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O29_I16_R0_C01_rom_inst (.q(O29_I16_R0_C0_SM1 ),.address(input_fmap_16[7:0]),.clk(clk),.d(0),.we(0));
//assign O29_I16_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O29_I16_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O29_I16_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O29_I16_R0_C01_rom_inst (.q(O29_I16_R0_C0_SM1 ),.address(input_fmap_16[7:0]),.clock  (clk));
logic [11-1:0] O29_I17_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O29_I17_R0_C02_rom_inst (.q(O29_I17_R0_C0_SM1 ),.address(input_fmap_17[7:0]),.clk(clk),.d(0),.we(0));
//assign O29_I17_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O29_I17_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O29_I17_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O29_I17_R0_C02_rom_inst (.q(O29_I17_R0_C0_SM1 ),.address(input_fmap_17[7:0]),.clock  (clk));
logic [10-1:0] O29_I19_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O29_I19_R0_C01_rom_inst (.q(O29_I19_R0_C0_SM1 ),.address(input_fmap_19[7:0]),.clk(clk),.d(0),.we(0));
//assign O29_I19_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O29_I19_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O29_I19_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O29_I19_R0_C01_rom_inst (.q(O29_I19_R0_C0_SM1 ),.address(input_fmap_19[7:0]),.clock  (clk));
logic [10-1:0] O29_I20_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O29_I20_R0_C01_rom_inst (.q(O29_I20_R0_C0_SM1 ),.address(input_fmap_20[7:0]),.clk(clk),.d(0),.we(0));
//assign O29_I20_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O29_I20_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O29_I20_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O29_I20_R0_C01_rom_inst (.q(O29_I20_R0_C0_SM1 ),.address(input_fmap_20[7:0]),.clock  (clk));
logic [10-1:0] O29_I21_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O29_I21_R0_C01_rom_inst (.q(O29_I21_R0_C0_SM1 ),.address(input_fmap_21[7:0]),.clk(clk),.d(0),.we(0));
//assign O29_I21_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O29_I21_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O29_I21_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O29_I21_R0_C01_rom_inst (.q(O29_I21_R0_C0_SM1 ),.address(input_fmap_21[7:0]),.clock  (clk));
logic [11-1:0] O29_I24_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O29_I24_R0_C02_rom_inst (.q(O29_I24_R0_C0_SM1 ),.address(input_fmap_24[7:0]),.clk(clk),.d(0),.we(0));
//assign O29_I24_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O29_I24_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O29_I24_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O29_I24_R0_C02_rom_inst (.q(O29_I24_R0_C0_SM1 ),.address(input_fmap_24[7:0]),.clock  (clk));
logic [10-1:0] O29_I26_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O29_I26_R0_C01_rom_inst (.q(O29_I26_R0_C0_SM1 ),.address(input_fmap_26[7:0]),.clk(clk),.d(0),.we(0));
//assign O29_I26_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O29_I26_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O29_I26_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O29_I26_R0_C01_rom_inst (.q(O29_I26_R0_C0_SM1 ),.address(input_fmap_26[7:0]),.clock  (clk));
logic [10-1:0] O29_I27_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O29_I27_R0_C01_rom_inst (.q(O29_I27_R0_C0_SM1 ),.address(input_fmap_27[7:0]),.clk(clk),.d(0),.we(0));
//assign O29_I27_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O29_I27_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O29_I27_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O29_I27_R0_C01_rom_inst (.q(O29_I27_R0_C0_SM1 ),.address(input_fmap_27[7:0]),.clock  (clk));
logic [10-1:0] O29_I29_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O29_I29_R0_C01_rom_inst (.q(O29_I29_R0_C0_SM1 ),.address(input_fmap_29[7:0]),.clk(clk),.d(0),.we(0));
//assign O29_I29_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O29_I29_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O29_I29_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O29_I29_R0_C01_rom_inst (.q(O29_I29_R0_C0_SM1 ),.address(input_fmap_29[7:0]),.clock  (clk));
logic [10-1:0] O29_I30_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O29_I30_R0_C01_rom_inst (.q(O29_I30_R0_C0_SM1 ),.address(input_fmap_30[7:0]),.clk(clk),.d(0),.we(0));
//assign O29_I30_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O29_I30_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O29_I30_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O29_I30_R0_C01_rom_inst (.q(O29_I30_R0_C0_SM1 ),.address(input_fmap_30[7:0]),.clock  (clk));
logic [10-1:0] O29_I31_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O29_I31_R0_C01_rom_inst (.q(O29_I31_R0_C0_SM1 ),.address(input_fmap_31[7:0]),.clk(clk),.d(0),.we(0));
//assign O29_I31_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O29_I31_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O29_I31_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O29_I31_R0_C01_rom_inst (.q(O29_I31_R0_C0_SM1 ),.address(input_fmap_31[7:0]),.clock  (clk));
logic [11-1:0] O30_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O30_I0_R0_C02_rom_inst (.q(O30_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O30_I0_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O30_I0_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O30_I0_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O30_I0_R0_C02_rom_inst (.q(O30_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [10-1:0] O30_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O30_I1_R0_C01_rom_inst (.q(O30_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O30_I1_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O30_I1_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O30_I1_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O30_I1_R0_C01_rom_inst (.q(O30_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [10-1:0] O30_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O30_I2_R0_C01_rom_inst (.q(O30_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O30_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O30_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O30_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O30_I2_R0_C01_rom_inst (.q(O30_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [10-1:0] O30_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O30_I3_R0_C01_rom_inst (.q(O30_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O30_I3_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O30_I3_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O30_I3_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O30_I3_R0_C01_rom_inst (.q(O30_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [10-1:0] O30_I5_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O30_I5_R0_C01_rom_inst (.q(O30_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clk(clk),.d(0),.we(0));
//assign O30_I5_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O30_I5_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O30_I5_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O30_I5_R0_C01_rom_inst (.q(O30_I5_R0_C0_SM1 ),.address(input_fmap_5[7:0]),.clock  (clk));
logic [10-1:0] O30_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O30_I6_R0_C01_rom_inst (.q(O30_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O30_I6_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O30_I6_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O30_I6_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O30_I6_R0_C01_rom_inst (.q(O30_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [10-1:0] O30_I10_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O30_I10_R0_C01_rom_inst (.q(O30_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clk(clk),.d(0),.we(0));
//assign O30_I10_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O30_I10_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O30_I10_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O30_I10_R0_C01_rom_inst (.q(O30_I10_R0_C0_SM1 ),.address(input_fmap_10[7:0]),.clock  (clk));
logic [10-1:0] O30_I11_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O30_I11_R0_C01_rom_inst (.q(O30_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clk(clk),.d(0),.we(0));
//assign O30_I11_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O30_I11_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O30_I11_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O30_I11_R0_C01_rom_inst (.q(O30_I11_R0_C0_SM1 ),.address(input_fmap_11[7:0]),.clock  (clk));
logic [10-1:0] O30_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O30_I13_R0_C01_rom_inst (.q(O30_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O30_I13_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O30_I13_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O30_I13_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O30_I13_R0_C01_rom_inst (.q(O30_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [11-1:0] O30_I14_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O30_I14_R0_C02_rom_inst (.q(O30_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clk(clk),.d(0),.we(0));
//assign O30_I14_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O30_I14_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O30_I14_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O30_I14_R0_C02_rom_inst (.q(O30_I14_R0_C0_SM1 ),.address(input_fmap_14[7:0]),.clock  (clk));
logic [10-1:0] O30_I15_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O30_I15_R0_C01_rom_inst (.q(O30_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clk(clk),.d(0),.we(0));
//assign O30_I15_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O30_I15_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O30_I15_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O30_I15_R0_C01_rom_inst (.q(O30_I15_R0_C0_SM1 ),.address(input_fmap_15[7:0]),.clock  (clk));
logic [10-1:0] O30_I16_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O30_I16_R0_C01_rom_inst (.q(O30_I16_R0_C0_SM1 ),.address(input_fmap_16[7:0]),.clk(clk),.d(0),.we(0));
//assign O30_I16_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O30_I16_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O30_I16_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O30_I16_R0_C01_rom_inst (.q(O30_I16_R0_C0_SM1 ),.address(input_fmap_16[7:0]),.clock  (clk));
logic [11-1:0] O30_I17_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O30_I17_R0_C03_rom_inst (.q(O30_I17_R0_C0_SM1 ),.address(input_fmap_17[7:0]),.clk(clk),.d(0),.we(0));
//assign O30_I17_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O30_I17_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O30_I17_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O30_I17_R0_C03_rom_inst (.q(O30_I17_R0_C0_SM1 ),.address(input_fmap_17[7:0]),.clock  (clk));
logic [10-1:0] O30_I18_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O30_I18_R0_C01_rom_inst (.q(O30_I18_R0_C0_SM1 ),.address(input_fmap_18[7:0]),.clk(clk),.d(0),.we(0));
//assign O30_I18_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O30_I18_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O30_I18_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O30_I18_R0_C01_rom_inst (.q(O30_I18_R0_C0_SM1 ),.address(input_fmap_18[7:0]),.clock  (clk));
logic [10-1:0] O30_I21_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O30_I21_R0_C01_rom_inst (.q(O30_I21_R0_C0_SM1 ),.address(input_fmap_21[7:0]),.clk(clk),.d(0),.we(0));
//assign O30_I21_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O30_I21_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O30_I21_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O30_I21_R0_C01_rom_inst (.q(O30_I21_R0_C0_SM1 ),.address(input_fmap_21[7:0]),.clock  (clk));
logic [11-1:0] O30_I22_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O30_I22_R0_C02_rom_inst (.q(O30_I22_R0_C0_SM1 ),.address(input_fmap_22[7:0]),.clk(clk),.d(0),.we(0));
//assign O30_I22_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O30_I22_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O30_I22_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O30_I22_R0_C02_rom_inst (.q(O30_I22_R0_C0_SM1 ),.address(input_fmap_22[7:0]),.clock  (clk));
logic [10-1:0] O30_I24_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O30_I24_R0_C01_rom_inst (.q(O30_I24_R0_C0_SM1 ),.address(input_fmap_24[7:0]),.clk(clk),.d(0),.we(0));
//assign O30_I24_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O30_I24_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O30_I24_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O30_I24_R0_C01_rom_inst (.q(O30_I24_R0_C0_SM1 ),.address(input_fmap_24[7:0]),.clock  (clk));
logic [10-1:0] O30_I25_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O30_I25_R0_C01_rom_inst (.q(O30_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clk(clk),.d(0),.we(0));
//assign O30_I25_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O30_I25_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O30_I25_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O30_I25_R0_C01_rom_inst (.q(O30_I25_R0_C0_SM1 ),.address(input_fmap_25[7:0]),.clock  (clk));
logic [11-1:0] O30_I27_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O30_I27_R0_C03_rom_inst (.q(O30_I27_R0_C0_SM1 ),.address(input_fmap_27[7:0]),.clk(clk),.d(0),.we(0));
//assign O30_I27_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O30_I27_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O30_I27_R0_C03_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O30_I27_R0_C03_rom_inst (.q(O30_I27_R0_C0_SM1 ),.address(input_fmap_27[7:0]),.clock  (clk));
logic [10-1:0] O30_I29_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O30_I29_R0_C01_rom_inst (.q(O30_I29_R0_C0_SM1 ),.address(input_fmap_29[7:0]),.clk(clk),.d(0),.we(0));
//assign O30_I29_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O30_I29_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O30_I29_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O30_I29_R0_C01_rom_inst (.q(O30_I29_R0_C0_SM1 ),.address(input_fmap_29[7:0]),.clock  (clk));
logic [10-1:0] O30_I31_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O30_I31_R0_C01_rom_inst (.q(O30_I31_R0_C0_SM1 ),.address(input_fmap_31[7:0]),.clk(clk),.d(0),.we(0));
//assign O30_I31_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O30_I31_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O30_I31_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O30_I31_R0_C01_rom_inst (.q(O30_I31_R0_C0_SM1 ),.address(input_fmap_31[7:0]),.clock  (clk));
logic [10-1:0] O31_I0_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O31_I0_R0_C01_rom_inst (.q(O31_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clk(clk),.d(0),.we(0));
//assign O31_I0_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O31_I0_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O31_I0_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O31_I0_R0_C01_rom_inst (.q(O31_I0_R0_C0_SM1 ),.address(input_fmap_0[7:0]),.clock  (clk));
logic [10-1:0] O31_I1_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O31_I1_R0_C01_rom_inst (.q(O31_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clk(clk),.d(0),.we(0));
//assign O31_I1_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O31_I1_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O31_I1_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O31_I1_R0_C01_rom_inst (.q(O31_I1_R0_C0_SM1 ),.address(input_fmap_1[7:0]),.clock  (clk));
logic [10-1:0] O31_I2_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O31_I2_R0_C01_rom_inst (.q(O31_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clk(clk),.d(0),.we(0));
//assign O31_I2_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O31_I2_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O31_I2_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O31_I2_R0_C01_rom_inst (.q(O31_I2_R0_C0_SM1 ),.address(input_fmap_2[7:0]),.clock  (clk));
logic [10-1:0] O31_I3_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O31_I3_R0_C01_rom_inst (.q(O31_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clk(clk),.d(0),.we(0));
//assign O31_I3_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O31_I3_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O31_I3_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O31_I3_R0_C01_rom_inst (.q(O31_I3_R0_C0_SM1 ),.address(input_fmap_3[7:0]),.clock  (clk));
logic [10-1:0] O31_I4_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O31_I4_R0_C01_rom_inst (.q(O31_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clk(clk),.d(0),.we(0));
//assign O31_I4_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O31_I4_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O31_I4_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O31_I4_R0_C01_rom_inst (.q(O31_I4_R0_C0_SM1 ),.address(input_fmap_4[7:0]),.clock  (clk));
logic [10-1:0] O31_I6_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O31_I6_R0_C01_rom_inst (.q(O31_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clk(clk),.d(0),.we(0));
//assign O31_I6_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O31_I6_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O31_I6_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O31_I6_R0_C01_rom_inst (.q(O31_I6_R0_C0_SM1 ),.address(input_fmap_6[7:0]),.clock  (clk));
logic [10-1:0] O31_I7_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O31_I7_R0_C01_rom_inst (.q(O31_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clk(clk),.d(0),.we(0));
//assign O31_I7_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O31_I7_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O31_I7_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O31_I7_R0_C01_rom_inst (.q(O31_I7_R0_C0_SM1 ),.address(input_fmap_7[7:0]),.clock  (clk));
logic [10-1:0] O31_I12_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O31_I12_R0_C01_rom_inst (.q(O31_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clk(clk),.d(0),.we(0));
//assign O31_I12_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O31_I12_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O31_I12_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O31_I12_R0_C01_rom_inst (.q(O31_I12_R0_C0_SM1 ),.address(input_fmap_12[7:0]),.clock  (clk));
logic [11-1:0] O31_I13_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(11),.INIT_FILE("deepfreeze_rom/deepfreeze_8_11.txt"))
    conv5_pw_O31_I13_R0_C02_rom_inst (.q(O31_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clk(clk),.d(0),.we(0));
//assign O31_I13_R0_C0_SM1  = 11'h1234;
//always@(posedge clk) begin 
//O31_I13_R0_C0_SM1  <= 11'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O31_I13_R0_C02_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(11))
//    conv5_pw_O31_I13_R0_C02_rom_inst (.q(O31_I13_R0_C0_SM1 ),.address(input_fmap_13[7:0]),.clock  (clk));
logic [10-1:0] O31_I16_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O31_I16_R0_C01_rom_inst (.q(O31_I16_R0_C0_SM1 ),.address(input_fmap_16[7:0]),.clk(clk),.d(0),.we(0));
//assign O31_I16_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O31_I16_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O31_I16_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O31_I16_R0_C01_rom_inst (.q(O31_I16_R0_C0_SM1 ),.address(input_fmap_16[7:0]),.clock  (clk));
logic [10-1:0] O31_I17_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O31_I17_R0_C01_rom_inst (.q(O31_I17_R0_C0_SM1 ),.address(input_fmap_17[7:0]),.clk(clk),.d(0),.we(0));
//assign O31_I17_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O31_I17_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O31_I17_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O31_I17_R0_C01_rom_inst (.q(O31_I17_R0_C0_SM1 ),.address(input_fmap_17[7:0]),.clock  (clk));
logic [10-1:0] O31_I19_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O31_I19_R0_C01_rom_inst (.q(O31_I19_R0_C0_SM1 ),.address(input_fmap_19[7:0]),.clk(clk),.d(0),.we(0));
//assign O31_I19_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O31_I19_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O31_I19_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O31_I19_R0_C01_rom_inst (.q(O31_I19_R0_C0_SM1 ),.address(input_fmap_19[7:0]),.clock  (clk));
logic [10-1:0] O31_I28_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O31_I28_R0_C01_rom_inst (.q(O31_I28_R0_C0_SM1 ),.address(input_fmap_28[7:0]),.clk(clk),.d(0),.we(0));
//assign O31_I28_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O31_I28_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O31_I28_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O31_I28_R0_C01_rom_inst (.q(O31_I28_R0_C0_SM1 ),.address(input_fmap_28[7:0]),.clock  (clk));
logic [10-1:0] O31_I30_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O31_I30_R0_C01_rom_inst (.q(O31_I30_R0_C0_SM1 ),.address(input_fmap_30[7:0]),.clk(clk),.d(0),.we(0));
//assign O31_I30_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O31_I30_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O31_I30_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O31_I30_R0_C01_rom_inst (.q(O31_I30_R0_C0_SM1 ),.address(input_fmap_30[7:0]),.clock  (clk));
logic [10-1:0] O31_I31_R0_C0_SM1 ;
ram_single # (.WORDS(256),.A_WIDTH(8),.D_WIDTH(10),.INIT_FILE("deepfreeze_rom/deepfreeze_8_10.txt"))
    conv5_pw_O31_I31_R0_C01_rom_inst (.q(O31_I31_R0_C0_SM1 ),.address(input_fmap_31[7:0]),.clk(clk),.d(0),.we(0));
//assign O31_I31_R0_C0_SM1  = 10'h1234;
//always@(posedge clk) begin 
//O31_I31_R0_C0_SM1  <= 10'h1234; 
//end
// singleport_rom # (.INIT_FILE("/home/data1/karan/DeepFreeze/DeepFreeze/DeepFreeze/examples/mobilenet_trained/ROM_init_files/conv5_pw_O31_I31_R0_C01_rom.mif"),.WORDS(256),.A_WIDTH(8),.D_WIDTH(10))
//    conv5_pw_O31_I31_R0_C01_rom_inst (.q(O31_I31_R0_C0_SM1 ),.address(input_fmap_31[7:0]),.clock  (clk));
logic signed [31:0] conv_mac_0;
logic signed [31:0] O0_N0_S0;		always @(posedge clk) O0_N0_S0 <=     O0_I0_R0_C0_SM1   +  O0_I2_R0_C0_SM1  ;
 logic signed [31:0] O0_N2_S0;		always @(posedge clk) O0_N2_S0 <=     O0_I4_R0_C0_SM1   +  O0_I5_R0_C0_SM1  ;
 logic signed [31:0] O0_N4_S0;		always @(posedge clk) O0_N4_S0 <=     O0_I6_R0_C0_SM1   +  O0_I7_R0_C0_SM1  ;
 logic signed [31:0] O0_N6_S0;		always @(posedge clk) O0_N6_S0 <=     O0_I8_R0_C0_SM1   +  O0_I9_R0_C0_SM1  ;
 logic signed [31:0] O0_N8_S0;		always @(posedge clk) O0_N8_S0 <=     O0_I11_R0_C0_SM1   +  O0_I13_R0_C0_SM1  ;
 logic signed [31:0] O0_N10_S0;		always @(posedge clk) O0_N10_S0 <=     O0_I17_R0_C0_SM1   +  O0_I19_R0_C0_SM1  ;
 logic signed [31:0] O0_N12_S0;		always @(posedge clk) O0_N12_S0 <=     O0_I20_R0_C0_SM1   +  O0_I23_R0_C0_SM1  ;
 logic signed [31:0] O0_N14_S0;		always @(posedge clk) O0_N14_S0 <=     O0_I25_R0_C0_SM1   +  O0_I29_R0_C0_SM1  ;
 logic signed [31:0] O0_N16_S0;		always @(posedge clk) O0_N16_S0 <=     O0_I31_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O0_N0_S1;		always @(posedge clk) O0_N0_S1 <=     O0_N0_S0  +  O0_N2_S0 ;
 logic signed [31:0] O0_N2_S1;		always @(posedge clk) O0_N2_S1 <=     O0_N4_S0  +  O0_N6_S0 ;
 logic signed [31:0] O0_N4_S1;		always @(posedge clk) O0_N4_S1 <=     O0_N8_S0  +  O0_N10_S0 ;
 logic signed [31:0] O0_N6_S1;		always @(posedge clk) O0_N6_S1 <=     O0_N12_S0  +  O0_N14_S0 ;
 logic signed [31:0] O0_N8_S1;		always @(posedge clk) O0_N8_S1 <=     O0_N16_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O0_N0_S2;		always @(posedge clk) O0_N0_S2 <=     O0_N0_S1  +  O0_N2_S1 ;
 logic signed [31:0] O0_N2_S2;		always @(posedge clk) O0_N2_S2 <=     O0_N4_S1  +  O0_N6_S1 ;
 logic signed [31:0] O0_N4_S2;		always @(posedge clk) O0_N4_S2 <=     O0_N8_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O0_N0_S3;		always @(posedge clk) O0_N0_S3 <=     O0_N0_S2  +  O0_N2_S2 ;
 logic signed [31:0] O0_N2_S3;		always @(posedge clk) O0_N2_S3 <=     O0_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O0_N0_S4;		always @(posedge clk) O0_N0_S4 <=     O0_N0_S3  +  O0_N2_S3 ;
 assign conv_mac_0 = O0_N0_S4;

logic signed [31:0] conv_mac_1;
logic signed [31:0] O1_N0_S0;		always @(posedge clk) O1_N0_S0 <=     O1_I9_R0_C0_SM1   +  O1_I11_R0_C0_SM1  ;
 logic signed [31:0] O1_N2_S0;		always @(posedge clk) O1_N2_S0 <=     O1_I23_R0_C0_SM1   +  O1_I26_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O1_N0_S1;		always @(posedge clk) O1_N0_S1 <=     O1_N0_S0  +  O1_N2_S0 ;
 assign conv_mac_1 = O1_N0_S1;

logic signed [31:0] conv_mac_2;
logic signed [31:0] O2_N0_S0;		always @(posedge clk) O2_N0_S0 <=     O2_I3_R0_C0_SM1   +  O2_I7_R0_C0_SM1  ;
 logic signed [31:0] O2_N2_S0;		always @(posedge clk) O2_N2_S0 <=     O2_I9_R0_C0_SM1   +  O2_I10_R0_C0_SM1  ;
 logic signed [31:0] O2_N4_S0;		always @(posedge clk) O2_N4_S0 <=     O2_I14_R0_C0_SM1   +  O2_I23_R0_C0_SM1  ;
 logic signed [31:0] O2_N6_S0;		always @(posedge clk) O2_N6_S0 <=     O2_I25_R0_C0_SM1   +  O2_I28_R0_C0_SM1  ;
 logic signed [31:0] O2_N8_S0;		always @(posedge clk) O2_N8_S0 <=     O2_I29_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O2_N0_S1;		always @(posedge clk) O2_N0_S1 <=     O2_N0_S0  +  O2_N2_S0 ;
 logic signed [31:0] O2_N2_S1;		always @(posedge clk) O2_N2_S1 <=     O2_N4_S0  +  O2_N6_S0 ;
 logic signed [31:0] O2_N4_S1;		always @(posedge clk) O2_N4_S1 <=     O2_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O2_N0_S2;		always @(posedge clk) O2_N0_S2 <=     O2_N0_S1  +  O2_N2_S1 ;
 logic signed [31:0] O2_N2_S2;		always @(posedge clk) O2_N2_S2 <=     O2_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O2_N0_S3;		always @(posedge clk) O2_N0_S3 <=     O2_N0_S2  +  O2_N2_S2 ;
 assign conv_mac_2 = O2_N0_S3;

logic signed [31:0] conv_mac_3;
logic signed [31:0] O3_N0_S0;		always @(posedge clk) O3_N0_S0 <=     O3_I1_R0_C0_SM1   +  O3_I2_R0_C0_SM1  ;
 logic signed [31:0] O3_N2_S0;		always @(posedge clk) O3_N2_S0 <=     O3_I3_R0_C0_SM1   +  O3_I5_R0_C0_SM1  ;
 logic signed [31:0] O3_N4_S0;		always @(posedge clk) O3_N4_S0 <=     O3_I6_R0_C0_SM1   +  O3_I7_R0_C0_SM1  ;
 logic signed [31:0] O3_N6_S0;		always @(posedge clk) O3_N6_S0 <=     O3_I8_R0_C0_SM1   +  O3_I9_R0_C0_SM1  ;
 logic signed [31:0] O3_N8_S0;		always @(posedge clk) O3_N8_S0 <=     O3_I10_R0_C0_SM1   +  O3_I12_R0_C0_SM1  ;
 logic signed [31:0] O3_N10_S0;		always @(posedge clk) O3_N10_S0 <=     O3_I13_R0_C0_SM1   +  O3_I14_R0_C0_SM1  ;
 logic signed [31:0] O3_N12_S0;		always @(posedge clk) O3_N12_S0 <=     O3_I15_R0_C0_SM1   +  O3_I16_R0_C0_SM1  ;
 logic signed [31:0] O3_N14_S0;		always @(posedge clk) O3_N14_S0 <=     O3_I18_R0_C0_SM1   +  O3_I21_R0_C0_SM1  ;
 logic signed [31:0] O3_N16_S0;		always @(posedge clk) O3_N16_S0 <=     O3_I22_R0_C0_SM1   +  O3_I23_R0_C0_SM1  ;
 logic signed [31:0] O3_N18_S0;		always @(posedge clk) O3_N18_S0 <=     O3_I24_R0_C0_SM1   +  O3_I25_R0_C0_SM1  ;
 logic signed [31:0] O3_N20_S0;		always @(posedge clk) O3_N20_S0 <=     O3_I29_R0_C0_SM1   +  O3_I30_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O3_N0_S1;		always @(posedge clk) O3_N0_S1 <=     O3_N0_S0  +  O3_N2_S0 ;
 logic signed [31:0] O3_N2_S1;		always @(posedge clk) O3_N2_S1 <=     O3_N4_S0  +  O3_N6_S0 ;
 logic signed [31:0] O3_N4_S1;		always @(posedge clk) O3_N4_S1 <=     O3_N8_S0  +  O3_N10_S0 ;
 logic signed [31:0] O3_N6_S1;		always @(posedge clk) O3_N6_S1 <=     O3_N12_S0  +  O3_N14_S0 ;
 logic signed [31:0] O3_N8_S1;		always @(posedge clk) O3_N8_S1 <=     O3_N16_S0  +  O3_N18_S0 ;
 logic signed [31:0] O3_N10_S1;		always @(posedge clk) O3_N10_S1 <=     O3_N20_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O3_N0_S2;		always @(posedge clk) O3_N0_S2 <=     O3_N0_S1  +  O3_N2_S1 ;
 logic signed [31:0] O3_N2_S2;		always @(posedge clk) O3_N2_S2 <=     O3_N4_S1  +  O3_N6_S1 ;
 logic signed [31:0] O3_N4_S2;		always @(posedge clk) O3_N4_S2 <=     O3_N8_S1  +  O3_N10_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O3_N0_S3;		always @(posedge clk) O3_N0_S3 <=     O3_N0_S2  +  O3_N2_S2 ;
 logic signed [31:0] O3_N2_S3;		always @(posedge clk) O3_N2_S3 <=     O3_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O3_N0_S4;		always @(posedge clk) O3_N0_S4 <=     O3_N0_S3  +  O3_N2_S3 ;
 assign conv_mac_3 = O3_N0_S4;

logic signed [31:0] conv_mac_4;
logic signed [31:0] O4_N0_S0;		always @(posedge clk) O4_N0_S0 <=     O4_I0_R0_C0_SM1   +  O4_I3_R0_C0_SM1  ;
 logic signed [31:0] O4_N2_S0;		always @(posedge clk) O4_N2_S0 <=     O4_I4_R0_C0_SM1   +  O4_I5_R0_C0_SM1  ;
 logic signed [31:0] O4_N4_S0;		always @(posedge clk) O4_N4_S0 <=     O4_I8_R0_C0_SM1   +  O4_I10_R0_C0_SM1  ;
 logic signed [31:0] O4_N6_S0;		always @(posedge clk) O4_N6_S0 <=     O4_I11_R0_C0_SM1   +  O4_I12_R0_C0_SM1  ;
 logic signed [31:0] O4_N8_S0;		always @(posedge clk) O4_N8_S0 <=     O4_I14_R0_C0_SM1   +  O4_I16_R0_C0_SM1  ;
 logic signed [31:0] O4_N10_S0;		always @(posedge clk) O4_N10_S0 <=     O4_I17_R0_C0_SM1   +  O4_I18_R0_C0_SM1  ;
 logic signed [31:0] O4_N12_S0;		always @(posedge clk) O4_N12_S0 <=     O4_I19_R0_C0_SM1   +  O4_I20_R0_C0_SM1  ;
 logic signed [31:0] O4_N14_S0;		always @(posedge clk) O4_N14_S0 <=     O4_I21_R0_C0_SM1   +  O4_I25_R0_C0_SM1  ;
 logic signed [31:0] O4_N16_S0;		always @(posedge clk) O4_N16_S0 <=     O4_I26_R0_C0_SM1   +  O4_I27_R0_C0_SM1  ;
 logic signed [31:0] O4_N18_S0;		always @(posedge clk) O4_N18_S0 <=     O4_I29_R0_C0_SM1   +  O4_I30_R0_C0_SM1  ;
 logic signed [31:0] O4_N20_S0;		always @(posedge clk) O4_N20_S0 <=     O4_I31_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O4_N0_S1;		always @(posedge clk) O4_N0_S1 <=     O4_N0_S0  +  O4_N2_S0 ;
 logic signed [31:0] O4_N2_S1;		always @(posedge clk) O4_N2_S1 <=     O4_N4_S0  +  O4_N6_S0 ;
 logic signed [31:0] O4_N4_S1;		always @(posedge clk) O4_N4_S1 <=     O4_N8_S0  +  O4_N10_S0 ;
 logic signed [31:0] O4_N6_S1;		always @(posedge clk) O4_N6_S1 <=     O4_N12_S0  +  O4_N14_S0 ;
 logic signed [31:0] O4_N8_S1;		always @(posedge clk) O4_N8_S1 <=     O4_N16_S0  +  O4_N18_S0 ;
 logic signed [31:0] O4_N10_S1;		always @(posedge clk) O4_N10_S1 <=     O4_N20_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O4_N0_S2;		always @(posedge clk) O4_N0_S2 <=     O4_N0_S1  +  O4_N2_S1 ;
 logic signed [31:0] O4_N2_S2;		always @(posedge clk) O4_N2_S2 <=     O4_N4_S1  +  O4_N6_S1 ;
 logic signed [31:0] O4_N4_S2;		always @(posedge clk) O4_N4_S2 <=     O4_N8_S1  +  O4_N10_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O4_N0_S3;		always @(posedge clk) O4_N0_S3 <=     O4_N0_S2  +  O4_N2_S2 ;
 logic signed [31:0] O4_N2_S3;		always @(posedge clk) O4_N2_S3 <=     O4_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O4_N0_S4;		always @(posedge clk) O4_N0_S4 <=     O4_N0_S3  +  O4_N2_S3 ;
 assign conv_mac_4 = O4_N0_S4;

logic signed [31:0] conv_mac_5;
logic signed [31:0] O5_N0_S0;		always @(posedge clk) O5_N0_S0 <=     O5_I0_R0_C0_SM1   +  O5_I1_R0_C0_SM1  ;
 logic signed [31:0] O5_N2_S0;		always @(posedge clk) O5_N2_S0 <=     O5_I2_R0_C0_SM1   +  O5_I5_R0_C0_SM1  ;
 logic signed [31:0] O5_N4_S0;		always @(posedge clk) O5_N4_S0 <=     O5_I9_R0_C0_SM1   +  O5_I12_R0_C0_SM1  ;
 logic signed [31:0] O5_N6_S0;		always @(posedge clk) O5_N6_S0 <=     O5_I19_R0_C0_SM1   +  O5_I20_R0_C0_SM1  ;
 logic signed [31:0] O5_N8_S0;		always @(posedge clk) O5_N8_S0 <=     O5_I23_R0_C0_SM1   +  O5_I24_R0_C0_SM1  ;
 logic signed [31:0] O5_N10_S0;		always @(posedge clk) O5_N10_S0 <=     O5_I25_R0_C0_SM1   +  O5_I28_R0_C0_SM1  ;
 logic signed [31:0] O5_N12_S0;		always @(posedge clk) O5_N12_S0 <=     O5_I30_R0_C0_SM1   +  O5_I31_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O5_N0_S1;		always @(posedge clk) O5_N0_S1 <=     O5_N0_S0  +  O5_N2_S0 ;
 logic signed [31:0] O5_N2_S1;		always @(posedge clk) O5_N2_S1 <=     O5_N4_S0  +  O5_N6_S0 ;
 logic signed [31:0] O5_N4_S1;		always @(posedge clk) O5_N4_S1 <=     O5_N8_S0  +  O5_N10_S0 ;
 logic signed [31:0] O5_N6_S1;		always @(posedge clk) O5_N6_S1 <=     O5_N12_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O5_N0_S2;		always @(posedge clk) O5_N0_S2 <=     O5_N0_S1  +  O5_N2_S1 ;
 logic signed [31:0] O5_N2_S2;		always @(posedge clk) O5_N2_S2 <=     O5_N4_S1  +  O5_N6_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O5_N0_S3;		always @(posedge clk) O5_N0_S3 <=     O5_N0_S2  +  O5_N2_S2 ;
 assign conv_mac_5 = O5_N0_S3;

logic signed [31:0] conv_mac_6;
logic signed [31:0] O6_N0_S0;		always @(posedge clk) O6_N0_S0 <=     O6_I0_R0_C0_SM1   +  O6_I1_R0_C0_SM1  ;
 logic signed [31:0] O6_N2_S0;		always @(posedge clk) O6_N2_S0 <=     O6_I2_R0_C0_SM1   +  O6_I4_R0_C0_SM1  ;
 logic signed [31:0] O6_N4_S0;		always @(posedge clk) O6_N4_S0 <=     O6_I6_R0_C0_SM1   +  O6_I7_R0_C0_SM1  ;
 logic signed [31:0] O6_N6_S0;		always @(posedge clk) O6_N6_S0 <=     O6_I8_R0_C0_SM1   +  O6_I10_R0_C0_SM1  ;
 logic signed [31:0] O6_N8_S0;		always @(posedge clk) O6_N8_S0 <=     O6_I14_R0_C0_SM1   +  O6_I15_R0_C0_SM1  ;
 logic signed [31:0] O6_N10_S0;		always @(posedge clk) O6_N10_S0 <=     O6_I16_R0_C0_SM1   +  O6_I17_R0_C0_SM1  ;
 logic signed [31:0] O6_N12_S0;		always @(posedge clk) O6_N12_S0 <=     O6_I19_R0_C0_SM1   +  O6_I20_R0_C0_SM1  ;
 logic signed [31:0] O6_N14_S0;		always @(posedge clk) O6_N14_S0 <=     O6_I21_R0_C0_SM1   +  O6_I22_R0_C0_SM1  ;
 logic signed [31:0] O6_N16_S0;		always @(posedge clk) O6_N16_S0 <=     O6_I23_R0_C0_SM1   +  O6_I24_R0_C0_SM1  ;
 logic signed [31:0] O6_N18_S0;		always @(posedge clk) O6_N18_S0 <=     O6_I25_R0_C0_SM1   +  O6_I26_R0_C0_SM1  ;
 logic signed [31:0] O6_N20_S0;		always @(posedge clk) O6_N20_S0 <=     O6_I27_R0_C0_SM1   +  O6_I28_R0_C0_SM1  ;
 logic signed [31:0] O6_N22_S0;		always @(posedge clk) O6_N22_S0 <=     O6_I29_R0_C0_SM1   +  O6_I31_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O6_N0_S1;		always @(posedge clk) O6_N0_S1 <=     O6_N0_S0  +  O6_N2_S0 ;
 logic signed [31:0] O6_N2_S1;		always @(posedge clk) O6_N2_S1 <=     O6_N4_S0  +  O6_N6_S0 ;
 logic signed [31:0] O6_N4_S1;		always @(posedge clk) O6_N4_S1 <=     O6_N8_S0  +  O6_N10_S0 ;
 logic signed [31:0] O6_N6_S1;		always @(posedge clk) O6_N6_S1 <=     O6_N12_S0  +  O6_N14_S0 ;
 logic signed [31:0] O6_N8_S1;		always @(posedge clk) O6_N8_S1 <=     O6_N16_S0  +  O6_N18_S0 ;
 logic signed [31:0] O6_N10_S1;		always @(posedge clk) O6_N10_S1 <=     O6_N20_S0  +  O6_N22_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O6_N0_S2;		always @(posedge clk) O6_N0_S2 <=     O6_N0_S1  +  O6_N2_S1 ;
 logic signed [31:0] O6_N2_S2;		always @(posedge clk) O6_N2_S2 <=     O6_N4_S1  +  O6_N6_S1 ;
 logic signed [31:0] O6_N4_S2;		always @(posedge clk) O6_N4_S2 <=     O6_N8_S1  +  O6_N10_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O6_N0_S3;		always @(posedge clk) O6_N0_S3 <=     O6_N0_S2  +  O6_N2_S2 ;
 logic signed [31:0] O6_N2_S3;		always @(posedge clk) O6_N2_S3 <=     O6_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O6_N0_S4;		always @(posedge clk) O6_N0_S4 <=     O6_N0_S3  +  O6_N2_S3 ;
 assign conv_mac_6 = O6_N0_S4;

logic signed [31:0] conv_mac_7;
logic signed [31:0] O7_N0_S0;		always @(posedge clk) O7_N0_S0 <=     O7_I3_R0_C0_SM1   +  O7_I9_R0_C0_SM1  ;
 logic signed [31:0] O7_N2_S0;		always @(posedge clk) O7_N2_S0 <=     O7_I14_R0_C0_SM1   +  O7_I15_R0_C0_SM1  ;
 logic signed [31:0] O7_N4_S0;		always @(posedge clk) O7_N4_S0 <=     O7_I18_R0_C0_SM1   +  O7_I23_R0_C0_SM1  ;
 logic signed [31:0] O7_N6_S0;		always @(posedge clk) O7_N6_S0 <=     O7_I27_R0_C0_SM1   +  O7_I28_R0_C0_SM1  ;
 logic signed [31:0] O7_N8_S0;		always @(posedge clk) O7_N8_S0 <=     O7_I29_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O7_N0_S1;		always @(posedge clk) O7_N0_S1 <=     O7_N0_S0  +  O7_N2_S0 ;
 logic signed [31:0] O7_N2_S1;		always @(posedge clk) O7_N2_S1 <=     O7_N4_S0  +  O7_N6_S0 ;
 logic signed [31:0] O7_N4_S1;		always @(posedge clk) O7_N4_S1 <=     O7_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O7_N0_S2;		always @(posedge clk) O7_N0_S2 <=     O7_N0_S1  +  O7_N2_S1 ;
 logic signed [31:0] O7_N2_S2;		always @(posedge clk) O7_N2_S2 <=     O7_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O7_N0_S3;		always @(posedge clk) O7_N0_S3 <=     O7_N0_S2  +  O7_N2_S2 ;
 assign conv_mac_7 = O7_N0_S3;

logic signed [31:0] conv_mac_8;
logic signed [31:0] O8_N0_S0;		always @(posedge clk) O8_N0_S0 <=     O8_I2_R0_C0_SM1   +  O8_I4_R0_C0_SM1  ;
 logic signed [31:0] O8_N2_S0;		always @(posedge clk) O8_N2_S0 <=     O8_I5_R0_C0_SM1   +  O8_I6_R0_C0_SM1  ;
 logic signed [31:0] O8_N4_S0;		always @(posedge clk) O8_N4_S0 <=     O8_I7_R0_C0_SM1   +  O8_I9_R0_C0_SM1  ;
 logic signed [31:0] O8_N6_S0;		always @(posedge clk) O8_N6_S0 <=     O8_I10_R0_C0_SM1   +  O8_I13_R0_C0_SM1  ;
 logic signed [31:0] O8_N8_S0;		always @(posedge clk) O8_N8_S0 <=     O8_I14_R0_C0_SM1   +  O8_I15_R0_C0_SM1  ;
 logic signed [31:0] O8_N10_S0;		always @(posedge clk) O8_N10_S0 <=     O8_I16_R0_C0_SM1   +  O8_I17_R0_C0_SM1  ;
 logic signed [31:0] O8_N12_S0;		always @(posedge clk) O8_N12_S0 <=     O8_I18_R0_C0_SM1   +  O8_I20_R0_C0_SM1  ;
 logic signed [31:0] O8_N14_S0;		always @(posedge clk) O8_N14_S0 <=     O8_I21_R0_C0_SM1   +  O8_I24_R0_C0_SM1  ;
 logic signed [31:0] O8_N16_S0;		always @(posedge clk) O8_N16_S0 <=     O8_I25_R0_C0_SM1   +  O8_I26_R0_C0_SM1  ;
 logic signed [31:0] O8_N18_S0;		always @(posedge clk) O8_N18_S0 <=     O8_I27_R0_C0_SM1   +  O8_I29_R0_C0_SM1  ;
 logic signed [31:0] O8_N20_S0;		always @(posedge clk) O8_N20_S0 <=     O8_I31_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O8_N0_S1;		always @(posedge clk) O8_N0_S1 <=     O8_N0_S0  +  O8_N2_S0 ;
 logic signed [31:0] O8_N2_S1;		always @(posedge clk) O8_N2_S1 <=     O8_N4_S0  +  O8_N6_S0 ;
 logic signed [31:0] O8_N4_S1;		always @(posedge clk) O8_N4_S1 <=     O8_N8_S0  +  O8_N10_S0 ;
 logic signed [31:0] O8_N6_S1;		always @(posedge clk) O8_N6_S1 <=     O8_N12_S0  +  O8_N14_S0 ;
 logic signed [31:0] O8_N8_S1;		always @(posedge clk) O8_N8_S1 <=     O8_N16_S0  +  O8_N18_S0 ;
 logic signed [31:0] O8_N10_S1;		always @(posedge clk) O8_N10_S1 <=     O8_N20_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O8_N0_S2;		always @(posedge clk) O8_N0_S2 <=     O8_N0_S1  +  O8_N2_S1 ;
 logic signed [31:0] O8_N2_S2;		always @(posedge clk) O8_N2_S2 <=     O8_N4_S1  +  O8_N6_S1 ;
 logic signed [31:0] O8_N4_S2;		always @(posedge clk) O8_N4_S2 <=     O8_N8_S1  +  O8_N10_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O8_N0_S3;		always @(posedge clk) O8_N0_S3 <=     O8_N0_S2  +  O8_N2_S2 ;
 logic signed [31:0] O8_N2_S3;		always @(posedge clk) O8_N2_S3 <=     O8_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O8_N0_S4;		always @(posedge clk) O8_N0_S4 <=     O8_N0_S3  +  O8_N2_S3 ;
 assign conv_mac_8 = O8_N0_S4;

logic signed [31:0] conv_mac_9;
logic signed [31:0] O9_N0_S0;		always @(posedge clk) O9_N0_S0 <=     O9_I0_R0_C0_SM1   +  O9_I1_R0_C0_SM1  ;
 logic signed [31:0] O9_N2_S0;		always @(posedge clk) O9_N2_S0 <=     O9_I2_R0_C0_SM1   +  O9_I5_R0_C0_SM1  ;
 logic signed [31:0] O9_N4_S0;		always @(posedge clk) O9_N4_S0 <=     O9_I6_R0_C0_SM1   +  O9_I9_R0_C0_SM1  ;
 logic signed [31:0] O9_N6_S0;		always @(posedge clk) O9_N6_S0 <=     O9_I10_R0_C0_SM1   +  O9_I11_R0_C0_SM1  ;
 logic signed [31:0] O9_N8_S0;		always @(posedge clk) O9_N8_S0 <=     O9_I13_R0_C0_SM1   +  O9_I14_R0_C0_SM1  ;
 logic signed [31:0] O9_N10_S0;		always @(posedge clk) O9_N10_S0 <=     O9_I16_R0_C0_SM1   +  O9_I17_R0_C0_SM1  ;
 logic signed [31:0] O9_N12_S0;		always @(posedge clk) O9_N12_S0 <=     O9_I19_R0_C0_SM1   +  O9_I24_R0_C0_SM1  ;
 logic signed [31:0] O9_N14_S0;		always @(posedge clk) O9_N14_S0 <=     O9_I25_R0_C0_SM1   +  O9_I26_R0_C0_SM1  ;
 logic signed [31:0] O9_N16_S0;		always @(posedge clk) O9_N16_S0 <=     O9_I28_R0_C0_SM1   +  O9_I31_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O9_N0_S1;		always @(posedge clk) O9_N0_S1 <=     O9_N0_S0  +  O9_N2_S0 ;
 logic signed [31:0] O9_N2_S1;		always @(posedge clk) O9_N2_S1 <=     O9_N4_S0  +  O9_N6_S0 ;
 logic signed [31:0] O9_N4_S1;		always @(posedge clk) O9_N4_S1 <=     O9_N8_S0  +  O9_N10_S0 ;
 logic signed [31:0] O9_N6_S1;		always @(posedge clk) O9_N6_S1 <=     O9_N12_S0  +  O9_N14_S0 ;
 logic signed [31:0] O9_N8_S1;		always @(posedge clk) O9_N8_S1 <=     O9_N16_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O9_N0_S2;		always @(posedge clk) O9_N0_S2 <=     O9_N0_S1  +  O9_N2_S1 ;
 logic signed [31:0] O9_N2_S2;		always @(posedge clk) O9_N2_S2 <=     O9_N4_S1  +  O9_N6_S1 ;
 logic signed [31:0] O9_N4_S2;		always @(posedge clk) O9_N4_S2 <=     O9_N8_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O9_N0_S3;		always @(posedge clk) O9_N0_S3 <=     O9_N0_S2  +  O9_N2_S2 ;
 logic signed [31:0] O9_N2_S3;		always @(posedge clk) O9_N2_S3 <=     O9_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O9_N0_S4;		always @(posedge clk) O9_N0_S4 <=     O9_N0_S3  +  O9_N2_S3 ;
 assign conv_mac_9 = O9_N0_S4;

logic signed [31:0] conv_mac_10;
logic signed [31:0] O10_N0_S0;		always @(posedge clk) O10_N0_S0 <=     O10_I1_R0_C0_SM1   +  O10_I2_R0_C0_SM1  ;
 logic signed [31:0] O10_N2_S0;		always @(posedge clk) O10_N2_S0 <=     O10_I4_R0_C0_SM1   +  O10_I8_R0_C0_SM1  ;
 logic signed [31:0] O10_N4_S0;		always @(posedge clk) O10_N4_S0 <=     O10_I9_R0_C0_SM1   +  O10_I11_R0_C0_SM1  ;
 logic signed [31:0] O10_N6_S0;		always @(posedge clk) O10_N6_S0 <=     O10_I12_R0_C0_SM1   +  O10_I16_R0_C0_SM1  ;
 logic signed [31:0] O10_N8_S0;		always @(posedge clk) O10_N8_S0 <=     O10_I19_R0_C0_SM1   +  O10_I20_R0_C0_SM1  ;
 logic signed [31:0] O10_N10_S0;		always @(posedge clk) O10_N10_S0 <=     O10_I23_R0_C0_SM1   +  O10_I25_R0_C0_SM1  ;
 logic signed [31:0] O10_N12_S0;		always @(posedge clk) O10_N12_S0 <=     O10_I26_R0_C0_SM1   +  O10_I28_R0_C0_SM1  ;
 logic signed [31:0] O10_N14_S0;		always @(posedge clk) O10_N14_S0 <=     O10_I30_R0_C0_SM1   +  O10_I31_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O10_N0_S1;		always @(posedge clk) O10_N0_S1 <=     O10_N0_S0  +  O10_N2_S0 ;
 logic signed [31:0] O10_N2_S1;		always @(posedge clk) O10_N2_S1 <=     O10_N4_S0  +  O10_N6_S0 ;
 logic signed [31:0] O10_N4_S1;		always @(posedge clk) O10_N4_S1 <=     O10_N8_S0  +  O10_N10_S0 ;
 logic signed [31:0] O10_N6_S1;		always @(posedge clk) O10_N6_S1 <=     O10_N12_S0  +  O10_N14_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O10_N0_S2;		always @(posedge clk) O10_N0_S2 <=     O10_N0_S1  +  O10_N2_S1 ;
 logic signed [31:0] O10_N2_S2;		always @(posedge clk) O10_N2_S2 <=     O10_N4_S1  +  O10_N6_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O10_N0_S3;		always @(posedge clk) O10_N0_S3 <=     O10_N0_S2  +  O10_N2_S2 ;
 assign conv_mac_10 = O10_N0_S3;

logic signed [31:0] conv_mac_11;
logic signed [31:0] O11_N0_S0;		always @(posedge clk) O11_N0_S0 <=     O11_I0_R0_C0_SM1   +  O11_I1_R0_C0_SM1  ;
 logic signed [31:0] O11_N2_S0;		always @(posedge clk) O11_N2_S0 <=     O11_I5_R0_C0_SM1   +  O11_I7_R0_C0_SM1  ;
 logic signed [31:0] O11_N4_S0;		always @(posedge clk) O11_N4_S0 <=     O11_I8_R0_C0_SM1   +  O11_I10_R0_C0_SM1  ;
 logic signed [31:0] O11_N6_S0;		always @(posedge clk) O11_N6_S0 <=     O11_I11_R0_C0_SM1   +  O11_I12_R0_C0_SM1  ;
 logic signed [31:0] O11_N8_S0;		always @(posedge clk) O11_N8_S0 <=     O11_I13_R0_C0_SM1   +  O11_I16_R0_C0_SM1  ;
 logic signed [31:0] O11_N10_S0;		always @(posedge clk) O11_N10_S0 <=     O11_I19_R0_C0_SM1   +  O11_I20_R0_C0_SM1  ;
 logic signed [31:0] O11_N12_S0;		always @(posedge clk) O11_N12_S0 <=     O11_I22_R0_C0_SM1   +  O11_I24_R0_C0_SM1  ;
 logic signed [31:0] O11_N14_S0;		always @(posedge clk) O11_N14_S0 <=     O11_I25_R0_C0_SM1   +  O11_I26_R0_C0_SM1  ;
 logic signed [31:0] O11_N16_S0;		always @(posedge clk) O11_N16_S0 <=     O11_I27_R0_C0_SM1   +  O11_I30_R0_C0_SM1  ;
 logic signed [31:0] O11_N18_S0;		always @(posedge clk) O11_N18_S0 <=     O11_I31_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O11_N0_S1;		always @(posedge clk) O11_N0_S1 <=     O11_N0_S0  +  O11_N2_S0 ;
 logic signed [31:0] O11_N2_S1;		always @(posedge clk) O11_N2_S1 <=     O11_N4_S0  +  O11_N6_S0 ;
 logic signed [31:0] O11_N4_S1;		always @(posedge clk) O11_N4_S1 <=     O11_N8_S0  +  O11_N10_S0 ;
 logic signed [31:0] O11_N6_S1;		always @(posedge clk) O11_N6_S1 <=     O11_N12_S0  +  O11_N14_S0 ;
 logic signed [31:0] O11_N8_S1;		always @(posedge clk) O11_N8_S1 <=     O11_N16_S0  +  O11_N18_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O11_N0_S2;		always @(posedge clk) O11_N0_S2 <=     O11_N0_S1  +  O11_N2_S1 ;
 logic signed [31:0] O11_N2_S2;		always @(posedge clk) O11_N2_S2 <=     O11_N4_S1  +  O11_N6_S1 ;
 logic signed [31:0] O11_N4_S2;		always @(posedge clk) O11_N4_S2 <=     O11_N8_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O11_N0_S3;		always @(posedge clk) O11_N0_S3 <=     O11_N0_S2  +  O11_N2_S2 ;
 logic signed [31:0] O11_N2_S3;		always @(posedge clk) O11_N2_S3 <=     O11_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O11_N0_S4;		always @(posedge clk) O11_N0_S4 <=     O11_N0_S3  +  O11_N2_S3 ;
 assign conv_mac_11 = O11_N0_S4;

logic signed [31:0] conv_mac_12;
logic signed [31:0] O12_N0_S0;		always @(posedge clk) O12_N0_S0 <=     O12_I0_R0_C0_SM1   +  O12_I1_R0_C0_SM1  ;
 logic signed [31:0] O12_N2_S0;		always @(posedge clk) O12_N2_S0 <=     O12_I2_R0_C0_SM1   +  O12_I3_R0_C0_SM1  ;
 logic signed [31:0] O12_N4_S0;		always @(posedge clk) O12_N4_S0 <=     O12_I5_R0_C0_SM1   +  O12_I6_R0_C0_SM1  ;
 logic signed [31:0] O12_N6_S0;		always @(posedge clk) O12_N6_S0 <=     O12_I7_R0_C0_SM1   +  O12_I9_R0_C0_SM1  ;
 logic signed [31:0] O12_N8_S0;		always @(posedge clk) O12_N8_S0 <=     O12_I10_R0_C0_SM1   +  O12_I11_R0_C0_SM1  ;
 logic signed [31:0] O12_N10_S0;		always @(posedge clk) O12_N10_S0 <=     O12_I12_R0_C0_SM1   +  O12_I13_R0_C0_SM1  ;
 logic signed [31:0] O12_N12_S0;		always @(posedge clk) O12_N12_S0 <=     O12_I14_R0_C0_SM1   +  O12_I15_R0_C0_SM1  ;
 logic signed [31:0] O12_N14_S0;		always @(posedge clk) O12_N14_S0 <=     O12_I17_R0_C0_SM1   +  O12_I18_R0_C0_SM1  ;
 logic signed [31:0] O12_N16_S0;		always @(posedge clk) O12_N16_S0 <=     O12_I20_R0_C0_SM1   +  O12_I24_R0_C0_SM1  ;
 logic signed [31:0] O12_N18_S0;		always @(posedge clk) O12_N18_S0 <=     O12_I25_R0_C0_SM1   +  O12_I27_R0_C0_SM1  ;
 logic signed [31:0] O12_N20_S0;		always @(posedge clk) O12_N20_S0 <=     O12_I29_R0_C0_SM1   +  O12_I30_R0_C0_SM1  ;
 logic signed [31:0] O12_N22_S0;		always @(posedge clk) O12_N22_S0 <=     O12_I31_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O12_N0_S1;		always @(posedge clk) O12_N0_S1 <=     O12_N0_S0  +  O12_N2_S0 ;
 logic signed [31:0] O12_N2_S1;		always @(posedge clk) O12_N2_S1 <=     O12_N4_S0  +  O12_N6_S0 ;
 logic signed [31:0] O12_N4_S1;		always @(posedge clk) O12_N4_S1 <=     O12_N8_S0  +  O12_N10_S0 ;
 logic signed [31:0] O12_N6_S1;		always @(posedge clk) O12_N6_S1 <=     O12_N12_S0  +  O12_N14_S0 ;
 logic signed [31:0] O12_N8_S1;		always @(posedge clk) O12_N8_S1 <=     O12_N16_S0  +  O12_N18_S0 ;
 logic signed [31:0] O12_N10_S1;		always @(posedge clk) O12_N10_S1 <=     O12_N20_S0  +  O12_N22_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O12_N0_S2;		always @(posedge clk) O12_N0_S2 <=     O12_N0_S1  +  O12_N2_S1 ;
 logic signed [31:0] O12_N2_S2;		always @(posedge clk) O12_N2_S2 <=     O12_N4_S1  +  O12_N6_S1 ;
 logic signed [31:0] O12_N4_S2;		always @(posedge clk) O12_N4_S2 <=     O12_N8_S1  +  O12_N10_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O12_N0_S3;		always @(posedge clk) O12_N0_S3 <=     O12_N0_S2  +  O12_N2_S2 ;
 logic signed [31:0] O12_N2_S3;		always @(posedge clk) O12_N2_S3 <=     O12_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O12_N0_S4;		always @(posedge clk) O12_N0_S4 <=     O12_N0_S3  +  O12_N2_S3 ;
 assign conv_mac_12 = O12_N0_S4;

logic signed [31:0] conv_mac_13;
logic signed [31:0] O13_N0_S0;		always @(posedge clk) O13_N0_S0 <=     O13_I1_R0_C0_SM1   +  O13_I2_R0_C0_SM1  ;
 logic signed [31:0] O13_N2_S0;		always @(posedge clk) O13_N2_S0 <=     O13_I4_R0_C0_SM1   +  O13_I5_R0_C0_SM1  ;
 logic signed [31:0] O13_N4_S0;		always @(posedge clk) O13_N4_S0 <=     O13_I9_R0_C0_SM1   +  O13_I11_R0_C0_SM1  ;
 logic signed [31:0] O13_N6_S0;		always @(posedge clk) O13_N6_S0 <=     O13_I15_R0_C0_SM1   +  O13_I16_R0_C0_SM1  ;
 logic signed [31:0] O13_N8_S0;		always @(posedge clk) O13_N8_S0 <=     O13_I20_R0_C0_SM1   +  O13_I21_R0_C0_SM1  ;
 logic signed [31:0] O13_N10_S0;		always @(posedge clk) O13_N10_S0 <=     O13_I22_R0_C0_SM1   +  O13_I25_R0_C0_SM1  ;
 logic signed [31:0] O13_N12_S0;		always @(posedge clk) O13_N12_S0 <=     O13_I27_R0_C0_SM1   +  O13_I28_R0_C0_SM1  ;
 logic signed [31:0] O13_N14_S0;		always @(posedge clk) O13_N14_S0 <=     O13_I30_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O13_N0_S1;		always @(posedge clk) O13_N0_S1 <=     O13_N0_S0  +  O13_N2_S0 ;
 logic signed [31:0] O13_N2_S1;		always @(posedge clk) O13_N2_S1 <=     O13_N4_S0  +  O13_N6_S0 ;
 logic signed [31:0] O13_N4_S1;		always @(posedge clk) O13_N4_S1 <=     O13_N8_S0  +  O13_N10_S0 ;
 logic signed [31:0] O13_N6_S1;		always @(posedge clk) O13_N6_S1 <=     O13_N12_S0  +  O13_N14_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O13_N0_S2;		always @(posedge clk) O13_N0_S2 <=     O13_N0_S1  +  O13_N2_S1 ;
 logic signed [31:0] O13_N2_S2;		always @(posedge clk) O13_N2_S2 <=     O13_N4_S1  +  O13_N6_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O13_N0_S3;		always @(posedge clk) O13_N0_S3 <=     O13_N0_S2  +  O13_N2_S2 ;
 assign conv_mac_13 = O13_N0_S3;

logic signed [31:0] conv_mac_14;
logic signed [31:0] O14_N0_S0;		always @(posedge clk) O14_N0_S0 <=     O14_I2_R0_C0_SM1   +  O14_I3_R0_C0_SM1  ;
 logic signed [31:0] O14_N2_S0;		always @(posedge clk) O14_N2_S0 <=     O14_I5_R0_C0_SM1   +  O14_I6_R0_C0_SM1  ;
 logic signed [31:0] O14_N4_S0;		always @(posedge clk) O14_N4_S0 <=     O14_I9_R0_C0_SM1   +  O14_I11_R0_C0_SM1  ;
 logic signed [31:0] O14_N6_S0;		always @(posedge clk) O14_N6_S0 <=     O14_I13_R0_C0_SM1   +  O14_I16_R0_C0_SM1  ;
 logic signed [31:0] O14_N8_S0;		always @(posedge clk) O14_N8_S0 <=     O14_I17_R0_C0_SM1   +  O14_I18_R0_C0_SM1  ;
 logic signed [31:0] O14_N10_S0;		always @(posedge clk) O14_N10_S0 <=     O14_I19_R0_C0_SM1   +  O14_I20_R0_C0_SM1  ;
 logic signed [31:0] O14_N12_S0;		always @(posedge clk) O14_N12_S0 <=     O14_I24_R0_C0_SM1   +  O14_I25_R0_C0_SM1  ;
 logic signed [31:0] O14_N14_S0;		always @(posedge clk) O14_N14_S0 <=     O14_I26_R0_C0_SM1   +  O14_I27_R0_C0_SM1  ;
 logic signed [31:0] O14_N16_S0;		always @(posedge clk) O14_N16_S0 <=     O14_I28_R0_C0_SM1   +  O14_I29_R0_C0_SM1  ;
 logic signed [31:0] O14_N18_S0;		always @(posedge clk) O14_N18_S0 <=     O14_I30_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O14_N0_S1;		always @(posedge clk) O14_N0_S1 <=     O14_N0_S0  +  O14_N2_S0 ;
 logic signed [31:0] O14_N2_S1;		always @(posedge clk) O14_N2_S1 <=     O14_N4_S0  +  O14_N6_S0 ;
 logic signed [31:0] O14_N4_S1;		always @(posedge clk) O14_N4_S1 <=     O14_N8_S0  +  O14_N10_S0 ;
 logic signed [31:0] O14_N6_S1;		always @(posedge clk) O14_N6_S1 <=     O14_N12_S0  +  O14_N14_S0 ;
 logic signed [31:0] O14_N8_S1;		always @(posedge clk) O14_N8_S1 <=     O14_N16_S0  +  O14_N18_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O14_N0_S2;		always @(posedge clk) O14_N0_S2 <=     O14_N0_S1  +  O14_N2_S1 ;
 logic signed [31:0] O14_N2_S2;		always @(posedge clk) O14_N2_S2 <=     O14_N4_S1  +  O14_N6_S1 ;
 logic signed [31:0] O14_N4_S2;		always @(posedge clk) O14_N4_S2 <=     O14_N8_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O14_N0_S3;		always @(posedge clk) O14_N0_S3 <=     O14_N0_S2  +  O14_N2_S2 ;
 logic signed [31:0] O14_N2_S3;		always @(posedge clk) O14_N2_S3 <=     O14_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O14_N0_S4;		always @(posedge clk) O14_N0_S4 <=     O14_N0_S3  +  O14_N2_S3 ;
 assign conv_mac_14 = O14_N0_S4;

logic signed [31:0] conv_mac_15;
logic signed [31:0] O15_N0_S0;		always @(posedge clk) O15_N0_S0 <=     O15_I0_R0_C0_SM1   +  O15_I2_R0_C0_SM1  ;
 logic signed [31:0] O15_N2_S0;		always @(posedge clk) O15_N2_S0 <=     O15_I4_R0_C0_SM1   +  O15_I5_R0_C0_SM1  ;
 logic signed [31:0] O15_N4_S0;		always @(posedge clk) O15_N4_S0 <=     O15_I6_R0_C0_SM1   +  O15_I7_R0_C0_SM1  ;
 logic signed [31:0] O15_N6_S0;		always @(posedge clk) O15_N6_S0 <=     O15_I8_R0_C0_SM1   +  O15_I9_R0_C0_SM1  ;
 logic signed [31:0] O15_N8_S0;		always @(posedge clk) O15_N8_S0 <=     O15_I10_R0_C0_SM1   +  O15_I11_R0_C0_SM1  ;
 logic signed [31:0] O15_N10_S0;		always @(posedge clk) O15_N10_S0 <=     O15_I12_R0_C0_SM1   +  O15_I13_R0_C0_SM1  ;
 logic signed [31:0] O15_N12_S0;		always @(posedge clk) O15_N12_S0 <=     O15_I15_R0_C0_SM1   +  O15_I16_R0_C0_SM1  ;
 logic signed [31:0] O15_N14_S0;		always @(posedge clk) O15_N14_S0 <=     O15_I18_R0_C0_SM1   +  O15_I19_R0_C0_SM1  ;
 logic signed [31:0] O15_N16_S0;		always @(posedge clk) O15_N16_S0 <=     O15_I20_R0_C0_SM1   +  O15_I21_R0_C0_SM1  ;
 logic signed [31:0] O15_N18_S0;		always @(posedge clk) O15_N18_S0 <=     O15_I22_R0_C0_SM1   +  O15_I23_R0_C0_SM1  ;
 logic signed [31:0] O15_N20_S0;		always @(posedge clk) O15_N20_S0 <=     O15_I24_R0_C0_SM1   +  O15_I25_R0_C0_SM1  ;
 logic signed [31:0] O15_N22_S0;		always @(posedge clk) O15_N22_S0 <=     O15_I26_R0_C0_SM1   +  O15_I28_R0_C0_SM1  ;
 logic signed [31:0] O15_N24_S0;		always @(posedge clk) O15_N24_S0 <=     O15_I30_R0_C0_SM1   +  O15_I31_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O15_N0_S1;		always @(posedge clk) O15_N0_S1 <=     O15_N0_S0  +  O15_N2_S0 ;
 logic signed [31:0] O15_N2_S1;		always @(posedge clk) O15_N2_S1 <=     O15_N4_S0  +  O15_N6_S0 ;
 logic signed [31:0] O15_N4_S1;		always @(posedge clk) O15_N4_S1 <=     O15_N8_S0  +  O15_N10_S0 ;
 logic signed [31:0] O15_N6_S1;		always @(posedge clk) O15_N6_S1 <=     O15_N12_S0  +  O15_N14_S0 ;
 logic signed [31:0] O15_N8_S1;		always @(posedge clk) O15_N8_S1 <=     O15_N16_S0  +  O15_N18_S0 ;
 logic signed [31:0] O15_N10_S1;		always @(posedge clk) O15_N10_S1 <=     O15_N20_S0  +  O15_N22_S0 ;
 logic signed [31:0] O15_N12_S1;		always @(posedge clk) O15_N12_S1 <=     O15_N24_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O15_N0_S2;		always @(posedge clk) O15_N0_S2 <=     O15_N0_S1  +  O15_N2_S1 ;
 logic signed [31:0] O15_N2_S2;		always @(posedge clk) O15_N2_S2 <=     O15_N4_S1  +  O15_N6_S1 ;
 logic signed [31:0] O15_N4_S2;		always @(posedge clk) O15_N4_S2 <=     O15_N8_S1  +  O15_N10_S1 ;
 logic signed [31:0] O15_N6_S2;		always @(posedge clk) O15_N6_S2 <=     O15_N12_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O15_N0_S3;		always @(posedge clk) O15_N0_S3 <=     O15_N0_S2  +  O15_N2_S2 ;
 logic signed [31:0] O15_N2_S3;		always @(posedge clk) O15_N2_S3 <=     O15_N4_S2  +  O15_N6_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O15_N0_S4;		always @(posedge clk) O15_N0_S4 <=     O15_N0_S3  +  O15_N2_S3 ;
 assign conv_mac_15 = O15_N0_S4;

logic signed [31:0] conv_mac_16;
logic signed [31:0] O16_N0_S0;		always @(posedge clk) O16_N0_S0 <=     O16_I1_R0_C0_SM1   +  O16_I4_R0_C0_SM1  ;
 logic signed [31:0] O16_N2_S0;		always @(posedge clk) O16_N2_S0 <=     O16_I5_R0_C0_SM1   +  O16_I7_R0_C0_SM1  ;
 logic signed [31:0] O16_N4_S0;		always @(posedge clk) O16_N4_S0 <=     O16_I8_R0_C0_SM1   +  O16_I10_R0_C0_SM1  ;
 logic signed [31:0] O16_N6_S0;		always @(posedge clk) O16_N6_S0 <=     O16_I11_R0_C0_SM1   +  O16_I12_R0_C0_SM1  ;
 logic signed [31:0] O16_N8_S0;		always @(posedge clk) O16_N8_S0 <=     O16_I14_R0_C0_SM1   +  O16_I15_R0_C0_SM1  ;
 logic signed [31:0] O16_N10_S0;		always @(posedge clk) O16_N10_S0 <=     O16_I17_R0_C0_SM1   +  O16_I18_R0_C0_SM1  ;
 logic signed [31:0] O16_N12_S0;		always @(posedge clk) O16_N12_S0 <=     O16_I19_R0_C0_SM1   +  O16_I20_R0_C0_SM1  ;
 logic signed [31:0] O16_N14_S0;		always @(posedge clk) O16_N14_S0 <=     O16_I23_R0_C0_SM1   +  O16_I25_R0_C0_SM1  ;
 logic signed [31:0] O16_N16_S0;		always @(posedge clk) O16_N16_S0 <=     O16_I26_R0_C0_SM1   +  O16_I27_R0_C0_SM1  ;
 logic signed [31:0] O16_N18_S0;		always @(posedge clk) O16_N18_S0 <=     O16_I28_R0_C0_SM1   +  O16_I29_R0_C0_SM1  ;
 logic signed [31:0] O16_N20_S0;		always @(posedge clk) O16_N20_S0 <=     O16_I30_R0_C0_SM1   +  O16_I31_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O16_N0_S1;		always @(posedge clk) O16_N0_S1 <=     O16_N0_S0  +  O16_N2_S0 ;
 logic signed [31:0] O16_N2_S1;		always @(posedge clk) O16_N2_S1 <=     O16_N4_S0  +  O16_N6_S0 ;
 logic signed [31:0] O16_N4_S1;		always @(posedge clk) O16_N4_S1 <=     O16_N8_S0  +  O16_N10_S0 ;
 logic signed [31:0] O16_N6_S1;		always @(posedge clk) O16_N6_S1 <=     O16_N12_S0  +  O16_N14_S0 ;
 logic signed [31:0] O16_N8_S1;		always @(posedge clk) O16_N8_S1 <=     O16_N16_S0  +  O16_N18_S0 ;
 logic signed [31:0] O16_N10_S1;		always @(posedge clk) O16_N10_S1 <=     O16_N20_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O16_N0_S2;		always @(posedge clk) O16_N0_S2 <=     O16_N0_S1  +  O16_N2_S1 ;
 logic signed [31:0] O16_N2_S2;		always @(posedge clk) O16_N2_S2 <=     O16_N4_S1  +  O16_N6_S1 ;
 logic signed [31:0] O16_N4_S2;		always @(posedge clk) O16_N4_S2 <=     O16_N8_S1  +  O16_N10_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O16_N0_S3;		always @(posedge clk) O16_N0_S3 <=     O16_N0_S2  +  O16_N2_S2 ;
 logic signed [31:0] O16_N2_S3;		always @(posedge clk) O16_N2_S3 <=     O16_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O16_N0_S4;		always @(posedge clk) O16_N0_S4 <=     O16_N0_S3  +  O16_N2_S3 ;
 assign conv_mac_16 = O16_N0_S4;

logic signed [31:0] conv_mac_17;
logic signed [31:0] O17_N0_S0;		always @(posedge clk) O17_N0_S0 <=     O17_I0_R0_C0_SM1   +  O17_I2_R0_C0_SM1  ;
 logic signed [31:0] O17_N2_S0;		always @(posedge clk) O17_N2_S0 <=     O17_I5_R0_C0_SM1   +  O17_I7_R0_C0_SM1  ;
 logic signed [31:0] O17_N4_S0;		always @(posedge clk) O17_N4_S0 <=     O17_I9_R0_C0_SM1   +  O17_I11_R0_C0_SM1  ;
 logic signed [31:0] O17_N6_S0;		always @(posedge clk) O17_N6_S0 <=     O17_I12_R0_C0_SM1   +  O17_I13_R0_C0_SM1  ;
 logic signed [31:0] O17_N8_S0;		always @(posedge clk) O17_N8_S0 <=     O17_I14_R0_C0_SM1   +  O17_I16_R0_C0_SM1  ;
 logic signed [31:0] O17_N10_S0;		always @(posedge clk) O17_N10_S0 <=     O17_I17_R0_C0_SM1   +  O17_I19_R0_C0_SM1  ;
 logic signed [31:0] O17_N12_S0;		always @(posedge clk) O17_N12_S0 <=     O17_I20_R0_C0_SM1   +  O17_I21_R0_C0_SM1  ;
 logic signed [31:0] O17_N14_S0;		always @(posedge clk) O17_N14_S0 <=     O17_I24_R0_C0_SM1   +  O17_I25_R0_C0_SM1  ;
 logic signed [31:0] O17_N16_S0;		always @(posedge clk) O17_N16_S0 <=     O17_I26_R0_C0_SM1   +  O17_I27_R0_C0_SM1  ;
 logic signed [31:0] O17_N18_S0;		always @(posedge clk) O17_N18_S0 <=     O17_I28_R0_C0_SM1   +  O17_I29_R0_C0_SM1  ;
 logic signed [31:0] O17_N20_S0;		always @(posedge clk) O17_N20_S0 <=     O17_I31_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O17_N0_S1;		always @(posedge clk) O17_N0_S1 <=     O17_N0_S0  +  O17_N2_S0 ;
 logic signed [31:0] O17_N2_S1;		always @(posedge clk) O17_N2_S1 <=     O17_N4_S0  +  O17_N6_S0 ;
 logic signed [31:0] O17_N4_S1;		always @(posedge clk) O17_N4_S1 <=     O17_N8_S0  +  O17_N10_S0 ;
 logic signed [31:0] O17_N6_S1;		always @(posedge clk) O17_N6_S1 <=     O17_N12_S0  +  O17_N14_S0 ;
 logic signed [31:0] O17_N8_S1;		always @(posedge clk) O17_N8_S1 <=     O17_N16_S0  +  O17_N18_S0 ;
 logic signed [31:0] O17_N10_S1;		always @(posedge clk) O17_N10_S1 <=     O17_N20_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O17_N0_S2;		always @(posedge clk) O17_N0_S2 <=     O17_N0_S1  +  O17_N2_S1 ;
 logic signed [31:0] O17_N2_S2;		always @(posedge clk) O17_N2_S2 <=     O17_N4_S1  +  O17_N6_S1 ;
 logic signed [31:0] O17_N4_S2;		always @(posedge clk) O17_N4_S2 <=     O17_N8_S1  +  O17_N10_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O17_N0_S3;		always @(posedge clk) O17_N0_S3 <=     O17_N0_S2  +  O17_N2_S2 ;
 logic signed [31:0] O17_N2_S3;		always @(posedge clk) O17_N2_S3 <=     O17_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O17_N0_S4;		always @(posedge clk) O17_N0_S4 <=     O17_N0_S3  +  O17_N2_S3 ;
 assign conv_mac_17 = O17_N0_S4;

logic signed [31:0] conv_mac_18;
logic signed [31:0] O18_N0_S0;		always @(posedge clk) O18_N0_S0 <=     O18_I2_R0_C0_SM1   +  O18_I4_R0_C0_SM1  ;
 logic signed [31:0] O18_N2_S0;		always @(posedge clk) O18_N2_S0 <=     O18_I5_R0_C0_SM1   +  O18_I6_R0_C0_SM1  ;
 logic signed [31:0] O18_N4_S0;		always @(posedge clk) O18_N4_S0 <=     O18_I7_R0_C0_SM1   +  O18_I9_R0_C0_SM1  ;
 logic signed [31:0] O18_N6_S0;		always @(posedge clk) O18_N6_S0 <=     O18_I11_R0_C0_SM1   +  O18_I12_R0_C0_SM1  ;
 logic signed [31:0] O18_N8_S0;		always @(posedge clk) O18_N8_S0 <=     O18_I17_R0_C0_SM1   +  O18_I19_R0_C0_SM1  ;
 logic signed [31:0] O18_N10_S0;		always @(posedge clk) O18_N10_S0 <=     O18_I21_R0_C0_SM1   +  O18_I22_R0_C0_SM1  ;
 logic signed [31:0] O18_N12_S0;		always @(posedge clk) O18_N12_S0 <=     O18_I23_R0_C0_SM1   +  O18_I26_R0_C0_SM1  ;
 logic signed [31:0] O18_N14_S0;		always @(posedge clk) O18_N14_S0 <=     O18_I28_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O18_N0_S1;		always @(posedge clk) O18_N0_S1 <=     O18_N0_S0  +  O18_N2_S0 ;
 logic signed [31:0] O18_N2_S1;		always @(posedge clk) O18_N2_S1 <=     O18_N4_S0  +  O18_N6_S0 ;
 logic signed [31:0] O18_N4_S1;		always @(posedge clk) O18_N4_S1 <=     O18_N8_S0  +  O18_N10_S0 ;
 logic signed [31:0] O18_N6_S1;		always @(posedge clk) O18_N6_S1 <=     O18_N12_S0  +  O18_N14_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O18_N0_S2;		always @(posedge clk) O18_N0_S2 <=     O18_N0_S1  +  O18_N2_S1 ;
 logic signed [31:0] O18_N2_S2;		always @(posedge clk) O18_N2_S2 <=     O18_N4_S1  +  O18_N6_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O18_N0_S3;		always @(posedge clk) O18_N0_S3 <=     O18_N0_S2  +  O18_N2_S2 ;
 assign conv_mac_18 = O18_N0_S3;

logic signed [31:0] conv_mac_19;
logic signed [31:0] O19_N0_S0;		always @(posedge clk) O19_N0_S0 <=     O19_I4_R0_C0_SM1   +  O19_I7_R0_C0_SM1  ;
 logic signed [31:0] O19_N2_S0;		always @(posedge clk) O19_N2_S0 <=     O19_I9_R0_C0_SM1   +  O19_I11_R0_C0_SM1  ;
 logic signed [31:0] O19_N4_S0;		always @(posedge clk) O19_N4_S0 <=     O19_I12_R0_C0_SM1   +  O19_I20_R0_C0_SM1  ;
 logic signed [31:0] O19_N6_S0;		always @(posedge clk) O19_N6_S0 <=     O19_I23_R0_C0_SM1   +  O19_I24_R0_C0_SM1  ;
 logic signed [31:0] O19_N8_S0;		always @(posedge clk) O19_N8_S0 <=     O19_I26_R0_C0_SM1   +  O19_I31_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O19_N0_S1;		always @(posedge clk) O19_N0_S1 <=     O19_N0_S0  +  O19_N2_S0 ;
 logic signed [31:0] O19_N2_S1;		always @(posedge clk) O19_N2_S1 <=     O19_N4_S0  +  O19_N6_S0 ;
 logic signed [31:0] O19_N4_S1;		always @(posedge clk) O19_N4_S1 <=     O19_N8_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O19_N0_S2;		always @(posedge clk) O19_N0_S2 <=     O19_N0_S1  +  O19_N2_S1 ;
 logic signed [31:0] O19_N2_S2;		always @(posedge clk) O19_N2_S2 <=     O19_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O19_N0_S3;		always @(posedge clk) O19_N0_S3 <=     O19_N0_S2  +  O19_N2_S2 ;
 assign conv_mac_19 = O19_N0_S3;

logic signed [31:0] conv_mac_20;
logic signed [31:0] O20_N0_S0;		always @(posedge clk) O20_N0_S0 <=     O20_I3_R0_C0_SM1   +  O20_I6_R0_C0_SM1  ;
 logic signed [31:0] O20_N2_S0;		always @(posedge clk) O20_N2_S0 <=     O20_I7_R0_C0_SM1   +  O20_I8_R0_C0_SM1  ;
 logic signed [31:0] O20_N4_S0;		always @(posedge clk) O20_N4_S0 <=     O20_I9_R0_C0_SM1   +  O20_I13_R0_C0_SM1  ;
 logic signed [31:0] O20_N6_S0;		always @(posedge clk) O20_N6_S0 <=     O20_I15_R0_C0_SM1   +  O20_I17_R0_C0_SM1  ;
 logic signed [31:0] O20_N8_S0;		always @(posedge clk) O20_N8_S0 <=     O20_I18_R0_C0_SM1   +  O20_I21_R0_C0_SM1  ;
 logic signed [31:0] O20_N10_S0;		always @(posedge clk) O20_N10_S0 <=     O20_I22_R0_C0_SM1   +  O20_I23_R0_C0_SM1  ;
 logic signed [31:0] O20_N12_S0;		always @(posedge clk) O20_N12_S0 <=     O20_I24_R0_C0_SM1   +  O20_I25_R0_C0_SM1  ;
 logic signed [31:0] O20_N14_S0;		always @(posedge clk) O20_N14_S0 <=     O20_I28_R0_C0_SM1   +  O20_I30_R0_C0_SM1  ;
 logic signed [31:0] O20_N16_S0;		always @(posedge clk) O20_N16_S0 <=     O20_I31_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O20_N0_S1;		always @(posedge clk) O20_N0_S1 <=     O20_N0_S0  +  O20_N2_S0 ;
 logic signed [31:0] O20_N2_S1;		always @(posedge clk) O20_N2_S1 <=     O20_N4_S0  +  O20_N6_S0 ;
 logic signed [31:0] O20_N4_S1;		always @(posedge clk) O20_N4_S1 <=     O20_N8_S0  +  O20_N10_S0 ;
 logic signed [31:0] O20_N6_S1;		always @(posedge clk) O20_N6_S1 <=     O20_N12_S0  +  O20_N14_S0 ;
 logic signed [31:0] O20_N8_S1;		always @(posedge clk) O20_N8_S1 <=     O20_N16_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O20_N0_S2;		always @(posedge clk) O20_N0_S2 <=     O20_N0_S1  +  O20_N2_S1 ;
 logic signed [31:0] O20_N2_S2;		always @(posedge clk) O20_N2_S2 <=     O20_N4_S1  +  O20_N6_S1 ;
 logic signed [31:0] O20_N4_S2;		always @(posedge clk) O20_N4_S2 <=     O20_N8_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O20_N0_S3;		always @(posedge clk) O20_N0_S3 <=     O20_N0_S2  +  O20_N2_S2 ;
 logic signed [31:0] O20_N2_S3;		always @(posedge clk) O20_N2_S3 <=     O20_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O20_N0_S4;		always @(posedge clk) O20_N0_S4 <=     O20_N0_S3  +  O20_N2_S3 ;
 assign conv_mac_20 = O20_N0_S4;

logic signed [31:0] conv_mac_21;
logic signed [31:0] O21_N0_S0;		always @(posedge clk) O21_N0_S0 <=     O21_I0_R0_C0_SM1   +  O21_I1_R0_C0_SM1  ;
 logic signed [31:0] O21_N2_S0;		always @(posedge clk) O21_N2_S0 <=     O21_I2_R0_C0_SM1   +  O21_I3_R0_C0_SM1  ;
 logic signed [31:0] O21_N4_S0;		always @(posedge clk) O21_N4_S0 <=     O21_I4_R0_C0_SM1   +  O21_I5_R0_C0_SM1  ;
 logic signed [31:0] O21_N6_S0;		always @(posedge clk) O21_N6_S0 <=     O21_I6_R0_C0_SM1   +  O21_I7_R0_C0_SM1  ;
 logic signed [31:0] O21_N8_S0;		always @(posedge clk) O21_N8_S0 <=     O21_I8_R0_C0_SM1   +  O21_I9_R0_C0_SM1  ;
 logic signed [31:0] O21_N10_S0;		always @(posedge clk) O21_N10_S0 <=     O21_I10_R0_C0_SM1   +  O21_I13_R0_C0_SM1  ;
 logic signed [31:0] O21_N12_S0;		always @(posedge clk) O21_N12_S0 <=     O21_I16_R0_C0_SM1   +  O21_I17_R0_C0_SM1  ;
 logic signed [31:0] O21_N14_S0;		always @(posedge clk) O21_N14_S0 <=     O21_I18_R0_C0_SM1   +  O21_I19_R0_C0_SM1  ;
 logic signed [31:0] O21_N16_S0;		always @(posedge clk) O21_N16_S0 <=     O21_I21_R0_C0_SM1   +  O21_I22_R0_C0_SM1  ;
 logic signed [31:0] O21_N18_S0;		always @(posedge clk) O21_N18_S0 <=     O21_I24_R0_C0_SM1   +  O21_I25_R0_C0_SM1  ;
 logic signed [31:0] O21_N20_S0;		always @(posedge clk) O21_N20_S0 <=     O21_I27_R0_C0_SM1   +  O21_I28_R0_C0_SM1  ;
 logic signed [31:0] O21_N22_S0;		always @(posedge clk) O21_N22_S0 <=     O21_I29_R0_C0_SM1   +  O21_I30_R0_C0_SM1  ;
 logic signed [31:0] O21_N24_S0;		always @(posedge clk) O21_N24_S0 <=     O21_I31_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O21_N0_S1;		always @(posedge clk) O21_N0_S1 <=     O21_N0_S0  +  O21_N2_S0 ;
 logic signed [31:0] O21_N2_S1;		always @(posedge clk) O21_N2_S1 <=     O21_N4_S0  +  O21_N6_S0 ;
 logic signed [31:0] O21_N4_S1;		always @(posedge clk) O21_N4_S1 <=     O21_N8_S0  +  O21_N10_S0 ;
 logic signed [31:0] O21_N6_S1;		always @(posedge clk) O21_N6_S1 <=     O21_N12_S0  +  O21_N14_S0 ;
 logic signed [31:0] O21_N8_S1;		always @(posedge clk) O21_N8_S1 <=     O21_N16_S0  +  O21_N18_S0 ;
 logic signed [31:0] O21_N10_S1;		always @(posedge clk) O21_N10_S1 <=     O21_N20_S0  +  O21_N22_S0 ;
 logic signed [31:0] O21_N12_S1;		always @(posedge clk) O21_N12_S1 <=     O21_N24_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O21_N0_S2;		always @(posedge clk) O21_N0_S2 <=     O21_N0_S1  +  O21_N2_S1 ;
 logic signed [31:0] O21_N2_S2;		always @(posedge clk) O21_N2_S2 <=     O21_N4_S1  +  O21_N6_S1 ;
 logic signed [31:0] O21_N4_S2;		always @(posedge clk) O21_N4_S2 <=     O21_N8_S1  +  O21_N10_S1 ;
 logic signed [31:0] O21_N6_S2;		always @(posedge clk) O21_N6_S2 <=     O21_N12_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O21_N0_S3;		always @(posedge clk) O21_N0_S3 <=     O21_N0_S2  +  O21_N2_S2 ;
 logic signed [31:0] O21_N2_S3;		always @(posedge clk) O21_N2_S3 <=     O21_N4_S2  +  O21_N6_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O21_N0_S4;		always @(posedge clk) O21_N0_S4 <=     O21_N0_S3  +  O21_N2_S3 ;
 assign conv_mac_21 = O21_N0_S4;

logic signed [31:0] conv_mac_22;
logic signed [31:0] O22_N0_S0;		always @(posedge clk) O22_N0_S0 <=     O22_I2_R0_C0_SM1   +  O22_I3_R0_C0_SM1  ;
 logic signed [31:0] O22_N2_S0;		always @(posedge clk) O22_N2_S0 <=     O22_I6_R0_C0_SM1   +  O22_I7_R0_C0_SM1  ;
 logic signed [31:0] O22_N4_S0;		always @(posedge clk) O22_N4_S0 <=     O22_I8_R0_C0_SM1   +  O22_I10_R0_C0_SM1  ;
 logic signed [31:0] O22_N6_S0;		always @(posedge clk) O22_N6_S0 <=     O22_I12_R0_C0_SM1   +  O22_I14_R0_C0_SM1  ;
 logic signed [31:0] O22_N8_S0;		always @(posedge clk) O22_N8_S0 <=     O22_I15_R0_C0_SM1   +  O22_I17_R0_C0_SM1  ;
 logic signed [31:0] O22_N10_S0;		always @(posedge clk) O22_N10_S0 <=     O22_I18_R0_C0_SM1   +  O22_I20_R0_C0_SM1  ;
 logic signed [31:0] O22_N12_S0;		always @(posedge clk) O22_N12_S0 <=     O22_I22_R0_C0_SM1   +  O22_I23_R0_C0_SM1  ;
 logic signed [31:0] O22_N14_S0;		always @(posedge clk) O22_N14_S0 <=     O22_I25_R0_C0_SM1   +  O22_I27_R0_C0_SM1  ;
 logic signed [31:0] O22_N16_S0;		always @(posedge clk) O22_N16_S0 <=     O22_I28_R0_C0_SM1   +  O22_I29_R0_C0_SM1  ;
 logic signed [31:0] O22_N18_S0;		always @(posedge clk) O22_N18_S0 <=     O22_I30_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O22_N0_S1;		always @(posedge clk) O22_N0_S1 <=     O22_N0_S0  +  O22_N2_S0 ;
 logic signed [31:0] O22_N2_S1;		always @(posedge clk) O22_N2_S1 <=     O22_N4_S0  +  O22_N6_S0 ;
 logic signed [31:0] O22_N4_S1;		always @(posedge clk) O22_N4_S1 <=     O22_N8_S0  +  O22_N10_S0 ;
 logic signed [31:0] O22_N6_S1;		always @(posedge clk) O22_N6_S1 <=     O22_N12_S0  +  O22_N14_S0 ;
 logic signed [31:0] O22_N8_S1;		always @(posedge clk) O22_N8_S1 <=     O22_N16_S0  +  O22_N18_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O22_N0_S2;		always @(posedge clk) O22_N0_S2 <=     O22_N0_S1  +  O22_N2_S1 ;
 logic signed [31:0] O22_N2_S2;		always @(posedge clk) O22_N2_S2 <=     O22_N4_S1  +  O22_N6_S1 ;
 logic signed [31:0] O22_N4_S2;		always @(posedge clk) O22_N4_S2 <=     O22_N8_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O22_N0_S3;		always @(posedge clk) O22_N0_S3 <=     O22_N0_S2  +  O22_N2_S2 ;
 logic signed [31:0] O22_N2_S3;		always @(posedge clk) O22_N2_S3 <=     O22_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O22_N0_S4;		always @(posedge clk) O22_N0_S4 <=     O22_N0_S3  +  O22_N2_S3 ;
 assign conv_mac_22 = O22_N0_S4;

logic signed [31:0] conv_mac_23;
logic signed [31:0] O23_N0_S0;		always @(posedge clk) O23_N0_S0 <=     O23_I3_R0_C0_SM1   +  O23_I10_R0_C0_SM1  ;
 logic signed [31:0] O23_N2_S0;		always @(posedge clk) O23_N2_S0 <=     O23_I15_R0_C0_SM1   +  O23_I17_R0_C0_SM1  ;
 logic signed [31:0] O23_N4_S0;		always @(posedge clk) O23_N4_S0 <=     O23_I18_R0_C0_SM1   +  O23_I22_R0_C0_SM1  ;
 logic signed [31:0] O23_N6_S0;		always @(posedge clk) O23_N6_S0 <=     O23_I25_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O23_N0_S1;		always @(posedge clk) O23_N0_S1 <=     O23_N0_S0  +  O23_N2_S0 ;
 logic signed [31:0] O23_N2_S1;		always @(posedge clk) O23_N2_S1 <=     O23_N4_S0  +  O23_N6_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O23_N0_S2;		always @(posedge clk) O23_N0_S2 <=     O23_N0_S1  +  O23_N2_S1 ;
 assign conv_mac_23 = O23_N0_S2;

logic signed [31:0] conv_mac_24;
logic signed [31:0] O24_N0_S0;		always @(posedge clk) O24_N0_S0 <=     O24_I0_R0_C0_SM1   +  O24_I1_R0_C0_SM1  ;
 logic signed [31:0] O24_N2_S0;		always @(posedge clk) O24_N2_S0 <=     O24_I2_R0_C0_SM1   +  O24_I8_R0_C0_SM1  ;
 logic signed [31:0] O24_N4_S0;		always @(posedge clk) O24_N4_S0 <=     O24_I10_R0_C0_SM1   +  O24_I13_R0_C0_SM1  ;
 logic signed [31:0] O24_N6_S0;		always @(posedge clk) O24_N6_S0 <=     O24_I14_R0_C0_SM1   +  O24_I17_R0_C0_SM1  ;
 logic signed [31:0] O24_N8_S0;		always @(posedge clk) O24_N8_S0 <=     O24_I23_R0_C0_SM1   +  O24_I25_R0_C0_SM1  ;
 logic signed [31:0] O24_N10_S0;		always @(posedge clk) O24_N10_S0 <=     O24_I27_R0_C0_SM1   +  O24_I30_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O24_N0_S1;		always @(posedge clk) O24_N0_S1 <=     O24_N0_S0  +  O24_N2_S0 ;
 logic signed [31:0] O24_N2_S1;		always @(posedge clk) O24_N2_S1 <=     O24_N4_S0  +  O24_N6_S0 ;
 logic signed [31:0] O24_N4_S1;		always @(posedge clk) O24_N4_S1 <=     O24_N8_S0  +  O24_N10_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O24_N0_S2;		always @(posedge clk) O24_N0_S2 <=     O24_N0_S1  +  O24_N2_S1 ;
 logic signed [31:0] O24_N2_S2;		always @(posedge clk) O24_N2_S2 <=     O24_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O24_N0_S3;		always @(posedge clk) O24_N0_S3 <=     O24_N0_S2  +  O24_N2_S2 ;
 assign conv_mac_24 = O24_N0_S3;

logic signed [31:0] conv_mac_25;
logic signed [31:0] O25_N0_S0;		always @(posedge clk) O25_N0_S0 <=     O25_I1_R0_C0_SM1   +  O25_I2_R0_C0_SM1  ;
 logic signed [31:0] O25_N2_S0;		always @(posedge clk) O25_N2_S0 <=     O25_I7_R0_C0_SM1   +  O25_I9_R0_C0_SM1  ;
 logic signed [31:0] O25_N4_S0;		always @(posedge clk) O25_N4_S0 <=     O25_I12_R0_C0_SM1   +  O25_I13_R0_C0_SM1  ;
 logic signed [31:0] O25_N6_S0;		always @(posedge clk) O25_N6_S0 <=     O25_I15_R0_C0_SM1   +  O25_I17_R0_C0_SM1  ;
 logic signed [31:0] O25_N8_S0;		always @(posedge clk) O25_N8_S0 <=     O25_I20_R0_C0_SM1   +  O25_I25_R0_C0_SM1  ;
 logic signed [31:0] O25_N10_S0;		always @(posedge clk) O25_N10_S0 <=     O25_I27_R0_C0_SM1   +  O25_I28_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O25_N0_S1;		always @(posedge clk) O25_N0_S1 <=     O25_N0_S0  +  O25_N2_S0 ;
 logic signed [31:0] O25_N2_S1;		always @(posedge clk) O25_N2_S1 <=     O25_N4_S0  +  O25_N6_S0 ;
 logic signed [31:0] O25_N4_S1;		always @(posedge clk) O25_N4_S1 <=     O25_N8_S0  +  O25_N10_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O25_N0_S2;		always @(posedge clk) O25_N0_S2 <=     O25_N0_S1  +  O25_N2_S1 ;
 logic signed [31:0] O25_N2_S2;		always @(posedge clk) O25_N2_S2 <=     O25_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O25_N0_S3;		always @(posedge clk) O25_N0_S3 <=     O25_N0_S2  +  O25_N2_S2 ;
 assign conv_mac_25 = O25_N0_S3;

logic signed [31:0] conv_mac_26;
logic signed [31:0] O26_N0_S0;		always @(posedge clk) O26_N0_S0 <=     O26_I0_R0_C0_SM1   +  O26_I2_R0_C0_SM1  ;
 logic signed [31:0] O26_N2_S0;		always @(posedge clk) O26_N2_S0 <=     O26_I3_R0_C0_SM1   +  O26_I4_R0_C0_SM1  ;
 logic signed [31:0] O26_N4_S0;		always @(posedge clk) O26_N4_S0 <=     O26_I8_R0_C0_SM1   +  O26_I9_R0_C0_SM1  ;
 logic signed [31:0] O26_N6_S0;		always @(posedge clk) O26_N6_S0 <=     O26_I11_R0_C0_SM1   +  O26_I12_R0_C0_SM1  ;
 logic signed [31:0] O26_N8_S0;		always @(posedge clk) O26_N8_S0 <=     O26_I16_R0_C0_SM1   +  O26_I17_R0_C0_SM1  ;
 logic signed [31:0] O26_N10_S0;		always @(posedge clk) O26_N10_S0 <=     O26_I19_R0_C0_SM1   +  O26_I20_R0_C0_SM1  ;
 logic signed [31:0] O26_N12_S0;		always @(posedge clk) O26_N12_S0 <=     O26_I22_R0_C0_SM1   +  O26_I25_R0_C0_SM1  ;
 logic signed [31:0] O26_N14_S0;		always @(posedge clk) O26_N14_S0 <=     O26_I26_R0_C0_SM1   +  O26_I29_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O26_N0_S1;		always @(posedge clk) O26_N0_S1 <=     O26_N0_S0  +  O26_N2_S0 ;
 logic signed [31:0] O26_N2_S1;		always @(posedge clk) O26_N2_S1 <=     O26_N4_S0  +  O26_N6_S0 ;
 logic signed [31:0] O26_N4_S1;		always @(posedge clk) O26_N4_S1 <=     O26_N8_S0  +  O26_N10_S0 ;
 logic signed [31:0] O26_N6_S1;		always @(posedge clk) O26_N6_S1 <=     O26_N12_S0  +  O26_N14_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O26_N0_S2;		always @(posedge clk) O26_N0_S2 <=     O26_N0_S1  +  O26_N2_S1 ;
 logic signed [31:0] O26_N2_S2;		always @(posedge clk) O26_N2_S2 <=     O26_N4_S1  +  O26_N6_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O26_N0_S3;		always @(posedge clk) O26_N0_S3 <=     O26_N0_S2  +  O26_N2_S2 ;
 assign conv_mac_26 = O26_N0_S3;

logic signed [31:0] conv_mac_27;
logic signed [31:0] O27_N0_S0;		always @(posedge clk) O27_N0_S0 <=     O27_I0_R0_C0_SM1   +  O27_I3_R0_C0_SM1  ;
 logic signed [31:0] O27_N2_S0;		always @(posedge clk) O27_N2_S0 <=     O27_I4_R0_C0_SM1   +  O27_I5_R0_C0_SM1  ;
 logic signed [31:0] O27_N4_S0;		always @(posedge clk) O27_N4_S0 <=     O27_I8_R0_C0_SM1   +  O27_I9_R0_C0_SM1  ;
 logic signed [31:0] O27_N6_S0;		always @(posedge clk) O27_N6_S0 <=     O27_I12_R0_C0_SM1   +  O27_I13_R0_C0_SM1  ;
 logic signed [31:0] O27_N8_S0;		always @(posedge clk) O27_N8_S0 <=     O27_I18_R0_C0_SM1   +  O27_I19_R0_C0_SM1  ;
 logic signed [31:0] O27_N10_S0;		always @(posedge clk) O27_N10_S0 <=     O27_I21_R0_C0_SM1   +  O27_I22_R0_C0_SM1  ;
 logic signed [31:0] O27_N12_S0;		always @(posedge clk) O27_N12_S0 <=     O27_I23_R0_C0_SM1   +  O27_I26_R0_C0_SM1  ;
 logic signed [31:0] O27_N14_S0;		always @(posedge clk) O27_N14_S0 <=     O27_I29_R0_C0_SM1   +  O27_I30_R0_C0_SM1  ;
 logic signed [31:0] O27_N16_S0;		always @(posedge clk) O27_N16_S0 <=     O27_I31_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O27_N0_S1;		always @(posedge clk) O27_N0_S1 <=     O27_N0_S0  +  O27_N2_S0 ;
 logic signed [31:0] O27_N2_S1;		always @(posedge clk) O27_N2_S1 <=     O27_N4_S0  +  O27_N6_S0 ;
 logic signed [31:0] O27_N4_S1;		always @(posedge clk) O27_N4_S1 <=     O27_N8_S0  +  O27_N10_S0 ;
 logic signed [31:0] O27_N6_S1;		always @(posedge clk) O27_N6_S1 <=     O27_N12_S0  +  O27_N14_S0 ;
 logic signed [31:0] O27_N8_S1;		always @(posedge clk) O27_N8_S1 <=     O27_N16_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O27_N0_S2;		always @(posedge clk) O27_N0_S2 <=     O27_N0_S1  +  O27_N2_S1 ;
 logic signed [31:0] O27_N2_S2;		always @(posedge clk) O27_N2_S2 <=     O27_N4_S1  +  O27_N6_S1 ;
 logic signed [31:0] O27_N4_S2;		always @(posedge clk) O27_N4_S2 <=     O27_N8_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O27_N0_S3;		always @(posedge clk) O27_N0_S3 <=     O27_N0_S2  +  O27_N2_S2 ;
 logic signed [31:0] O27_N2_S3;		always @(posedge clk) O27_N2_S3 <=     O27_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O27_N0_S4;		always @(posedge clk) O27_N0_S4 <=     O27_N0_S3  +  O27_N2_S3 ;
 assign conv_mac_27 = O27_N0_S4;

logic signed [31:0] conv_mac_28;
logic signed [31:0] O28_N0_S0;		always @(posedge clk) O28_N0_S0 <=     O28_I0_R0_C0_SM1   +  O28_I1_R0_C0_SM1  ;
 logic signed [31:0] O28_N2_S0;		always @(posedge clk) O28_N2_S0 <=     O28_I2_R0_C0_SM1   +  O28_I6_R0_C0_SM1  ;
 logic signed [31:0] O28_N4_S0;		always @(posedge clk) O28_N4_S0 <=     O28_I7_R0_C0_SM1   +  O28_I8_R0_C0_SM1  ;
 logic signed [31:0] O28_N6_S0;		always @(posedge clk) O28_N6_S0 <=     O28_I9_R0_C0_SM1   +  O28_I14_R0_C0_SM1  ;
 logic signed [31:0] O28_N8_S0;		always @(posedge clk) O28_N8_S0 <=     O28_I15_R0_C0_SM1   +  O28_I16_R0_C0_SM1  ;
 logic signed [31:0] O28_N10_S0;		always @(posedge clk) O28_N10_S0 <=     O28_I18_R0_C0_SM1   +  O28_I21_R0_C0_SM1  ;
 logic signed [31:0] O28_N12_S0;		always @(posedge clk) O28_N12_S0 <=     O28_I22_R0_C0_SM1   +  O28_I23_R0_C0_SM1  ;
 logic signed [31:0] O28_N14_S0;		always @(posedge clk) O28_N14_S0 <=     O28_I24_R0_C0_SM1   +  O28_I25_R0_C0_SM1  ;
 logic signed [31:0] O28_N16_S0;		always @(posedge clk) O28_N16_S0 <=     O28_I27_R0_C0_SM1   +  O28_I28_R0_C0_SM1  ;
 logic signed [31:0] O28_N18_S0;		always @(posedge clk) O28_N18_S0 <=     O28_I30_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O28_N0_S1;		always @(posedge clk) O28_N0_S1 <=     O28_N0_S0  +  O28_N2_S0 ;
 logic signed [31:0] O28_N2_S1;		always @(posedge clk) O28_N2_S1 <=     O28_N4_S0  +  O28_N6_S0 ;
 logic signed [31:0] O28_N4_S1;		always @(posedge clk) O28_N4_S1 <=     O28_N8_S0  +  O28_N10_S0 ;
 logic signed [31:0] O28_N6_S1;		always @(posedge clk) O28_N6_S1 <=     O28_N12_S0  +  O28_N14_S0 ;
 logic signed [31:0] O28_N8_S1;		always @(posedge clk) O28_N8_S1 <=     O28_N16_S0  +  O28_N18_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O28_N0_S2;		always @(posedge clk) O28_N0_S2 <=     O28_N0_S1  +  O28_N2_S1 ;
 logic signed [31:0] O28_N2_S2;		always @(posedge clk) O28_N2_S2 <=     O28_N4_S1  +  O28_N6_S1 ;
 logic signed [31:0] O28_N4_S2;		always @(posedge clk) O28_N4_S2 <=     O28_N8_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O28_N0_S3;		always @(posedge clk) O28_N0_S3 <=     O28_N0_S2  +  O28_N2_S2 ;
 logic signed [31:0] O28_N2_S3;		always @(posedge clk) O28_N2_S3 <=     O28_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O28_N0_S4;		always @(posedge clk) O28_N0_S4 <=     O28_N0_S3  +  O28_N2_S3 ;
 assign conv_mac_28 = O28_N0_S4;

logic signed [31:0] conv_mac_29;
logic signed [31:0] O29_N0_S0;		always @(posedge clk) O29_N0_S0 <=     O29_I0_R0_C0_SM1   +  O29_I1_R0_C0_SM1  ;
 logic signed [31:0] O29_N2_S0;		always @(posedge clk) O29_N2_S0 <=     O29_I2_R0_C0_SM1   +  O29_I3_R0_C0_SM1  ;
 logic signed [31:0] O29_N4_S0;		always @(posedge clk) O29_N4_S0 <=     O29_I4_R0_C0_SM1   +  O29_I5_R0_C0_SM1  ;
 logic signed [31:0] O29_N6_S0;		always @(posedge clk) O29_N6_S0 <=     O29_I6_R0_C0_SM1   +  O29_I8_R0_C0_SM1  ;
 logic signed [31:0] O29_N8_S0;		always @(posedge clk) O29_N8_S0 <=     O29_I11_R0_C0_SM1   +  O29_I12_R0_C0_SM1  ;
 logic signed [31:0] O29_N10_S0;		always @(posedge clk) O29_N10_S0 <=     O29_I13_R0_C0_SM1   +  O29_I16_R0_C0_SM1  ;
 logic signed [31:0] O29_N12_S0;		always @(posedge clk) O29_N12_S0 <=     O29_I17_R0_C0_SM1   +  O29_I19_R0_C0_SM1  ;
 logic signed [31:0] O29_N14_S0;		always @(posedge clk) O29_N14_S0 <=     O29_I20_R0_C0_SM1   +  O29_I21_R0_C0_SM1  ;
 logic signed [31:0] O29_N16_S0;		always @(posedge clk) O29_N16_S0 <=     O29_I24_R0_C0_SM1   +  O29_I26_R0_C0_SM1  ;
 logic signed [31:0] O29_N18_S0;		always @(posedge clk) O29_N18_S0 <=     O29_I27_R0_C0_SM1   +  O29_I29_R0_C0_SM1  ;
 logic signed [31:0] O29_N20_S0;		always @(posedge clk) O29_N20_S0 <=     O29_I30_R0_C0_SM1   +  O29_I31_R0_C0_SM1  ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O29_N0_S1;		always @(posedge clk) O29_N0_S1 <=     O29_N0_S0  +  O29_N2_S0 ;
 logic signed [31:0] O29_N2_S1;		always @(posedge clk) O29_N2_S1 <=     O29_N4_S0  +  O29_N6_S0 ;
 logic signed [31:0] O29_N4_S1;		always @(posedge clk) O29_N4_S1 <=     O29_N8_S0  +  O29_N10_S0 ;
 logic signed [31:0] O29_N6_S1;		always @(posedge clk) O29_N6_S1 <=     O29_N12_S0  +  O29_N14_S0 ;
 logic signed [31:0] O29_N8_S1;		always @(posedge clk) O29_N8_S1 <=     O29_N16_S0  +  O29_N18_S0 ;
 logic signed [31:0] O29_N10_S1;		always @(posedge clk) O29_N10_S1 <=     O29_N20_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O29_N0_S2;		always @(posedge clk) O29_N0_S2 <=     O29_N0_S1  +  O29_N2_S1 ;
 logic signed [31:0] O29_N2_S2;		always @(posedge clk) O29_N2_S2 <=     O29_N4_S1  +  O29_N6_S1 ;
 logic signed [31:0] O29_N4_S2;		always @(posedge clk) O29_N4_S2 <=     O29_N8_S1  +  O29_N10_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O29_N0_S3;		always @(posedge clk) O29_N0_S3 <=     O29_N0_S2  +  O29_N2_S2 ;
 logic signed [31:0] O29_N2_S3;		always @(posedge clk) O29_N2_S3 <=     O29_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O29_N0_S4;		always @(posedge clk) O29_N0_S4 <=     O29_N0_S3  +  O29_N2_S3 ;
 assign conv_mac_29 = O29_N0_S4;

logic signed [31:0] conv_mac_30;
logic signed [31:0] O30_N0_S0;		always @(posedge clk) O30_N0_S0 <=     O30_I0_R0_C0_SM1   +  O30_I1_R0_C0_SM1  ;
 logic signed [31:0] O30_N2_S0;		always @(posedge clk) O30_N2_S0 <=     O30_I2_R0_C0_SM1   +  O30_I3_R0_C0_SM1  ;
 logic signed [31:0] O30_N4_S0;		always @(posedge clk) O30_N4_S0 <=     O30_I5_R0_C0_SM1   +  O30_I6_R0_C0_SM1  ;
 logic signed [31:0] O30_N6_S0;		always @(posedge clk) O30_N6_S0 <=     O30_I10_R0_C0_SM1   +  O30_I11_R0_C0_SM1  ;
 logic signed [31:0] O30_N8_S0;		always @(posedge clk) O30_N8_S0 <=     O30_I13_R0_C0_SM1   +  O30_I14_R0_C0_SM1  ;
 logic signed [31:0] O30_N10_S0;		always @(posedge clk) O30_N10_S0 <=     O30_I15_R0_C0_SM1   +  O30_I16_R0_C0_SM1  ;
 logic signed [31:0] O30_N12_S0;		always @(posedge clk) O30_N12_S0 <=     O30_I17_R0_C0_SM1   +  O30_I18_R0_C0_SM1  ;
 logic signed [31:0] O30_N14_S0;		always @(posedge clk) O30_N14_S0 <=     O30_I21_R0_C0_SM1   +  O30_I22_R0_C0_SM1  ;
 logic signed [31:0] O30_N16_S0;		always @(posedge clk) O30_N16_S0 <=     O30_I24_R0_C0_SM1   +  O30_I25_R0_C0_SM1  ;
 logic signed [31:0] O30_N18_S0;		always @(posedge clk) O30_N18_S0 <=     O30_I27_R0_C0_SM1   +  O30_I29_R0_C0_SM1  ;
 logic signed [31:0] O30_N20_S0;		always @(posedge clk) O30_N20_S0 <=     O30_I31_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O30_N0_S1;		always @(posedge clk) O30_N0_S1 <=     O30_N0_S0  +  O30_N2_S0 ;
 logic signed [31:0] O30_N2_S1;		always @(posedge clk) O30_N2_S1 <=     O30_N4_S0  +  O30_N6_S0 ;
 logic signed [31:0] O30_N4_S1;		always @(posedge clk) O30_N4_S1 <=     O30_N8_S0  +  O30_N10_S0 ;
 logic signed [31:0] O30_N6_S1;		always @(posedge clk) O30_N6_S1 <=     O30_N12_S0  +  O30_N14_S0 ;
 logic signed [31:0] O30_N8_S1;		always @(posedge clk) O30_N8_S1 <=     O30_N16_S0  +  O30_N18_S0 ;
 logic signed [31:0] O30_N10_S1;		always @(posedge clk) O30_N10_S1 <=     O30_N20_S0     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O30_N0_S2;		always @(posedge clk) O30_N0_S2 <=     O30_N0_S1  +  O30_N2_S1 ;
 logic signed [31:0] O30_N2_S2;		always @(posedge clk) O30_N2_S2 <=     O30_N4_S1  +  O30_N6_S1 ;
 logic signed [31:0] O30_N4_S2;		always @(posedge clk) O30_N4_S2 <=     O30_N8_S1  +  O30_N10_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O30_N0_S3;		always @(posedge clk) O30_N0_S3 <=     O30_N0_S2  +  O30_N2_S2 ;
 logic signed [31:0] O30_N2_S3;		always @(posedge clk) O30_N2_S3 <=     O30_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O30_N0_S4;		always @(posedge clk) O30_N0_S4 <=     O30_N0_S3  +  O30_N2_S3 ;
 assign conv_mac_30 = O30_N0_S4;

logic signed [31:0] conv_mac_31;
logic signed [31:0] O31_N0_S0;		always @(posedge clk) O31_N0_S0 <=     O31_I0_R0_C0_SM1   +  O31_I1_R0_C0_SM1  ;
 logic signed [31:0] O31_N2_S0;		always @(posedge clk) O31_N2_S0 <=     O31_I2_R0_C0_SM1   +  O31_I3_R0_C0_SM1  ;
 logic signed [31:0] O31_N4_S0;		always @(posedge clk) O31_N4_S0 <=     O31_I4_R0_C0_SM1   +  O31_I6_R0_C0_SM1  ;
 logic signed [31:0] O31_N6_S0;		always @(posedge clk) O31_N6_S0 <=     O31_I7_R0_C0_SM1   +  O31_I12_R0_C0_SM1  ;
 logic signed [31:0] O31_N8_S0;		always @(posedge clk) O31_N8_S0 <=     O31_I13_R0_C0_SM1   +  O31_I16_R0_C0_SM1  ;
 logic signed [31:0] O31_N10_S0;		always @(posedge clk) O31_N10_S0 <=     O31_I17_R0_C0_SM1   +  O31_I19_R0_C0_SM1  ;
 logic signed [31:0] O31_N12_S0;		always @(posedge clk) O31_N12_S0 <=     O31_I28_R0_C0_SM1   +  O31_I30_R0_C0_SM1  ;
 logic signed [31:0] O31_N14_S0;		always @(posedge clk) O31_N14_S0 <=     O31_I31_R0_C0_SM1      ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O31_N0_S1;		always @(posedge clk) O31_N0_S1 <=     O31_N0_S0  +  O31_N2_S0 ;
 logic signed [31:0] O31_N2_S1;		always @(posedge clk) O31_N2_S1 <=     O31_N4_S0  +  O31_N6_S0 ;
 logic signed [31:0] O31_N4_S1;		always @(posedge clk) O31_N4_S1 <=     O31_N8_S0  +  O31_N10_S0 ;
 logic signed [31:0] O31_N6_S1;		always @(posedge clk) O31_N6_S1 <=     O31_N12_S0  +  O31_N14_S0 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O31_N0_S2;		always @(posedge clk) O31_N0_S2 <=     O31_N0_S1  +  O31_N2_S1 ;
 logic signed [31:0] O31_N2_S2;		always @(posedge clk) O31_N2_S2 <=     O31_N4_S1  +  O31_N6_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [31:0] O31_N0_S3;		always @(posedge clk) O31_N0_S3 <=     O31_N0_S2  +  O31_N2_S2 ;
 assign conv_mac_31 = O31_N0_S3;

logic valid_D1;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D1<= 0 ;
	else valid_D1<=valid;
end
logic valid_D2;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D2<= 0 ;
	else valid_D2<=valid_D1;
end
logic valid_D3;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D3<= 0 ;
	else valid_D3<=valid_D2;
end
logic valid_D4;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D4<= 0 ;
	else valid_D4<=valid_D3;
end
logic valid_D5;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D5<= 0 ;
	else valid_D5<=valid_D4;
end
logic valid_D6;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D6<= 0 ;
	else valid_D6<=valid_D5;
end
always_ff @(posedge clk) begin
	if (rstn == 0) ready <= 0 ;
	else ready <=valid_D6;
end
logic [31:0] bias_add_0;
assign bias_add_0 = conv_mac_0 + 6'd20;
logic [31:0] bias_add_1;
assign bias_add_1 = conv_mac_1 + 6'd18;
logic [31:0] bias_add_2;
assign bias_add_2 = conv_mac_2 + 6'd21;
logic [31:0] bias_add_3;
assign bias_add_3 = conv_mac_3 - 5'd10;
logic [31:0] bias_add_4;
assign bias_add_4 = conv_mac_4 - 4'd7;
logic [31:0] bias_add_5;
assign bias_add_5 = conv_mac_5 - 5'd11;
logic [31:0] bias_add_6;
assign bias_add_6 = conv_mac_6 + 5'd14;
logic [31:0] bias_add_7;
assign bias_add_7 = conv_mac_7 + 4'd6;
logic [31:0] bias_add_8;
assign bias_add_8 = conv_mac_8;
logic [31:0] bias_add_9;
assign bias_add_9 = conv_mac_9 - 6'd18;
logic [31:0] bias_add_10;
assign bias_add_10 = conv_mac_10 - 3'd2;
logic [31:0] bias_add_11;
assign bias_add_11 = conv_mac_11 - 6'd20;
logic [31:0] bias_add_12;
assign bias_add_12 = conv_mac_12 - 3'd3;
logic [31:0] bias_add_13;
assign bias_add_13 = conv_mac_13 + 6'd16;
logic [31:0] bias_add_14;
assign bias_add_14 = conv_mac_14 + 6'd21;
logic [31:0] bias_add_15;
assign bias_add_15 = conv_mac_15 + 4'd7;
logic [31:0] bias_add_16;
assign bias_add_16 = conv_mac_16 + 4'd6;
logic [31:0] bias_add_17;
assign bias_add_17 = conv_mac_17 + 7'd32;
logic [31:0] bias_add_18;
assign bias_add_18 = conv_mac_18 + 6'd16;
logic [31:0] bias_add_19;
assign bias_add_19 = conv_mac_19 + 6'd24;
logic [31:0] bias_add_20;
assign bias_add_20 = conv_mac_20 + 6'd30;
logic [31:0] bias_add_21;
assign bias_add_21 = conv_mac_21 - 5'd10;
logic [31:0] bias_add_22;
assign bias_add_22 = conv_mac_22 + 5'd13;
logic [31:0] bias_add_23;
assign bias_add_23 = conv_mac_23 + 4'd4;
logic [31:0] bias_add_24;
assign bias_add_24 = conv_mac_24 + 3'd3;
logic [31:0] bias_add_25;
assign bias_add_25 = conv_mac_25 + 6'd28;
logic [31:0] bias_add_26;
assign bias_add_26 = conv_mac_26 - 4'd5;
logic [31:0] bias_add_27;
assign bias_add_27 = conv_mac_27 + 3'd3;
logic [31:0] bias_add_28;
assign bias_add_28 = conv_mac_28 + 6'd29;
logic [31:0] bias_add_29;
assign bias_add_29 = conv_mac_29 - 6'd16;
logic [31:0] bias_add_30;
assign bias_add_30 = conv_mac_30 + 4'd6;
logic [31:0] bias_add_31;
assign bias_add_31 = conv_mac_31 + 5'd9;

logic [7:0] relu_0;
assign relu_0[7:0] = (bias_add_0[31]==0) ? ((bias_add_0<3'd6) ? {{bias_add_0[31],bias_add_0[10:4]}} :'d6) : '0;
logic [7:0] relu_1;
assign relu_1[7:0] = (bias_add_1[31]==0) ? ((bias_add_1<3'd6) ? {{bias_add_1[31],bias_add_1[10:4]}} :'d6) : '0;
logic [7:0] relu_2;
assign relu_2[7:0] = (bias_add_2[31]==0) ? ((bias_add_2<3'd6) ? {{bias_add_2[31],bias_add_2[10:4]}} :'d6) : '0;
logic [7:0] relu_3;
assign relu_3[7:0] = (bias_add_3[31]==0) ? ((bias_add_3<3'd6) ? {{bias_add_3[31],bias_add_3[10:4]}} :'d6) : '0;
logic [7:0] relu_4;
assign relu_4[7:0] = (bias_add_4[31]==0) ? ((bias_add_4<3'd6) ? {{bias_add_4[31],bias_add_4[10:4]}} :'d6) : '0;
logic [7:0] relu_5;
assign relu_5[7:0] = (bias_add_5[31]==0) ? ((bias_add_5<3'd6) ? {{bias_add_5[31],bias_add_5[10:4]}} :'d6) : '0;
logic [7:0] relu_6;
assign relu_6[7:0] = (bias_add_6[31]==0) ? ((bias_add_6<3'd6) ? {{bias_add_6[31],bias_add_6[10:4]}} :'d6) : '0;
logic [7:0] relu_7;
assign relu_7[7:0] = (bias_add_7[31]==0) ? ((bias_add_7<3'd6) ? {{bias_add_7[31],bias_add_7[10:4]}} :'d6) : '0;
logic [7:0] relu_8;
assign relu_8[7:0] = (bias_add_8[31]==0) ? ((bias_add_8<3'd6) ? {{bias_add_8[31],bias_add_8[10:4]}} :'d6) : '0;
logic [7:0] relu_9;
assign relu_9[7:0] = (bias_add_9[31]==0) ? ((bias_add_9<3'd6) ? {{bias_add_9[31],bias_add_9[10:4]}} :'d6) : '0;
logic [7:0] relu_10;
assign relu_10[7:0] = (bias_add_10[31]==0) ? ((bias_add_10<3'd6) ? {{bias_add_10[31],bias_add_10[10:4]}} :'d6) : '0;
logic [7:0] relu_11;
assign relu_11[7:0] = (bias_add_11[31]==0) ? ((bias_add_11<3'd6) ? {{bias_add_11[31],bias_add_11[10:4]}} :'d6) : '0;
logic [7:0] relu_12;
assign relu_12[7:0] = (bias_add_12[31]==0) ? ((bias_add_12<3'd6) ? {{bias_add_12[31],bias_add_12[10:4]}} :'d6) : '0;
logic [7:0] relu_13;
assign relu_13[7:0] = (bias_add_13[31]==0) ? ((bias_add_13<3'd6) ? {{bias_add_13[31],bias_add_13[10:4]}} :'d6) : '0;
logic [7:0] relu_14;
assign relu_14[7:0] = (bias_add_14[31]==0) ? ((bias_add_14<3'd6) ? {{bias_add_14[31],bias_add_14[10:4]}} :'d6) : '0;
logic [7:0] relu_15;
assign relu_15[7:0] = (bias_add_15[31]==0) ? ((bias_add_15<3'd6) ? {{bias_add_15[31],bias_add_15[10:4]}} :'d6) : '0;
logic [7:0] relu_16;
assign relu_16[7:0] = (bias_add_16[31]==0) ? ((bias_add_16<3'd6) ? {{bias_add_16[31],bias_add_16[10:4]}} :'d6) : '0;
logic [7:0] relu_17;
assign relu_17[7:0] = (bias_add_17[31]==0) ? ((bias_add_17<3'd6) ? {{bias_add_17[31],bias_add_17[10:4]}} :'d6) : '0;
logic [7:0] relu_18;
assign relu_18[7:0] = (bias_add_18[31]==0) ? ((bias_add_18<3'd6) ? {{bias_add_18[31],bias_add_18[10:4]}} :'d6) : '0;
logic [7:0] relu_19;
assign relu_19[7:0] = (bias_add_19[31]==0) ? ((bias_add_19<3'd6) ? {{bias_add_19[31],bias_add_19[10:4]}} :'d6) : '0;
logic [7:0] relu_20;
assign relu_20[7:0] = (bias_add_20[31]==0) ? ((bias_add_20<3'd6) ? {{bias_add_20[31],bias_add_20[10:4]}} :'d6) : '0;
logic [7:0] relu_21;
assign relu_21[7:0] = (bias_add_21[31]==0) ? ((bias_add_21<3'd6) ? {{bias_add_21[31],bias_add_21[10:4]}} :'d6) : '0;
logic [7:0] relu_22;
assign relu_22[7:0] = (bias_add_22[31]==0) ? ((bias_add_22<3'd6) ? {{bias_add_22[31],bias_add_22[10:4]}} :'d6) : '0;
logic [7:0] relu_23;
assign relu_23[7:0] = (bias_add_23[31]==0) ? ((bias_add_23<3'd6) ? {{bias_add_23[31],bias_add_23[10:4]}} :'d6) : '0;
logic [7:0] relu_24;
assign relu_24[7:0] = (bias_add_24[31]==0) ? ((bias_add_24<3'd6) ? {{bias_add_24[31],bias_add_24[10:4]}} :'d6) : '0;
logic [7:0] relu_25;
assign relu_25[7:0] = (bias_add_25[31]==0) ? ((bias_add_25<3'd6) ? {{bias_add_25[31],bias_add_25[10:4]}} :'d6) : '0;
logic [7:0] relu_26;
assign relu_26[7:0] = (bias_add_26[31]==0) ? ((bias_add_26<3'd6) ? {{bias_add_26[31],bias_add_26[10:4]}} :'d6) : '0;
logic [7:0] relu_27;
assign relu_27[7:0] = (bias_add_27[31]==0) ? ((bias_add_27<3'd6) ? {{bias_add_27[31],bias_add_27[10:4]}} :'d6) : '0;
logic [7:0] relu_28;
assign relu_28[7:0] = (bias_add_28[31]==0) ? ((bias_add_28<3'd6) ? {{bias_add_28[31],bias_add_28[10:4]}} :'d6) : '0;
logic [7:0] relu_29;
assign relu_29[7:0] = (bias_add_29[31]==0) ? ((bias_add_29<3'd6) ? {{bias_add_29[31],bias_add_29[10:4]}} :'d6) : '0;
logic [7:0] relu_30;
assign relu_30[7:0] = (bias_add_30[31]==0) ? ((bias_add_30<3'd6) ? {{bias_add_30[31],bias_add_30[10:4]}} :'d6) : '0;
logic [7:0] relu_31;
assign relu_31[7:0] = (bias_add_31[31]==0) ? ((bias_add_31<3'd6) ? {{bias_add_31[31],bias_add_31[10:4]}} :'d6) : '0;

assign output_act = {
	relu_31,
	relu_30,
	relu_29,
	relu_28,
	relu_27,
	relu_26,
	relu_25,
	relu_24,
	relu_23,
	relu_22,
	relu_21,
	relu_20,
	relu_19,
	relu_18,
	relu_17,
	relu_16,
	relu_15,
	relu_14,
	relu_13,
	relu_12,
	relu_11,
	relu_10,
	relu_9,
	relu_8,
	relu_7,
	relu_6,
	relu_5,
	relu_4,
	relu_3,
	relu_2,
	relu_1,
	relu_0
};

endmodule
module conv6_pw (
    input logic clk,
    input logic rstn,
    input logic valid,
    input logic [256-1:0] input_act,
    output logic [512-1:0] output_act,
    output logic ready
);
logic we;
logic [8:0] zero_number; 
assign zero_number = 9'd0; 
//1
logic [256-1:0] input_act_ff ;
always_ff @(posedge clk) begin
    if (rstn == 0) begin
        input_act_ff <= '0;
      //  ready <= '0;
    end
    else begin
        input_act_ff <= input_act;
     //   ready <= valid;
    end
end
logic [7:0] input_fmap_0;
assign input_fmap_0 = input_act_ff[7:0];
logic [7:0] input_fmap_1;
assign input_fmap_1 = input_act_ff[15:8];
logic [7:0] input_fmap_2;
assign input_fmap_2 = input_act_ff[23:16];
logic [7:0] input_fmap_3;
assign input_fmap_3 = input_act_ff[31:24];
logic [7:0] input_fmap_4;
assign input_fmap_4 = input_act_ff[39:32];
logic [7:0] input_fmap_5;
assign input_fmap_5 = input_act_ff[47:40];
logic [7:0] input_fmap_6;
assign input_fmap_6 = input_act_ff[55:48];
logic [7:0] input_fmap_7;
assign input_fmap_7 = input_act_ff[63:56];
logic [7:0] input_fmap_8;
assign input_fmap_8 = input_act_ff[71:64];
logic [7:0] input_fmap_9;
assign input_fmap_9 = input_act_ff[79:72];
logic [7:0] input_fmap_10;
assign input_fmap_10 = input_act_ff[87:80];
logic [7:0] input_fmap_11;
assign input_fmap_11 = input_act_ff[95:88];
logic [7:0] input_fmap_12;
assign input_fmap_12 = input_act_ff[103:96];
logic [7:0] input_fmap_13;
assign input_fmap_13 = input_act_ff[111:104];
logic [7:0] input_fmap_14;
assign input_fmap_14 = input_act_ff[119:112];
logic [7:0] input_fmap_15;
assign input_fmap_15 = input_act_ff[127:120];
logic [7:0] input_fmap_16;
assign input_fmap_16 = input_act_ff[135:128];
logic [7:0] input_fmap_17;
assign input_fmap_17 = input_act_ff[143:136];
logic [7:0] input_fmap_18;
assign input_fmap_18 = input_act_ff[151:144];
logic [7:0] input_fmap_19;
assign input_fmap_19 = input_act_ff[159:152];
logic [7:0] input_fmap_20;
assign input_fmap_20 = input_act_ff[167:160];
logic [7:0] input_fmap_21;
assign input_fmap_21 = input_act_ff[175:168];
logic [7:0] input_fmap_22;
assign input_fmap_22 = input_act_ff[183:176];
logic [7:0] input_fmap_23;
assign input_fmap_23 = input_act_ff[191:184];
logic [7:0] input_fmap_24;
assign input_fmap_24 = input_act_ff[199:192];
logic [7:0] input_fmap_25;
assign input_fmap_25 = input_act_ff[207:200];
logic [7:0] input_fmap_26;
assign input_fmap_26 = input_act_ff[215:208];
logic [7:0] input_fmap_27;
assign input_fmap_27 = input_act_ff[223:216];
logic [7:0] input_fmap_28;
assign input_fmap_28 = input_act_ff[231:224];
logic [7:0] input_fmap_29;
assign input_fmap_29 = input_act_ff[239:232];
logic [7:0] input_fmap_30;
assign input_fmap_30 = input_act_ff[247:240];
logic [7:0] input_fmap_31;
assign input_fmap_31 = input_act_ff[255:248];

logic signed [31:0] conv_mac_0;
logic signed [63:0] chainout_0_O0; 
logic signed [63:0] O0_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O0(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd4),.bx(input_fmap_1[7:0]),.by( 9'sd1),.cx(input_fmap_3[7:0]),.cy(-9'sd1),.dx(input_fmap_4[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O0_N0_S1),.chainout(chainout_0_O0));
logic signed [63:0] chainout_2_O0; 
logic signed [63:0] O0_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O0(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_5[7:0]),.ay( 9'sd1),.bx(input_fmap_6[7:0]),.by( 9'sd1),.cx(input_fmap_8[7:0]),.cy( 9'sd1),.dx(input_fmap_10[7:0]),.dy( 9'sd3),.chainin(63'd0),.result(O0_N2_S1),.chainout(chainout_2_O0));
logic signed [63:0] chainout_4_O0; 
logic signed [63:0] O0_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O0(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_11[7:0]),.ay(-9'sd5),.bx(input_fmap_13[7:0]),.by(-9'sd2),.cx(input_fmap_14[7:0]),.cy(-9'sd1),.dx(input_fmap_15[7:0]),.dy(-9'sd3),.chainin(63'd0),.result(O0_N4_S1),.chainout(chainout_4_O0));
logic signed [63:0] chainout_6_O0; 
logic signed [63:0] O0_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O0(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_20[7:0]),.ay( 9'sd1),.bx(input_fmap_21[7:0]),.by(-9'sd2),.cx(input_fmap_23[7:0]),.cy( 9'sd1),.dx(input_fmap_24[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O0_N6_S1),.chainout(chainout_6_O0));
logic signed [63:0] chainout_8_O0; 
logic signed [63:0] O0_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O0(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_26[7:0]),.ay( 9'sd5),.bx(input_fmap_27[7:0]),.by(-9'sd3),.cx(input_fmap_29[7:0]),.cy(-9'sd1),.dx(input_fmap_30[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O0_N8_S1),.chainout(chainout_8_O0));
logic signed [63:0] chainout_10_O0; 
logic signed [63:0] O0_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O0(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_31[7:0]),.ay(-9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O0_N10_S1),.chainout(chainout_10_O0));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O0_N0_S2;		always @(posedge clk) O0_N0_S2 <=     O0_N0_S1  +  O0_N2_S1 ;
 logic signed [21:0] O0_N2_S2;		always @(posedge clk) O0_N2_S2 <=     O0_N4_S1  +  O0_N6_S1 ;
 logic signed [21:0] O0_N4_S2;		always @(posedge clk) O0_N4_S2 <=     O0_N8_S1  +  O0_N10_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O0_N0_S3;		always @(posedge clk) O0_N0_S3 <=     O0_N0_S2  +  O0_N2_S2 ;
 logic signed [22:0] O0_N2_S3;		always @(posedge clk) O0_N2_S3 <=     O0_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O0_N0_S4;		always @(posedge clk) O0_N0_S4 <=     O0_N0_S3  +  O0_N2_S3 ;
 assign conv_mac_0 = O0_N0_S4;

logic signed [31:0] conv_mac_1;
logic signed [63:0] chainout_0_O1; 
logic signed [63:0] O1_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O1(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_2[7:0]),.ay( 9'sd1),.bx(input_fmap_3[7:0]),.by( 9'sd1),.cx(input_fmap_7[7:0]),.cy( 9'sd3),.dx(input_fmap_11[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O1_N0_S1),.chainout(chainout_0_O1));
logic signed [63:0] chainout_2_O1; 
logic signed [63:0] O1_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O1(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_12[7:0]),.ay( 9'sd1),.bx(input_fmap_17[7:0]),.by(-9'sd1),.cx(input_fmap_25[7:0]),.cy(-9'sd1),.dx(input_fmap_28[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O1_N2_S1),.chainout(chainout_2_O1));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O1_N0_S2;		always @(posedge clk) O1_N0_S2 <=     O1_N0_S1  +  O1_N2_S1 ;
 assign conv_mac_1 = O1_N0_S2;

logic signed [31:0] conv_mac_2;
logic signed [63:0] chainout_0_O2; 
logic signed [63:0] O2_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O2(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay(-9'sd1),.bx(input_fmap_7[7:0]),.by(-9'sd1),.cx(input_fmap_10[7:0]),.cy(-9'sd1),.dx(input_fmap_11[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O2_N0_S1),.chainout(chainout_0_O2));
logic signed [63:0] chainout_2_O2; 
logic signed [63:0] O2_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O2(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_12[7:0]),.ay(-9'sd1),.bx(input_fmap_13[7:0]),.by( 9'sd2),.cx(input_fmap_16[7:0]),.cy( 9'sd1),.dx(input_fmap_24[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O2_N2_S1),.chainout(chainout_2_O2));
logic signed [63:0] chainout_4_O2; 
logic signed [63:0] O2_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O2(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_25[7:0]),.ay( 9'sd1),.bx(input_fmap_27[7:0]),.by( 9'sd1),.cx(input_fmap_30[7:0]),.cy(-9'sd2),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O2_N4_S1),.chainout(chainout_4_O2));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O2_N0_S2;		always @(posedge clk) O2_N0_S2 <=     O2_N0_S1  +  O2_N2_S1 ;
 logic signed [21:0] O2_N2_S2;		always @(posedge clk) O2_N2_S2 <=     O2_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O2_N0_S3;		always @(posedge clk) O2_N0_S3 <=     O2_N0_S2  +  O2_N2_S2 ;
 assign conv_mac_2 = O2_N0_S3;

logic signed [31:0] conv_mac_3;
logic signed [63:0] chainout_0_O3; 
logic signed [63:0] O3_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O3(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay(-9'sd1),.bx(input_fmap_5[7:0]),.by(-9'sd1),.cx(input_fmap_7[7:0]),.cy( 9'sd1),.dx(input_fmap_12[7:0]),.dy( 9'sd3),.chainin(63'd0),.result(O3_N0_S1),.chainout(chainout_0_O3));
logic signed [63:0] chainout_2_O3; 
logic signed [63:0] O3_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O3(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_13[7:0]),.ay(-9'sd2),.bx(input_fmap_15[7:0]),.by(-9'sd1),.cx(input_fmap_16[7:0]),.cy(-9'sd1),.dx(input_fmap_23[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O3_N2_S1),.chainout(chainout_2_O3));
logic signed [63:0] chainout_4_O3; 
logic signed [63:0] O3_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O3(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_25[7:0]),.ay(-9'sd1),.bx(input_fmap_26[7:0]),.by( 9'sd1),.cx(input_fmap_27[7:0]),.cy( 9'sd1),.dx(input_fmap_29[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O3_N4_S1),.chainout(chainout_4_O3));
logic signed [63:0] chainout_6_O3; 
logic signed [63:0] O3_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O3(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_30[7:0]),.ay( 9'sd2),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O3_N6_S1),.chainout(chainout_6_O3));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O3_N0_S2;		always @(posedge clk) O3_N0_S2 <=     O3_N0_S1  +  O3_N2_S1 ;
 logic signed [21:0] O3_N2_S2;		always @(posedge clk) O3_N2_S2 <=     O3_N4_S1  +  O3_N6_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O3_N0_S3;		always @(posedge clk) O3_N0_S3 <=     O3_N0_S2  +  O3_N2_S2 ;
 assign conv_mac_3 = O3_N0_S3;

logic signed [31:0] conv_mac_4;
logic signed [63:0] chainout_0_O4; 
logic signed [63:0] O4_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O4(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd2),.bx(input_fmap_1[7:0]),.by( 9'sd1),.cx(input_fmap_3[7:0]),.cy(-9'sd1),.dx(input_fmap_4[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O4_N0_S1),.chainout(chainout_0_O4));
logic signed [63:0] chainout_2_O4; 
logic signed [63:0] O4_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O4(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_6[7:0]),.ay( 9'sd1),.bx(input_fmap_8[7:0]),.by( 9'sd1),.cx(input_fmap_10[7:0]),.cy(-9'sd1),.dx(input_fmap_11[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O4_N2_S1),.chainout(chainout_2_O4));
logic signed [63:0] chainout_4_O4; 
logic signed [63:0] O4_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O4(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_15[7:0]),.ay( 9'sd1),.bx(input_fmap_16[7:0]),.by(-9'sd1),.cx(input_fmap_18[7:0]),.cy( 9'sd2),.dx(input_fmap_19[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O4_N4_S1),.chainout(chainout_4_O4));
logic signed [63:0] chainout_6_O4; 
logic signed [63:0] O4_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O4(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_20[7:0]),.ay( 9'sd2),.bx(input_fmap_21[7:0]),.by(-9'sd1),.cx(input_fmap_25[7:0]),.cy(-9'sd1),.dx(input_fmap_26[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O4_N6_S1),.chainout(chainout_6_O4));
logic signed [63:0] chainout_8_O4; 
logic signed [63:0] O4_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O4(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_28[7:0]),.ay(-9'sd1),.bx(input_fmap_29[7:0]),.by(-9'sd1),.cx(input_fmap_30[7:0]),.cy(-9'sd1),.dx(input_fmap_31[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O4_N8_S1),.chainout(chainout_8_O4));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O4_N0_S2;		always @(posedge clk) O4_N0_S2 <=     O4_N0_S1  +  O4_N2_S1 ;
 logic signed [21:0] O4_N2_S2;		always @(posedge clk) O4_N2_S2 <=     O4_N4_S1  +  O4_N6_S1 ;
 logic signed [21:0] O4_N4_S2;		always @(posedge clk) O4_N4_S2 <=     O4_N8_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O4_N0_S3;		always @(posedge clk) O4_N0_S3 <=     O4_N0_S2  +  O4_N2_S2 ;
 logic signed [22:0] O4_N2_S3;		always @(posedge clk) O4_N2_S3 <=     O4_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O4_N0_S4;		always @(posedge clk) O4_N0_S4 <=     O4_N0_S3  +  O4_N2_S3 ;
 assign conv_mac_4 = O4_N0_S4;

logic signed [31:0] conv_mac_5;
logic signed [63:0] chainout_0_O5; 
logic signed [63:0] O5_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O5(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_4[7:0]),.ay(-9'sd1),.bx(input_fmap_5[7:0]),.by( 9'sd1),.cx(input_fmap_6[7:0]),.cy( 9'sd1),.dx(input_fmap_9[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O5_N0_S1),.chainout(chainout_0_O5));
logic signed [63:0] chainout_2_O5; 
logic signed [63:0] O5_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O5(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_13[7:0]),.ay(-9'sd1),.bx(input_fmap_15[7:0]),.by( 9'sd1),.cx(input_fmap_21[7:0]),.cy( 9'sd1),.dx(input_fmap_22[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O5_N2_S1),.chainout(chainout_2_O5));
logic signed [63:0] chainout_4_O5; 
logic signed [63:0] O5_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O5(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_24[7:0]),.ay( 9'sd1),.bx(input_fmap_25[7:0]),.by(-9'sd1),.cx(input_fmap_30[7:0]),.cy( 9'sd1),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O5_N4_S1),.chainout(chainout_4_O5));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O5_N0_S2;		always @(posedge clk) O5_N0_S2 <=     O5_N0_S1  +  O5_N2_S1 ;
 logic signed [21:0] O5_N2_S2;		always @(posedge clk) O5_N2_S2 <=     O5_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O5_N0_S3;		always @(posedge clk) O5_N0_S3 <=     O5_N0_S2  +  O5_N2_S2 ;
 assign conv_mac_5 = O5_N0_S3;

logic signed [31:0] conv_mac_6;
logic signed [63:0] chainout_0_O6; 
logic signed [63:0] O6_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O6(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay(-9'sd1),.bx(input_fmap_3[7:0]),.by(-9'sd1),.cx(input_fmap_6[7:0]),.cy( 9'sd1),.dx(input_fmap_8[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O6_N0_S1),.chainout(chainout_0_O6));
logic signed [63:0] chainout_2_O6; 
logic signed [63:0] O6_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O6(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_11[7:0]),.ay(-9'sd2),.bx(input_fmap_13[7:0]),.by(-9'sd3),.cx(input_fmap_14[7:0]),.cy(-9'sd1),.dx(input_fmap_17[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O6_N2_S1),.chainout(chainout_2_O6));
logic signed [63:0] chainout_4_O6; 
logic signed [63:0] O6_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O6(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_18[7:0]),.ay(-9'sd1),.bx(input_fmap_19[7:0]),.by( 9'sd1),.cx(input_fmap_21[7:0]),.cy(-9'sd1),.dx(input_fmap_25[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O6_N4_S1),.chainout(chainout_4_O6));
logic signed [63:0] chainout_6_O6; 
logic signed [63:0] O6_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O6(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_27[7:0]),.ay(-9'sd1),.bx(input_fmap_28[7:0]),.by(-9'sd1),.cx(input_fmap_29[7:0]),.cy( 9'sd2),.dx(input_fmap_30[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O6_N6_S1),.chainout(chainout_6_O6));
logic signed [63:0] chainout_8_O6; 
logic signed [63:0] O6_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O6(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_31[7:0]),.ay( 9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O6_N8_S1),.chainout(chainout_8_O6));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O6_N0_S2;		always @(posedge clk) O6_N0_S2 <=     O6_N0_S1  +  O6_N2_S1 ;
 logic signed [21:0] O6_N2_S2;		always @(posedge clk) O6_N2_S2 <=     O6_N4_S1  +  O6_N6_S1 ;
 logic signed [21:0] O6_N4_S2;		always @(posedge clk) O6_N4_S2 <=     O6_N8_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O6_N0_S3;		always @(posedge clk) O6_N0_S3 <=     O6_N0_S2  +  O6_N2_S2 ;
 logic signed [22:0] O6_N2_S3;		always @(posedge clk) O6_N2_S3 <=     O6_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O6_N0_S4;		always @(posedge clk) O6_N0_S4 <=     O6_N0_S3  +  O6_N2_S3 ;
 assign conv_mac_6 = O6_N0_S4;

logic signed [31:0] conv_mac_7;
logic signed [63:0] chainout_0_O7; 
logic signed [63:0] O7_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O7(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_4[7:0]),.ay( 9'sd1),.bx(input_fmap_5[7:0]),.by( 9'sd1),.cx(input_fmap_8[7:0]),.cy( 9'sd1),.dx(input_fmap_10[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O7_N0_S1),.chainout(chainout_0_O7));
logic signed [63:0] chainout_2_O7; 
logic signed [63:0] O7_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O7(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_14[7:0]),.ay(-9'sd1),.bx(input_fmap_15[7:0]),.by(-9'sd1),.cx(input_fmap_26[7:0]),.cy( 9'sd1),.dx(input_fmap_28[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O7_N2_S1),.chainout(chainout_2_O7));
logic signed [63:0] chainout_4_O7; 
logic signed [63:0] O7_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O7(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_29[7:0]),.ay(-9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O7_N4_S1),.chainout(chainout_4_O7));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O7_N0_S2;		always @(posedge clk) O7_N0_S2 <=     O7_N0_S1  +  O7_N2_S1 ;
 logic signed [21:0] O7_N2_S2;		always @(posedge clk) O7_N2_S2 <=     O7_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O7_N0_S3;		always @(posedge clk) O7_N0_S3 <=     O7_N0_S2  +  O7_N2_S2 ;
 assign conv_mac_7 = O7_N0_S3;

logic signed [31:0] conv_mac_8;
logic signed [63:0] chainout_0_O8; 
logic signed [63:0] O8_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O8(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay(-9'sd1),.bx(input_fmap_2[7:0]),.by( 9'sd1),.cx(input_fmap_6[7:0]),.cy(-9'sd1),.dx(input_fmap_8[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O8_N0_S1),.chainout(chainout_0_O8));
logic signed [63:0] chainout_2_O8; 
logic signed [63:0] O8_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O8(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_11[7:0]),.ay(-9'sd1),.bx(input_fmap_12[7:0]),.by(-9'sd1),.cx(input_fmap_13[7:0]),.cy( 9'sd1),.dx(input_fmap_16[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O8_N2_S1),.chainout(chainout_2_O8));
logic signed [63:0] chainout_4_O8; 
logic signed [63:0] O8_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O8(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_17[7:0]),.ay(-9'sd1),.bx(input_fmap_21[7:0]),.by(-9'sd1),.cx(input_fmap_22[7:0]),.cy( 9'sd1),.dx(input_fmap_23[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O8_N4_S1),.chainout(chainout_4_O8));
logic signed [63:0] chainout_6_O8; 
logic signed [63:0] O8_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O8(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_26[7:0]),.ay(-9'sd1),.bx(input_fmap_30[7:0]),.by(-9'sd2),.cx(input_fmap_31[7:0]),.cy(-9'sd2),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O8_N6_S1),.chainout(chainout_6_O8));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O8_N0_S2;		always @(posedge clk) O8_N0_S2 <=     O8_N0_S1  +  O8_N2_S1 ;
 logic signed [21:0] O8_N2_S2;		always @(posedge clk) O8_N2_S2 <=     O8_N4_S1  +  O8_N6_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O8_N0_S3;		always @(posedge clk) O8_N0_S3 <=     O8_N0_S2  +  O8_N2_S2 ;
 assign conv_mac_8 = O8_N0_S3;

logic signed [31:0] conv_mac_9;
logic signed [63:0] chainout_0_O9; 
logic signed [63:0] O9_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O9(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd1),.bx(input_fmap_4[7:0]),.by( 9'sd1),.cx(input_fmap_5[7:0]),.cy( 9'sd1),.dx(input_fmap_7[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O9_N0_S1),.chainout(chainout_0_O9));
logic signed [63:0] chainout_2_O9; 
logic signed [63:0] O9_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O9(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_8[7:0]),.ay( 9'sd1),.bx(input_fmap_10[7:0]),.by( 9'sd2),.cx(input_fmap_11[7:0]),.cy( 9'sd1),.dx(input_fmap_14[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O9_N2_S1),.chainout(chainout_2_O9));
logic signed [63:0] chainout_4_O9; 
logic signed [63:0] O9_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O9(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_15[7:0]),.ay(-9'sd2),.bx(input_fmap_16[7:0]),.by( 9'sd1),.cx(input_fmap_22[7:0]),.cy(-9'sd1),.dx(input_fmap_23[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O9_N4_S1),.chainout(chainout_4_O9));
logic signed [63:0] chainout_6_O9; 
logic signed [63:0] O9_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O9(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_24[7:0]),.ay(-9'sd1),.bx(input_fmap_26[7:0]),.by( 9'sd1),.cx(input_fmap_28[7:0]),.cy(-9'sd1),.dx(input_fmap_29[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O9_N6_S1),.chainout(chainout_6_O9));
logic signed [63:0] chainout_8_O9; 
logic signed [63:0] O9_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O9(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_30[7:0]),.ay( 9'sd1),.bx(input_fmap_31[7:0]),.by( 9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O9_N8_S1),.chainout(chainout_8_O9));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O9_N0_S2;		always @(posedge clk) O9_N0_S2 <=     O9_N0_S1  +  O9_N2_S1 ;
 logic signed [21:0] O9_N2_S2;		always @(posedge clk) O9_N2_S2 <=     O9_N4_S1  +  O9_N6_S1 ;
 logic signed [21:0] O9_N4_S2;		always @(posedge clk) O9_N4_S2 <=     O9_N8_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O9_N0_S3;		always @(posedge clk) O9_N0_S3 <=     O9_N0_S2  +  O9_N2_S2 ;
 logic signed [22:0] O9_N2_S3;		always @(posedge clk) O9_N2_S3 <=     O9_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O9_N0_S4;		always @(posedge clk) O9_N0_S4 <=     O9_N0_S3  +  O9_N2_S3 ;
 assign conv_mac_9 = O9_N0_S4;

logic signed [31:0] conv_mac_10;
logic signed [63:0] chainout_0_O10; 
logic signed [63:0] O10_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O10(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay(-9'sd1),.bx(input_fmap_2[7:0]),.by( 9'sd1),.cx(input_fmap_7[7:0]),.cy( 9'sd1),.dx(input_fmap_10[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O10_N0_S1),.chainout(chainout_0_O10));
logic signed [63:0] chainout_2_O10; 
logic signed [63:0] O10_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O10(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_12[7:0]),.ay(-9'sd1),.bx(input_fmap_13[7:0]),.by(-9'sd1),.cx(input_fmap_15[7:0]),.cy( 9'sd2),.dx(input_fmap_17[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O10_N2_S1),.chainout(chainout_2_O10));
logic signed [63:0] chainout_4_O10; 
logic signed [63:0] O10_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O10(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_18[7:0]),.ay(-9'sd2),.bx(input_fmap_19[7:0]),.by( 9'sd1),.cx(input_fmap_21[7:0]),.cy( 9'sd2),.dx(input_fmap_25[7:0]),.dy( 9'sd5),.chainin(63'd0),.result(O10_N4_S1),.chainout(chainout_4_O10));
logic signed [63:0] chainout_6_O10; 
logic signed [63:0] O10_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O10(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_26[7:0]),.ay(-9'sd1),.bx(input_fmap_28[7:0]),.by(-9'sd1),.cx(input_fmap_29[7:0]),.cy( 9'sd4),.dx(input_fmap_30[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O10_N6_S1),.chainout(chainout_6_O10));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O10_N0_S2;		always @(posedge clk) O10_N0_S2 <=     O10_N0_S1  +  O10_N2_S1 ;
 logic signed [21:0] O10_N2_S2;		always @(posedge clk) O10_N2_S2 <=     O10_N4_S1  +  O10_N6_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O10_N0_S3;		always @(posedge clk) O10_N0_S3 <=     O10_N0_S2  +  O10_N2_S2 ;
 assign conv_mac_10 = O10_N0_S3;

logic signed [31:0] conv_mac_11;
logic signed [63:0] chainout_0_O11; 
logic signed [63:0] O11_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O11(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd1),.bx(input_fmap_1[7:0]),.by( 9'sd2),.cx(input_fmap_5[7:0]),.cy( 9'sd2),.dx(input_fmap_6[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O11_N0_S1),.chainout(chainout_0_O11));
logic signed [63:0] chainout_2_O11; 
logic signed [63:0] O11_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O11(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_8[7:0]),.ay(-9'sd1),.bx(input_fmap_10[7:0]),.by( 9'sd1),.cx(input_fmap_13[7:0]),.cy( 9'sd1),.dx(input_fmap_14[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O11_N2_S1),.chainout(chainout_2_O11));
logic signed [63:0] chainout_4_O11; 
logic signed [63:0] O11_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O11(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_15[7:0]),.ay( 9'sd1),.bx(input_fmap_19[7:0]),.by(-9'sd1),.cx(input_fmap_20[7:0]),.cy( 9'sd1),.dx(input_fmap_21[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O11_N4_S1),.chainout(chainout_4_O11));
logic signed [63:0] chainout_6_O11; 
logic signed [63:0] O11_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O11(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_24[7:0]),.ay( 9'sd1),.bx(input_fmap_30[7:0]),.by( 9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O11_N6_S1),.chainout(chainout_6_O11));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O11_N0_S2;		always @(posedge clk) O11_N0_S2 <=     O11_N0_S1  +  O11_N2_S1 ;
 logic signed [21:0] O11_N2_S2;		always @(posedge clk) O11_N2_S2 <=     O11_N4_S1  +  O11_N6_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O11_N0_S3;		always @(posedge clk) O11_N0_S3 <=     O11_N0_S2  +  O11_N2_S2 ;
 assign conv_mac_11 = O11_N0_S3;

logic signed [31:0] conv_mac_12;
logic signed [63:0] chainout_0_O12; 
logic signed [63:0] O12_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O12(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay( 9'sd2),.bx(input_fmap_2[7:0]),.by( 9'sd2),.cx(input_fmap_8[7:0]),.cy( 9'sd1),.dx(input_fmap_9[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O12_N0_S1),.chainout(chainout_0_O12));
logic signed [63:0] chainout_2_O12; 
logic signed [63:0] O12_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O12(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_11[7:0]),.ay( 9'sd1),.bx(input_fmap_13[7:0]),.by( 9'sd2),.cx(input_fmap_16[7:0]),.cy( 9'sd1),.dx(input_fmap_17[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O12_N2_S1),.chainout(chainout_2_O12));
logic signed [63:0] chainout_4_O12; 
logic signed [63:0] O12_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O12(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_20[7:0]),.ay(-9'sd1),.bx(input_fmap_23[7:0]),.by( 9'sd1),.cx(input_fmap_29[7:0]),.cy(-9'sd1),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O12_N4_S1),.chainout(chainout_4_O12));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O12_N0_S2;		always @(posedge clk) O12_N0_S2 <=     O12_N0_S1  +  O12_N2_S1 ;
 logic signed [21:0] O12_N2_S2;		always @(posedge clk) O12_N2_S2 <=     O12_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O12_N0_S3;		always @(posedge clk) O12_N0_S3 <=     O12_N0_S2  +  O12_N2_S2 ;
 assign conv_mac_12 = O12_N0_S3;

logic signed [31:0] conv_mac_13;
logic signed [63:0] chainout_0_O13; 
logic signed [63:0] O13_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O13(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd2),.bx(input_fmap_1[7:0]),.by( 9'sd1),.cx(input_fmap_2[7:0]),.cy( 9'sd1),.dx(input_fmap_3[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O13_N0_S1),.chainout(chainout_0_O13));
logic signed [63:0] chainout_2_O13; 
logic signed [63:0] O13_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O13(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_4[7:0]),.ay(-9'sd1),.bx(input_fmap_7[7:0]),.by( 9'sd1),.cx(input_fmap_8[7:0]),.cy(-9'sd1),.dx(input_fmap_14[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O13_N2_S1),.chainout(chainout_2_O13));
logic signed [63:0] chainout_4_O13; 
logic signed [63:0] O13_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O13(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_16[7:0]),.ay(-9'sd2),.bx(input_fmap_19[7:0]),.by(-9'sd1),.cx(input_fmap_20[7:0]),.cy(-9'sd1),.dx(input_fmap_21[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O13_N4_S1),.chainout(chainout_4_O13));
logic signed [63:0] chainout_6_O13; 
logic signed [63:0] O13_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O13(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_22[7:0]),.ay( 9'sd1),.bx(input_fmap_24[7:0]),.by( 9'sd1),.cx(input_fmap_25[7:0]),.cy(-9'sd1),.dx(input_fmap_26[7:0]),.dy( 9'sd3),.chainin(63'd0),.result(O13_N6_S1),.chainout(chainout_6_O13));
logic signed [63:0] chainout_8_O13; 
logic signed [63:0] O13_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O13(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_27[7:0]),.ay(-9'sd2),.bx(input_fmap_28[7:0]),.by( 9'sd1),.cx(input_fmap_29[7:0]),.cy( 9'sd2),.dx(input_fmap_30[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O13_N8_S1),.chainout(chainout_8_O13));
logic signed [63:0] chainout_10_O13; 
logic signed [63:0] O13_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O13(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_31[7:0]),.ay(-9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O13_N10_S1),.chainout(chainout_10_O13));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O13_N0_S2;		always @(posedge clk) O13_N0_S2 <=     O13_N0_S1  +  O13_N2_S1 ;
 logic signed [21:0] O13_N2_S2;		always @(posedge clk) O13_N2_S2 <=     O13_N4_S1  +  O13_N6_S1 ;
 logic signed [21:0] O13_N4_S2;		always @(posedge clk) O13_N4_S2 <=     O13_N8_S1  +  O13_N10_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O13_N0_S3;		always @(posedge clk) O13_N0_S3 <=     O13_N0_S2  +  O13_N2_S2 ;
 logic signed [22:0] O13_N2_S3;		always @(posedge clk) O13_N2_S3 <=     O13_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O13_N0_S4;		always @(posedge clk) O13_N0_S4 <=     O13_N0_S3  +  O13_N2_S3 ;
 assign conv_mac_13 = O13_N0_S4;

logic signed [31:0] conv_mac_14;
logic signed [63:0] chainout_0_O14; 
logic signed [63:0] O14_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O14(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd2),.bx(input_fmap_2[7:0]),.by( 9'sd3),.cx(input_fmap_3[7:0]),.cy( 9'sd1),.dx(input_fmap_4[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O14_N0_S1),.chainout(chainout_0_O14));
logic signed [63:0] chainout_2_O14; 
logic signed [63:0] O14_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O14(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_5[7:0]),.ay(-9'sd1),.bx(input_fmap_7[7:0]),.by(-9'sd2),.cx(input_fmap_11[7:0]),.cy(-9'sd1),.dx(input_fmap_12[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O14_N2_S1),.chainout(chainout_2_O14));
logic signed [63:0] chainout_4_O14; 
logic signed [63:0] O14_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O14(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_13[7:0]),.ay(-9'sd3),.bx(input_fmap_15[7:0]),.by(-9'sd1),.cx(input_fmap_16[7:0]),.cy( 9'sd3),.dx(input_fmap_21[7:0]),.dy( 9'sd4),.chainin(63'd0),.result(O14_N4_S1),.chainout(chainout_4_O14));
logic signed [63:0] chainout_6_O14; 
logic signed [63:0] O14_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O14(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_22[7:0]),.ay( 9'sd2),.bx(input_fmap_23[7:0]),.by( 9'sd1),.cx(input_fmap_26[7:0]),.cy( 9'sd1),.dx(input_fmap_28[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O14_N6_S1),.chainout(chainout_6_O14));
logic signed [63:0] chainout_8_O14; 
logic signed [63:0] O14_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O14(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_29[7:0]),.ay(-9'sd1),.bx(input_fmap_31[7:0]),.by(-9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O14_N8_S1),.chainout(chainout_8_O14));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O14_N0_S2;		always @(posedge clk) O14_N0_S2 <=     O14_N0_S1  +  O14_N2_S1 ;
 logic signed [21:0] O14_N2_S2;		always @(posedge clk) O14_N2_S2 <=     O14_N4_S1  +  O14_N6_S1 ;
 logic signed [21:0] O14_N4_S2;		always @(posedge clk) O14_N4_S2 <=     O14_N8_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O14_N0_S3;		always @(posedge clk) O14_N0_S3 <=     O14_N0_S2  +  O14_N2_S2 ;
 logic signed [22:0] O14_N2_S3;		always @(posedge clk) O14_N2_S3 <=     O14_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O14_N0_S4;		always @(posedge clk) O14_N0_S4 <=     O14_N0_S3  +  O14_N2_S3 ;
 assign conv_mac_14 = O14_N0_S4;

logic signed [31:0] conv_mac_15;
logic signed [63:0] chainout_0_O15; 
logic signed [63:0] O15_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O15(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd1),.bx(input_fmap_1[7:0]),.by(-9'sd1),.cx(input_fmap_3[7:0]),.cy( 9'sd4),.dx(input_fmap_4[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O15_N0_S1),.chainout(chainout_0_O15));
logic signed [63:0] chainout_2_O15; 
logic signed [63:0] O15_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O15(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_5[7:0]),.ay( 9'sd1),.bx(input_fmap_6[7:0]),.by( 9'sd2),.cx(input_fmap_8[7:0]),.cy( 9'sd2),.dx(input_fmap_16[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O15_N2_S1),.chainout(chainout_2_O15));
logic signed [63:0] chainout_4_O15; 
logic signed [63:0] O15_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O15(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_17[7:0]),.ay( 9'sd1),.bx(input_fmap_18[7:0]),.by( 9'sd1),.cx(input_fmap_21[7:0]),.cy( 9'sd2),.dx(input_fmap_22[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O15_N4_S1),.chainout(chainout_4_O15));
logic signed [63:0] chainout_6_O15; 
logic signed [63:0] O15_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O15(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_25[7:0]),.ay(-9'sd1),.bx(input_fmap_27[7:0]),.by( 9'sd1),.cx(input_fmap_28[7:0]),.cy(-9'sd1),.dx(input_fmap_31[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O15_N6_S1),.chainout(chainout_6_O15));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O15_N0_S2;		always @(posedge clk) O15_N0_S2 <=     O15_N0_S1  +  O15_N2_S1 ;
 logic signed [21:0] O15_N2_S2;		always @(posedge clk) O15_N2_S2 <=     O15_N4_S1  +  O15_N6_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O15_N0_S3;		always @(posedge clk) O15_N0_S3 <=     O15_N0_S2  +  O15_N2_S2 ;
 assign conv_mac_15 = O15_N0_S3;

logic signed [31:0] conv_mac_16;
logic signed [63:0] chainout_0_O16; 
logic signed [63:0] O16_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O16(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay( 9'sd1),.bx(input_fmap_2[7:0]),.by(-9'sd1),.cx(input_fmap_6[7:0]),.cy(-9'sd1),.dx(input_fmap_14[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O16_N0_S1),.chainout(chainout_0_O16));
logic signed [63:0] chainout_2_O16; 
logic signed [63:0] O16_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O16(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_17[7:0]),.ay( 9'sd2),.bx(input_fmap_18[7:0]),.by( 9'sd1),.cx(input_fmap_22[7:0]),.cy(-9'sd1),.dx(input_fmap_23[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O16_N2_S1),.chainout(chainout_2_O16));
logic signed [63:0] chainout_4_O16; 
logic signed [63:0] O16_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O16(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_27[7:0]),.ay( 9'sd2),.bx(input_fmap_29[7:0]),.by(-9'sd1),.cx(input_fmap_30[7:0]),.cy( 9'sd1),.dx(input_fmap_31[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O16_N4_S1),.chainout(chainout_4_O16));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O16_N0_S2;		always @(posedge clk) O16_N0_S2 <=     O16_N0_S1  +  O16_N2_S1 ;
 logic signed [21:0] O16_N2_S2;		always @(posedge clk) O16_N2_S2 <=     O16_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O16_N0_S3;		always @(posedge clk) O16_N0_S3 <=     O16_N0_S2  +  O16_N2_S2 ;
 assign conv_mac_16 = O16_N0_S3;

logic signed [31:0] conv_mac_17;
logic signed [63:0] chainout_0_O17; 
logic signed [63:0] O17_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O17(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_9[7:0]),.ay( 9'sd1),.bx(input_fmap_10[7:0]),.by(-9'sd1),.cx(input_fmap_17[7:0]),.cy(-9'sd1),.dx(input_fmap_24[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O17_N0_S1),.chainout(chainout_0_O17));
logic signed [63:0] chainout_2_O17; 
logic signed [63:0] O17_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O17(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_31[7:0]),.ay( 9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O17_N2_S1),.chainout(chainout_2_O17));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O17_N0_S2;		always @(posedge clk) O17_N0_S2 <=     O17_N0_S1  +  O17_N2_S1 ;
 assign conv_mac_17 = O17_N0_S2;

logic signed [31:0] conv_mac_18;
logic signed [63:0] chainout_0_O18; 
logic signed [63:0] O18_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O18(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd1),.bx(input_fmap_1[7:0]),.by( 9'sd1),.cx(input_fmap_2[7:0]),.cy(-9'sd1),.dx(input_fmap_3[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O18_N0_S1),.chainout(chainout_0_O18));
logic signed [63:0] chainout_2_O18; 
logic signed [63:0] O18_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O18(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_5[7:0]),.ay(-9'sd1),.bx(input_fmap_6[7:0]),.by(-9'sd2),.cx(input_fmap_10[7:0]),.cy(-9'sd1),.dx(input_fmap_11[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O18_N2_S1),.chainout(chainout_2_O18));
logic signed [63:0] chainout_4_O18; 
logic signed [63:0] O18_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O18(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_12[7:0]),.ay( 9'sd1),.bx(input_fmap_13[7:0]),.by(-9'sd1),.cx(input_fmap_14[7:0]),.cy( 9'sd1),.dx(input_fmap_15[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O18_N4_S1),.chainout(chainout_4_O18));
logic signed [63:0] chainout_6_O18; 
logic signed [63:0] O18_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O18(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_17[7:0]),.ay( 9'sd1),.bx(input_fmap_20[7:0]),.by(-9'sd1),.cx(input_fmap_21[7:0]),.cy( 9'sd1),.dx(input_fmap_22[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O18_N6_S1),.chainout(chainout_6_O18));
logic signed [63:0] chainout_8_O18; 
logic signed [63:0] O18_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O18(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_23[7:0]),.ay(-9'sd1),.bx(input_fmap_25[7:0]),.by( 9'sd1),.cx(input_fmap_26[7:0]),.cy( 9'sd1),.dx(input_fmap_27[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O18_N8_S1),.chainout(chainout_8_O18));
logic signed [63:0] chainout_10_O18; 
logic signed [63:0] O18_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O18(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_29[7:0]),.ay(-9'sd1),.bx(input_fmap_30[7:0]),.by(-9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O18_N10_S1),.chainout(chainout_10_O18));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O18_N0_S2;		always @(posedge clk) O18_N0_S2 <=     O18_N0_S1  +  O18_N2_S1 ;
 logic signed [21:0] O18_N2_S2;		always @(posedge clk) O18_N2_S2 <=     O18_N4_S1  +  O18_N6_S1 ;
 logic signed [21:0] O18_N4_S2;		always @(posedge clk) O18_N4_S2 <=     O18_N8_S1  +  O18_N10_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O18_N0_S3;		always @(posedge clk) O18_N0_S3 <=     O18_N0_S2  +  O18_N2_S2 ;
 logic signed [22:0] O18_N2_S3;		always @(posedge clk) O18_N2_S3 <=     O18_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O18_N0_S4;		always @(posedge clk) O18_N0_S4 <=     O18_N0_S3  +  O18_N2_S3 ;
 assign conv_mac_18 = O18_N0_S4;

logic signed [31:0] conv_mac_19;
logic signed [63:0] chainout_0_O19; 
logic signed [63:0] O19_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O19(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd1),.bx(input_fmap_1[7:0]),.by( 9'sd1),.cx(input_fmap_4[7:0]),.cy( 9'sd1),.dx(input_fmap_8[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O19_N0_S1),.chainout(chainout_0_O19));
logic signed [63:0] chainout_2_O19; 
logic signed [63:0] O19_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O19(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_12[7:0]),.ay( 9'sd1),.bx(input_fmap_14[7:0]),.by(-9'sd1),.cx(input_fmap_15[7:0]),.cy( 9'sd1),.dx(input_fmap_16[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O19_N2_S1),.chainout(chainout_2_O19));
logic signed [63:0] chainout_4_O19; 
logic signed [63:0] O19_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O19(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_17[7:0]),.ay(-9'sd1),.bx(input_fmap_19[7:0]),.by(-9'sd1),.cx(input_fmap_24[7:0]),.cy(-9'sd1),.dx(input_fmap_26[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O19_N4_S1),.chainout(chainout_4_O19));
logic signed [63:0] chainout_6_O19; 
logic signed [63:0] O19_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O19(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_27[7:0]),.ay( 9'sd3),.bx(input_fmap_31[7:0]),.by(-9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O19_N6_S1),.chainout(chainout_6_O19));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O19_N0_S2;		always @(posedge clk) O19_N0_S2 <=     O19_N0_S1  +  O19_N2_S1 ;
 logic signed [21:0] O19_N2_S2;		always @(posedge clk) O19_N2_S2 <=     O19_N4_S1  +  O19_N6_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O19_N0_S3;		always @(posedge clk) O19_N0_S3 <=     O19_N0_S2  +  O19_N2_S2 ;
 assign conv_mac_19 = O19_N0_S3;

logic signed [31:0] conv_mac_20;
logic signed [63:0] chainout_0_O20; 
logic signed [63:0] O20_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O20(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay(-9'sd1),.bx(input_fmap_2[7:0]),.by( 9'sd4),.cx(input_fmap_3[7:0]),.cy(-9'sd1),.dx(input_fmap_6[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O20_N0_S1),.chainout(chainout_0_O20));
logic signed [63:0] chainout_2_O20; 
logic signed [63:0] O20_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O20(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_9[7:0]),.ay( 9'sd1),.bx(input_fmap_11[7:0]),.by(-9'sd1),.cx(input_fmap_16[7:0]),.cy( 9'sd3),.dx(input_fmap_23[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O20_N2_S1),.chainout(chainout_2_O20));
logic signed [63:0] chainout_4_O20; 
logic signed [63:0] O20_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O20(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_25[7:0]),.ay( 9'sd1),.bx(input_fmap_26[7:0]),.by( 9'sd1),.cx(input_fmap_27[7:0]),.cy(-9'sd1),.dx(input_fmap_30[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O20_N4_S1),.chainout(chainout_4_O20));
logic signed [63:0] chainout_6_O20; 
logic signed [63:0] O20_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O20(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_31[7:0]),.ay(-9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O20_N6_S1),.chainout(chainout_6_O20));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O20_N0_S2;		always @(posedge clk) O20_N0_S2 <=     O20_N0_S1  +  O20_N2_S1 ;
 logic signed [21:0] O20_N2_S2;		always @(posedge clk) O20_N2_S2 <=     O20_N4_S1  +  O20_N6_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O20_N0_S3;		always @(posedge clk) O20_N0_S3 <=     O20_N0_S2  +  O20_N2_S2 ;
 assign conv_mac_20 = O20_N0_S3;

logic signed [31:0] conv_mac_21;
logic signed [63:0] chainout_0_O21; 
logic signed [63:0] O21_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O21(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_2[7:0]),.ay(-9'sd1),.bx(input_fmap_3[7:0]),.by(-9'sd1),.cx(input_fmap_5[7:0]),.cy(-9'sd2),.dx(input_fmap_6[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O21_N0_S1),.chainout(chainout_0_O21));
logic signed [63:0] chainout_2_O21; 
logic signed [63:0] O21_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O21(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_10[7:0]),.ay(-9'sd2),.bx(input_fmap_11[7:0]),.by(-9'sd1),.cx(input_fmap_13[7:0]),.cy(-9'sd2),.dx(input_fmap_14[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O21_N2_S1),.chainout(chainout_2_O21));
logic signed [63:0] chainout_4_O21; 
logic signed [63:0] O21_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O21(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_15[7:0]),.ay(-9'sd1),.bx(input_fmap_17[7:0]),.by(-9'sd1),.cx(input_fmap_18[7:0]),.cy(-9'sd1),.dx(input_fmap_19[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O21_N4_S1),.chainout(chainout_4_O21));
logic signed [63:0] chainout_6_O21; 
logic signed [63:0] O21_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O21(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_20[7:0]),.ay(-9'sd1),.bx(input_fmap_21[7:0]),.by(-9'sd1),.cx(input_fmap_23[7:0]),.cy(-9'sd1),.dx(input_fmap_24[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O21_N6_S1),.chainout(chainout_6_O21));
logic signed [63:0] chainout_8_O21; 
logic signed [63:0] O21_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O21(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_25[7:0]),.ay( 9'sd2),.bx(input_fmap_26[7:0]),.by(-9'sd1),.cx(input_fmap_27[7:0]),.cy( 9'sd1),.dx(input_fmap_28[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O21_N8_S1),.chainout(chainout_8_O21));
logic signed [63:0] chainout_10_O21; 
logic signed [63:0] O21_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O21(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_30[7:0]),.ay( 9'sd1),.bx(input_fmap_31[7:0]),.by( 9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O21_N10_S1),.chainout(chainout_10_O21));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O21_N0_S2;		always @(posedge clk) O21_N0_S2 <=     O21_N0_S1  +  O21_N2_S1 ;
 logic signed [21:0] O21_N2_S2;		always @(posedge clk) O21_N2_S2 <=     O21_N4_S1  +  O21_N6_S1 ;
 logic signed [21:0] O21_N4_S2;		always @(posedge clk) O21_N4_S2 <=     O21_N8_S1  +  O21_N10_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O21_N0_S3;		always @(posedge clk) O21_N0_S3 <=     O21_N0_S2  +  O21_N2_S2 ;
 logic signed [22:0] O21_N2_S3;		always @(posedge clk) O21_N2_S3 <=     O21_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O21_N0_S4;		always @(posedge clk) O21_N0_S4 <=     O21_N0_S3  +  O21_N2_S3 ;
 assign conv_mac_21 = O21_N0_S4;

logic signed [31:0] conv_mac_22;
logic signed [63:0] chainout_0_O22; 
logic signed [63:0] O22_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O22(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay( 9'sd1),.bx(input_fmap_2[7:0]),.by(-9'sd2),.cx(input_fmap_3[7:0]),.cy( 9'sd1),.dx(input_fmap_4[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O22_N0_S1),.chainout(chainout_0_O22));
logic signed [63:0] chainout_2_O22; 
logic signed [63:0] O22_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O22(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_6[7:0]),.ay(-9'sd1),.bx(input_fmap_7[7:0]),.by(-9'sd1),.cx(input_fmap_8[7:0]),.cy(-9'sd1),.dx(input_fmap_9[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O22_N2_S1),.chainout(chainout_2_O22));
logic signed [63:0] chainout_4_O22; 
logic signed [63:0] O22_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O22(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_10[7:0]),.ay( 9'sd1),.bx(input_fmap_12[7:0]),.by(-9'sd1),.cx(input_fmap_13[7:0]),.cy(-9'sd2),.dx(input_fmap_16[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O22_N4_S1),.chainout(chainout_4_O22));
logic signed [63:0] chainout_6_O22; 
logic signed [63:0] O22_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O22(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_17[7:0]),.ay( 9'sd1),.bx(input_fmap_18[7:0]),.by(-9'sd1),.cx(input_fmap_21[7:0]),.cy(-9'sd1),.dx(input_fmap_22[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O22_N6_S1),.chainout(chainout_6_O22));
logic signed [63:0] chainout_8_O22; 
logic signed [63:0] O22_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O22(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_23[7:0]),.ay(-9'sd1),.bx(input_fmap_25[7:0]),.by( 9'sd1),.cx(input_fmap_26[7:0]),.cy(-9'sd1),.dx(input_fmap_27[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O22_N8_S1),.chainout(chainout_8_O22));
logic signed [63:0] chainout_10_O22; 
logic signed [63:0] O22_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O22(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_30[7:0]),.ay( 9'sd2),.bx(input_fmap_31[7:0]),.by( 9'sd2),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O22_N10_S1),.chainout(chainout_10_O22));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O22_N0_S2;		always @(posedge clk) O22_N0_S2 <=     O22_N0_S1  +  O22_N2_S1 ;
 logic signed [21:0] O22_N2_S2;		always @(posedge clk) O22_N2_S2 <=     O22_N4_S1  +  O22_N6_S1 ;
 logic signed [21:0] O22_N4_S2;		always @(posedge clk) O22_N4_S2 <=     O22_N8_S1  +  O22_N10_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O22_N0_S3;		always @(posedge clk) O22_N0_S3 <=     O22_N0_S2  +  O22_N2_S2 ;
 logic signed [22:0] O22_N2_S3;		always @(posedge clk) O22_N2_S3 <=     O22_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O22_N0_S4;		always @(posedge clk) O22_N0_S4 <=     O22_N0_S3  +  O22_N2_S3 ;
 assign conv_mac_22 = O22_N0_S4;

logic signed [31:0] conv_mac_23;
logic signed [63:0] chainout_0_O23; 
logic signed [63:0] O23_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O23(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd1),.bx(input_fmap_2[7:0]),.by( 9'sd1),.cx(input_fmap_7[7:0]),.cy( 9'sd1),.dx(input_fmap_10[7:0]),.dy( 9'sd3),.chainin(63'd0),.result(O23_N0_S1),.chainout(chainout_0_O23));
logic signed [63:0] chainout_2_O23; 
logic signed [63:0] O23_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O23(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_11[7:0]),.ay(-9'sd1),.bx(input_fmap_14[7:0]),.by(-9'sd1),.cx(input_fmap_16[7:0]),.cy( 9'sd1),.dx(input_fmap_17[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O23_N2_S1),.chainout(chainout_2_O23));
logic signed [63:0] chainout_4_O23; 
logic signed [63:0] O23_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O23(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_18[7:0]),.ay( 9'sd1),.bx(input_fmap_20[7:0]),.by(-9'sd1),.cx(input_fmap_21[7:0]),.cy( 9'sd1),.dx(input_fmap_24[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O23_N4_S1),.chainout(chainout_4_O23));
logic signed [63:0] chainout_6_O23; 
logic signed [63:0] O23_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O23(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_25[7:0]),.ay( 9'sd1),.bx(input_fmap_27[7:0]),.by( 9'sd1),.cx(input_fmap_28[7:0]),.cy( 9'sd1),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O23_N6_S1),.chainout(chainout_6_O23));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O23_N0_S2;		always @(posedge clk) O23_N0_S2 <=     O23_N0_S1  +  O23_N2_S1 ;
 logic signed [21:0] O23_N2_S2;		always @(posedge clk) O23_N2_S2 <=     O23_N4_S1  +  O23_N6_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O23_N0_S3;		always @(posedge clk) O23_N0_S3 <=     O23_N0_S2  +  O23_N2_S2 ;
 assign conv_mac_23 = O23_N0_S3;

logic signed [31:0] conv_mac_24;
logic signed [63:0] chainout_0_O24; 
logic signed [63:0] O24_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O24(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay(-9'sd1),.bx(input_fmap_2[7:0]),.by( 9'sd2),.cx(input_fmap_3[7:0]),.cy( 9'sd1),.dx(input_fmap_7[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O24_N0_S1),.chainout(chainout_0_O24));
logic signed [63:0] chainout_2_O24; 
logic signed [63:0] O24_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O24(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_10[7:0]),.ay(-9'sd1),.bx(input_fmap_16[7:0]),.by(-9'sd1),.cx(input_fmap_20[7:0]),.cy(-9'sd1),.dx(input_fmap_22[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O24_N2_S1),.chainout(chainout_2_O24));
logic signed [63:0] chainout_4_O24; 
logic signed [63:0] O24_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O24(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_23[7:0]),.ay( 9'sd3),.bx(input_fmap_26[7:0]),.by(-9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O24_N4_S1),.chainout(chainout_4_O24));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O24_N0_S2;		always @(posedge clk) O24_N0_S2 <=     O24_N0_S1  +  O24_N2_S1 ;
 logic signed [21:0] O24_N2_S2;		always @(posedge clk) O24_N2_S2 <=     O24_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O24_N0_S3;		always @(posedge clk) O24_N0_S3 <=     O24_N0_S2  +  O24_N2_S2 ;
 assign conv_mac_24 = O24_N0_S3;

logic signed [31:0] conv_mac_25;
logic signed [63:0] chainout_0_O25; 
logic signed [63:0] O25_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O25(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_2[7:0]),.ay(-9'sd2),.bx(input_fmap_7[7:0]),.by( 9'sd2),.cx(input_fmap_22[7:0]),.cy(-9'sd1),.dx(input_fmap_23[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O25_N0_S1),.chainout(chainout_0_O25));
assign conv_mac_25 = O25_N0_S1;

logic signed [31:0] conv_mac_26;
logic signed [63:0] chainout_0_O26; 
logic signed [63:0] O26_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O26(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay( 9'sd1),.bx(input_fmap_7[7:0]),.by(-9'sd1),.cx(input_fmap_9[7:0]),.cy( 9'sd1),.dx(input_fmap_13[7:0]),.dy( 9'sd3),.chainin(63'd0),.result(O26_N0_S1),.chainout(chainout_0_O26));
logic signed [63:0] chainout_2_O26; 
logic signed [63:0] O26_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O26(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_19[7:0]),.ay( 9'sd1),.bx(input_fmap_22[7:0]),.by( 9'sd1),.cx(input_fmap_23[7:0]),.cy(-9'sd1),.dx(input_fmap_25[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O26_N2_S1),.chainout(chainout_2_O26));
logic signed [63:0] chainout_4_O26; 
logic signed [63:0] O26_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O26(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_30[7:0]),.ay(-9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O26_N4_S1),.chainout(chainout_4_O26));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O26_N0_S2;		always @(posedge clk) O26_N0_S2 <=     O26_N0_S1  +  O26_N2_S1 ;
 logic signed [21:0] O26_N2_S2;		always @(posedge clk) O26_N2_S2 <=     O26_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O26_N0_S3;		always @(posedge clk) O26_N0_S3 <=     O26_N0_S2  +  O26_N2_S2 ;
 assign conv_mac_26 = O26_N0_S3;

logic signed [31:0] conv_mac_27;
logic signed [63:0] chainout_0_O27; 
logic signed [63:0] O27_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O27(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_3[7:0]),.ay( 9'sd1),.bx(input_fmap_4[7:0]),.by( 9'sd1),.cx(input_fmap_5[7:0]),.cy( 9'sd1),.dx(input_fmap_6[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O27_N0_S1),.chainout(chainout_0_O27));
logic signed [63:0] chainout_2_O27; 
logic signed [63:0] O27_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O27(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_7[7:0]),.ay(-9'sd1),.bx(input_fmap_8[7:0]),.by( 9'sd1),.cx(input_fmap_9[7:0]),.cy( 9'sd1),.dx(input_fmap_11[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O27_N2_S1),.chainout(chainout_2_O27));
logic signed [63:0] chainout_4_O27; 
logic signed [63:0] O27_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O27(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_14[7:0]),.ay( 9'sd1),.bx(input_fmap_17[7:0]),.by( 9'sd1),.cx(input_fmap_22[7:0]),.cy(-9'sd1),.dx(input_fmap_24[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O27_N4_S1),.chainout(chainout_4_O27));
logic signed [63:0] chainout_6_O27; 
logic signed [63:0] O27_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O27(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_25[7:0]),.ay( 9'sd1),.bx(input_fmap_28[7:0]),.by(-9'sd1),.cx(input_fmap_29[7:0]),.cy( 9'sd1),.dx(input_fmap_31[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O27_N6_S1),.chainout(chainout_6_O27));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O27_N0_S2;		always @(posedge clk) O27_N0_S2 <=     O27_N0_S1  +  O27_N2_S1 ;
 logic signed [21:0] O27_N2_S2;		always @(posedge clk) O27_N2_S2 <=     O27_N4_S1  +  O27_N6_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O27_N0_S3;		always @(posedge clk) O27_N0_S3 <=     O27_N0_S2  +  O27_N2_S2 ;
 assign conv_mac_27 = O27_N0_S3;

logic signed [31:0] conv_mac_28;
logic signed [63:0] chainout_0_O28; 
logic signed [63:0] O28_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O28(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd1),.bx(input_fmap_1[7:0]),.by(-9'sd1),.cx(input_fmap_3[7:0]),.cy( 9'sd1),.dx(input_fmap_4[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O28_N0_S1),.chainout(chainout_0_O28));
logic signed [63:0] chainout_2_O28; 
logic signed [63:0] O28_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O28(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_5[7:0]),.ay( 9'sd2),.bx(input_fmap_8[7:0]),.by( 9'sd1),.cx(input_fmap_10[7:0]),.cy( 9'sd1),.dx(input_fmap_14[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O28_N2_S1),.chainout(chainout_2_O28));
logic signed [63:0] chainout_4_O28; 
logic signed [63:0] O28_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O28(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_15[7:0]),.ay(-9'sd1),.bx(input_fmap_16[7:0]),.by( 9'sd1),.cx(input_fmap_17[7:0]),.cy( 9'sd2),.dx(input_fmap_18[7:0]),.dy( 9'sd4),.chainin(63'd0),.result(O28_N4_S1),.chainout(chainout_4_O28));
logic signed [63:0] chainout_6_O28; 
logic signed [63:0] O28_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O28(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_19[7:0]),.ay( 9'sd2),.bx(input_fmap_20[7:0]),.by( 9'sd1),.cx(input_fmap_21[7:0]),.cy(-9'sd1),.dx(input_fmap_24[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O28_N6_S1),.chainout(chainout_6_O28));
logic signed [63:0] chainout_8_O28; 
logic signed [63:0] O28_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O28(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_25[7:0]),.ay(-9'sd2),.bx(input_fmap_27[7:0]),.by(-9'sd1),.cx(input_fmap_29[7:0]),.cy(-9'sd1),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O28_N8_S1),.chainout(chainout_8_O28));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O28_N0_S2;		always @(posedge clk) O28_N0_S2 <=     O28_N0_S1  +  O28_N2_S1 ;
 logic signed [21:0] O28_N2_S2;		always @(posedge clk) O28_N2_S2 <=     O28_N4_S1  +  O28_N6_S1 ;
 logic signed [21:0] O28_N4_S2;		always @(posedge clk) O28_N4_S2 <=     O28_N8_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O28_N0_S3;		always @(posedge clk) O28_N0_S3 <=     O28_N0_S2  +  O28_N2_S2 ;
 logic signed [22:0] O28_N2_S3;		always @(posedge clk) O28_N2_S3 <=     O28_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O28_N0_S4;		always @(posedge clk) O28_N0_S4 <=     O28_N0_S3  +  O28_N2_S3 ;
 assign conv_mac_28 = O28_N0_S4;

logic signed [31:0] conv_mac_29;
logic signed [63:0] chainout_0_O29; 
logic signed [63:0] O29_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O29(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd1),.bx(input_fmap_1[7:0]),.by( 9'sd1),.cx(input_fmap_5[7:0]),.cy( 9'sd1),.dx(input_fmap_6[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O29_N0_S1),.chainout(chainout_0_O29));
logic signed [63:0] chainout_2_O29; 
logic signed [63:0] O29_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O29(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_7[7:0]),.ay(-9'sd1),.bx(input_fmap_13[7:0]),.by(-9'sd1),.cx(input_fmap_16[7:0]),.cy(-9'sd1),.dx(input_fmap_18[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O29_N2_S1),.chainout(chainout_2_O29));
logic signed [63:0] chainout_4_O29; 
logic signed [63:0] O29_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O29(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_20[7:0]),.ay( 9'sd1),.bx(input_fmap_23[7:0]),.by(-9'sd1),.cx(input_fmap_26[7:0]),.cy(-9'sd1),.dx(input_fmap_27[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O29_N4_S1),.chainout(chainout_4_O29));
logic signed [63:0] chainout_6_O29; 
logic signed [63:0] O29_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O29(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_28[7:0]),.ay(-9'sd1),.bx(input_fmap_29[7:0]),.by(-9'sd1),.cx(input_fmap_30[7:0]),.cy(-9'sd1),.dx(input_fmap_31[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O29_N6_S1),.chainout(chainout_6_O29));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O29_N0_S2;		always @(posedge clk) O29_N0_S2 <=     O29_N0_S1  +  O29_N2_S1 ;
 logic signed [21:0] O29_N2_S2;		always @(posedge clk) O29_N2_S2 <=     O29_N4_S1  +  O29_N6_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O29_N0_S3;		always @(posedge clk) O29_N0_S3 <=     O29_N0_S2  +  O29_N2_S2 ;
 assign conv_mac_29 = O29_N0_S3;

logic signed [31:0] conv_mac_30;
logic signed [63:0] chainout_0_O30; 
logic signed [63:0] O30_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O30(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_6[7:0]),.ay( 9'sd1),.bx(input_fmap_7[7:0]),.by(-9'sd1),.cx(input_fmap_9[7:0]),.cy(-9'sd1),.dx(input_fmap_12[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O30_N0_S1),.chainout(chainout_0_O30));
logic signed [63:0] chainout_2_O30; 
logic signed [63:0] O30_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O30(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_14[7:0]),.ay( 9'sd1),.bx(input_fmap_16[7:0]),.by( 9'sd2),.cx(input_fmap_20[7:0]),.cy(-9'sd1),.dx(input_fmap_22[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O30_N2_S1),.chainout(chainout_2_O30));
logic signed [63:0] chainout_4_O30; 
logic signed [63:0] O30_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O30(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_23[7:0]),.ay( 9'sd1),.bx(input_fmap_27[7:0]),.by( 9'sd1),.cx(input_fmap_30[7:0]),.cy( 9'sd2),.dx(input_fmap_31[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O30_N4_S1),.chainout(chainout_4_O30));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O30_N0_S2;		always @(posedge clk) O30_N0_S2 <=     O30_N0_S1  +  O30_N2_S1 ;
 logic signed [21:0] O30_N2_S2;		always @(posedge clk) O30_N2_S2 <=     O30_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O30_N0_S3;		always @(posedge clk) O30_N0_S3 <=     O30_N0_S2  +  O30_N2_S2 ;
 assign conv_mac_30 = O30_N0_S3;

logic signed [31:0] conv_mac_31;
logic signed [63:0] chainout_0_O31; 
logic signed [63:0] O31_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O31(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd1),.bx(input_fmap_1[7:0]),.by( 9'sd1),.cx(input_fmap_5[7:0]),.cy( 9'sd1),.dx(input_fmap_6[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O31_N0_S1),.chainout(chainout_0_O31));
logic signed [63:0] chainout_2_O31; 
logic signed [63:0] O31_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O31(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_13[7:0]),.ay( 9'sd1),.bx(input_fmap_17[7:0]),.by(-9'sd1),.cx(input_fmap_19[7:0]),.cy(-9'sd1),.dx(input_fmap_25[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O31_N2_S1),.chainout(chainout_2_O31));
logic signed [63:0] chainout_4_O31; 
logic signed [63:0] O31_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O31(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_26[7:0]),.ay( 9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O31_N4_S1),.chainout(chainout_4_O31));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O31_N0_S2;		always @(posedge clk) O31_N0_S2 <=     O31_N0_S1  +  O31_N2_S1 ;
 logic signed [21:0] O31_N2_S2;		always @(posedge clk) O31_N2_S2 <=     O31_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O31_N0_S3;		always @(posedge clk) O31_N0_S3 <=     O31_N0_S2  +  O31_N2_S2 ;
 assign conv_mac_31 = O31_N0_S3;

logic signed [31:0] conv_mac_32;
logic signed [63:0] chainout_0_O32; 
logic signed [63:0] O32_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O32(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd1),.bx(input_fmap_1[7:0]),.by(-9'sd2),.cx(input_fmap_3[7:0]),.cy(-9'sd1),.dx(input_fmap_5[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O32_N0_S1),.chainout(chainout_0_O32));
logic signed [63:0] chainout_2_O32; 
logic signed [63:0] O32_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O32(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_9[7:0]),.ay( 9'sd1),.bx(input_fmap_10[7:0]),.by( 9'sd1),.cx(input_fmap_11[7:0]),.cy(-9'sd1),.dx(input_fmap_12[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O32_N2_S1),.chainout(chainout_2_O32));
logic signed [63:0] chainout_4_O32; 
logic signed [63:0] O32_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O32(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_17[7:0]),.ay( 9'sd2),.bx(input_fmap_18[7:0]),.by( 9'sd2),.cx(input_fmap_19[7:0]),.cy( 9'sd1),.dx(input_fmap_21[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O32_N4_S1),.chainout(chainout_4_O32));
logic signed [63:0] chainout_6_O32; 
logic signed [63:0] O32_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O32(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_23[7:0]),.ay(-9'sd1),.bx(input_fmap_25[7:0]),.by(-9'sd1),.cx(input_fmap_26[7:0]),.cy(-9'sd2),.dx(input_fmap_28[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O32_N6_S1),.chainout(chainout_6_O32));
logic signed [63:0] chainout_8_O32; 
logic signed [63:0] O32_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O32(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_29[7:0]),.ay(-9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O32_N8_S1),.chainout(chainout_8_O32));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O32_N0_S2;		always @(posedge clk) O32_N0_S2 <=     O32_N0_S1  +  O32_N2_S1 ;
 logic signed [21:0] O32_N2_S2;		always @(posedge clk) O32_N2_S2 <=     O32_N4_S1  +  O32_N6_S1 ;
 logic signed [21:0] O32_N4_S2;		always @(posedge clk) O32_N4_S2 <=     O32_N8_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O32_N0_S3;		always @(posedge clk) O32_N0_S3 <=     O32_N0_S2  +  O32_N2_S2 ;
 logic signed [22:0] O32_N2_S3;		always @(posedge clk) O32_N2_S3 <=     O32_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O32_N0_S4;		always @(posedge clk) O32_N0_S4 <=     O32_N0_S3  +  O32_N2_S3 ;
 assign conv_mac_32 = O32_N0_S4;

logic signed [31:0] conv_mac_33;
logic signed [63:0] chainout_0_O33; 
logic signed [63:0] O33_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O33(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay( 9'sd2),.bx(input_fmap_7[7:0]),.by(-9'sd1),.cx(input_fmap_11[7:0]),.cy(-9'sd1),.dx(input_fmap_16[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O33_N0_S1),.chainout(chainout_0_O33));
logic signed [63:0] chainout_2_O33; 
logic signed [63:0] O33_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O33(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_18[7:0]),.ay( 9'sd1),.bx(input_fmap_22[7:0]),.by( 9'sd1),.cx(input_fmap_23[7:0]),.cy(-9'sd1),.dx(input_fmap_27[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O33_N2_S1),.chainout(chainout_2_O33));
logic signed [63:0] chainout_4_O33; 
logic signed [63:0] O33_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O33(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_28[7:0]),.ay(-9'sd1),.bx(input_fmap_31[7:0]),.by(-9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O33_N4_S1),.chainout(chainout_4_O33));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O33_N0_S2;		always @(posedge clk) O33_N0_S2 <=     O33_N0_S1  +  O33_N2_S1 ;
 logic signed [21:0] O33_N2_S2;		always @(posedge clk) O33_N2_S2 <=     O33_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O33_N0_S3;		always @(posedge clk) O33_N0_S3 <=     O33_N0_S2  +  O33_N2_S2 ;
 assign conv_mac_33 = O33_N0_S3;

logic signed [31:0] conv_mac_34;
logic signed [63:0] chainout_0_O34; 
logic signed [63:0] O34_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O34(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay(-9'sd1),.bx(input_fmap_4[7:0]),.by(-9'sd1),.cx(input_fmap_5[7:0]),.cy( 9'sd1),.dx(input_fmap_7[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O34_N0_S1),.chainout(chainout_0_O34));
logic signed [63:0] chainout_2_O34; 
logic signed [63:0] O34_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O34(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_11[7:0]),.ay( 9'sd5),.bx(input_fmap_12[7:0]),.by(-9'sd1),.cx(input_fmap_13[7:0]),.cy( 9'sd1),.dx(input_fmap_15[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O34_N2_S1),.chainout(chainout_2_O34));
logic signed [63:0] chainout_4_O34; 
logic signed [63:0] O34_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O34(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_16[7:0]),.ay( 9'sd1),.bx(input_fmap_18[7:0]),.by(-9'sd1),.cx(input_fmap_20[7:0]),.cy(-9'sd2),.dx(input_fmap_23[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O34_N4_S1),.chainout(chainout_4_O34));
logic signed [63:0] chainout_6_O34; 
logic signed [63:0] O34_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O34(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_25[7:0]),.ay( 9'sd1),.bx(input_fmap_27[7:0]),.by(-9'sd1),.cx(input_fmap_28[7:0]),.cy( 9'sd1),.dx(input_fmap_29[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O34_N6_S1),.chainout(chainout_6_O34));
logic signed [63:0] chainout_8_O34; 
logic signed [63:0] O34_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O34(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_30[7:0]),.ay( 9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O34_N8_S1),.chainout(chainout_8_O34));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O34_N0_S2;		always @(posedge clk) O34_N0_S2 <=     O34_N0_S1  +  O34_N2_S1 ;
 logic signed [21:0] O34_N2_S2;		always @(posedge clk) O34_N2_S2 <=     O34_N4_S1  +  O34_N6_S1 ;
 logic signed [21:0] O34_N4_S2;		always @(posedge clk) O34_N4_S2 <=     O34_N8_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O34_N0_S3;		always @(posedge clk) O34_N0_S3 <=     O34_N0_S2  +  O34_N2_S2 ;
 logic signed [22:0] O34_N2_S3;		always @(posedge clk) O34_N2_S3 <=     O34_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O34_N0_S4;		always @(posedge clk) O34_N0_S4 <=     O34_N0_S3  +  O34_N2_S3 ;
 assign conv_mac_34 = O34_N0_S4;

logic signed [31:0] conv_mac_35;
logic signed [63:0] chainout_0_O35; 
logic signed [63:0] O35_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O35(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd2),.bx(input_fmap_1[7:0]),.by(-9'sd1),.cx(input_fmap_2[7:0]),.cy( 9'sd1),.dx(input_fmap_6[7:0]),.dy(-9'sd3),.chainin(63'd0),.result(O35_N0_S1),.chainout(chainout_0_O35));
logic signed [63:0] chainout_2_O35; 
logic signed [63:0] O35_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O35(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_7[7:0]),.ay(-9'sd2),.bx(input_fmap_8[7:0]),.by(-9'sd1),.cx(input_fmap_10[7:0]),.cy(-9'sd1),.dx(input_fmap_11[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O35_N2_S1),.chainout(chainout_2_O35));
logic signed [63:0] chainout_4_O35; 
logic signed [63:0] O35_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O35(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_12[7:0]),.ay( 9'sd1),.bx(input_fmap_13[7:0]),.by(-9'sd1),.cx(input_fmap_15[7:0]),.cy( 9'sd1),.dx(input_fmap_16[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O35_N4_S1),.chainout(chainout_4_O35));
logic signed [63:0] chainout_6_O35; 
logic signed [63:0] O35_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O35(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_17[7:0]),.ay( 9'sd2),.bx(input_fmap_18[7:0]),.by( 9'sd2),.cx(input_fmap_19[7:0]),.cy( 9'sd1),.dx(input_fmap_21[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O35_N6_S1),.chainout(chainout_6_O35));
logic signed [63:0] chainout_8_O35; 
logic signed [63:0] O35_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O35(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_22[7:0]),.ay( 9'sd1),.bx(input_fmap_23[7:0]),.by( 9'sd1),.cx(input_fmap_26[7:0]),.cy(-9'sd1),.dx(input_fmap_27[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O35_N8_S1),.chainout(chainout_8_O35));
logic signed [63:0] chainout_10_O35; 
logic signed [63:0] O35_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O35(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_28[7:0]),.ay(-9'sd1),.bx(input_fmap_30[7:0]),.by(-9'sd2),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O35_N10_S1),.chainout(chainout_10_O35));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O35_N0_S2;		always @(posedge clk) O35_N0_S2 <=     O35_N0_S1  +  O35_N2_S1 ;
 logic signed [21:0] O35_N2_S2;		always @(posedge clk) O35_N2_S2 <=     O35_N4_S1  +  O35_N6_S1 ;
 logic signed [21:0] O35_N4_S2;		always @(posedge clk) O35_N4_S2 <=     O35_N8_S1  +  O35_N10_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O35_N0_S3;		always @(posedge clk) O35_N0_S3 <=     O35_N0_S2  +  O35_N2_S2 ;
 logic signed [22:0] O35_N2_S3;		always @(posedge clk) O35_N2_S3 <=     O35_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O35_N0_S4;		always @(posedge clk) O35_N0_S4 <=     O35_N0_S3  +  O35_N2_S3 ;
 assign conv_mac_35 = O35_N0_S4;

logic signed [31:0] conv_mac_36;
logic signed [63:0] chainout_0_O36; 
logic signed [63:0] O36_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O36(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd1),.bx(input_fmap_2[7:0]),.by(-9'sd1),.cx(input_fmap_11[7:0]),.cy(-9'sd1),.dx(input_fmap_12[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O36_N0_S1),.chainout(chainout_0_O36));
logic signed [63:0] chainout_2_O36; 
logic signed [63:0] O36_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O36(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_13[7:0]),.ay( 9'sd2),.bx(input_fmap_17[7:0]),.by(-9'sd1),.cx(input_fmap_23[7:0]),.cy( 9'sd2),.dx(input_fmap_25[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O36_N2_S1),.chainout(chainout_2_O36));
logic signed [63:0] chainout_4_O36; 
logic signed [63:0] O36_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O36(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_27[7:0]),.ay( 9'sd1),.bx(input_fmap_28[7:0]),.by(-9'sd1),.cx(input_fmap_30[7:0]),.cy(-9'sd1),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O36_N4_S1),.chainout(chainout_4_O36));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O36_N0_S2;		always @(posedge clk) O36_N0_S2 <=     O36_N0_S1  +  O36_N2_S1 ;
 logic signed [21:0] O36_N2_S2;		always @(posedge clk) O36_N2_S2 <=     O36_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O36_N0_S3;		always @(posedge clk) O36_N0_S3 <=     O36_N0_S2  +  O36_N2_S2 ;
 assign conv_mac_36 = O36_N0_S3;

logic signed [31:0] conv_mac_37;
logic signed [63:0] chainout_0_O37; 
logic signed [63:0] O37_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O37(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_2[7:0]),.ay(-9'sd1),.bx(input_fmap_7[7:0]),.by( 9'sd2),.cx(input_fmap_13[7:0]),.cy( 9'sd1),.dx(input_fmap_16[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O37_N0_S1),.chainout(chainout_0_O37));
logic signed [63:0] chainout_2_O37; 
logic signed [63:0] O37_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O37(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_17[7:0]),.ay( 9'sd1),.bx(input_fmap_22[7:0]),.by(-9'sd1),.cx(input_fmap_23[7:0]),.cy( 9'sd3),.dx(input_fmap_30[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O37_N2_S1),.chainout(chainout_2_O37));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O37_N0_S2;		always @(posedge clk) O37_N0_S2 <=     O37_N0_S1  +  O37_N2_S1 ;
 assign conv_mac_37 = O37_N0_S2;

logic signed [31:0] conv_mac_38;
logic signed [63:0] chainout_0_O38; 
logic signed [63:0] O38_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O38(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay( 9'sd1),.bx(input_fmap_2[7:0]),.by(-9'sd3),.cx(input_fmap_3[7:0]),.cy(-9'sd1),.dx(input_fmap_5[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O38_N0_S1),.chainout(chainout_0_O38));
logic signed [63:0] chainout_2_O38; 
logic signed [63:0] O38_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O38(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_8[7:0]),.ay(-9'sd1),.bx(input_fmap_14[7:0]),.by(-9'sd1),.cx(input_fmap_15[7:0]),.cy( 9'sd1),.dx(input_fmap_16[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O38_N2_S1),.chainout(chainout_2_O38));
logic signed [63:0] chainout_4_O38; 
logic signed [63:0] O38_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O38(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_19[7:0]),.ay(-9'sd1),.bx(input_fmap_22[7:0]),.by( 9'sd2),.cx(input_fmap_23[7:0]),.cy(-9'sd4),.dx(input_fmap_25[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O38_N4_S1),.chainout(chainout_4_O38));
logic signed [63:0] chainout_6_O38; 
logic signed [63:0] O38_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O38(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_27[7:0]),.ay( 9'sd1),.bx(input_fmap_28[7:0]),.by(-9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O38_N6_S1),.chainout(chainout_6_O38));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O38_N0_S2;		always @(posedge clk) O38_N0_S2 <=     O38_N0_S1  +  O38_N2_S1 ;
 logic signed [21:0] O38_N2_S2;		always @(posedge clk) O38_N2_S2 <=     O38_N4_S1  +  O38_N6_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O38_N0_S3;		always @(posedge clk) O38_N0_S3 <=     O38_N0_S2  +  O38_N2_S2 ;
 assign conv_mac_38 = O38_N0_S3;

logic signed [31:0] conv_mac_39;
logic signed [63:0] chainout_0_O39; 
logic signed [63:0] O39_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O39(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd2),.bx(input_fmap_1[7:0]),.by( 9'sd4),.cx(input_fmap_4[7:0]),.cy( 9'sd1),.dx(input_fmap_7[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O39_N0_S1),.chainout(chainout_0_O39));
logic signed [63:0] chainout_2_O39; 
logic signed [63:0] O39_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O39(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_9[7:0]),.ay( 9'sd1),.bx(input_fmap_10[7:0]),.by( 9'sd1),.cx(input_fmap_11[7:0]),.cy(-9'sd2),.dx(input_fmap_13[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O39_N2_S1),.chainout(chainout_2_O39));
logic signed [63:0] chainout_4_O39; 
logic signed [63:0] O39_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O39(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_14[7:0]),.ay( 9'sd1),.bx(input_fmap_16[7:0]),.by(-9'sd1),.cx(input_fmap_17[7:0]),.cy(-9'sd1),.dx(input_fmap_18[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O39_N4_S1),.chainout(chainout_4_O39));
logic signed [63:0] chainout_6_O39; 
logic signed [63:0] O39_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O39(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_19[7:0]),.ay(-9'sd2),.bx(input_fmap_23[7:0]),.by(-9'sd1),.cx(input_fmap_25[7:0]),.cy(-9'sd1),.dx(input_fmap_26[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O39_N6_S1),.chainout(chainout_6_O39));
logic signed [63:0] chainout_8_O39; 
logic signed [63:0] O39_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O39(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_29[7:0]),.ay(-9'sd1),.bx(input_fmap_30[7:0]),.by(-9'sd1),.cx(input_fmap_31[7:0]),.cy( 9'sd1),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O39_N8_S1),.chainout(chainout_8_O39));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O39_N0_S2;		always @(posedge clk) O39_N0_S2 <=     O39_N0_S1  +  O39_N2_S1 ;
 logic signed [21:0] O39_N2_S2;		always @(posedge clk) O39_N2_S2 <=     O39_N4_S1  +  O39_N6_S1 ;
 logic signed [21:0] O39_N4_S2;		always @(posedge clk) O39_N4_S2 <=     O39_N8_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O39_N0_S3;		always @(posedge clk) O39_N0_S3 <=     O39_N0_S2  +  O39_N2_S2 ;
 logic signed [22:0] O39_N2_S3;		always @(posedge clk) O39_N2_S3 <=     O39_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O39_N0_S4;		always @(posedge clk) O39_N0_S4 <=     O39_N0_S3  +  O39_N2_S3 ;
 assign conv_mac_39 = O39_N0_S4;

logic signed [31:0] conv_mac_40;
logic signed [63:0] chainout_0_O40; 
logic signed [63:0] O40_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O40(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_7[7:0]),.ay( 9'sd1),.bx(input_fmap_13[7:0]),.by( 9'sd3),.cx(input_fmap_23[7:0]),.cy( 9'sd2),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O40_N0_S1),.chainout(chainout_0_O40));
assign conv_mac_40 = O40_N0_S1;

logic signed [31:0] conv_mac_41;
logic signed [63:0] chainout_0_O41; 
logic signed [63:0] O41_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O41(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd1),.bx(input_fmap_5[7:0]),.by(-9'sd1),.cx(input_fmap_7[7:0]),.cy(-9'sd1),.dx(input_fmap_11[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O41_N0_S1),.chainout(chainout_0_O41));
logic signed [63:0] chainout_2_O41; 
logic signed [63:0] O41_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O41(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_13[7:0]),.ay(-9'sd1),.bx(input_fmap_18[7:0]),.by(-9'sd1),.cx(input_fmap_22[7:0]),.cy(-9'sd1),.dx(input_fmap_23[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O41_N2_S1),.chainout(chainout_2_O41));
logic signed [63:0] chainout_4_O41; 
logic signed [63:0] O41_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O41(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_25[7:0]),.ay(-9'sd1),.bx(input_fmap_27[7:0]),.by( 9'sd2),.cx(input_fmap_28[7:0]),.cy(-9'sd2),.dx(input_fmap_29[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O41_N4_S1),.chainout(chainout_4_O41));
logic signed [63:0] chainout_6_O41; 
logic signed [63:0] O41_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O41(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_30[7:0]),.ay( 9'sd2),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O41_N6_S1),.chainout(chainout_6_O41));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O41_N0_S2;		always @(posedge clk) O41_N0_S2 <=     O41_N0_S1  +  O41_N2_S1 ;
 logic signed [21:0] O41_N2_S2;		always @(posedge clk) O41_N2_S2 <=     O41_N4_S1  +  O41_N6_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O41_N0_S3;		always @(posedge clk) O41_N0_S3 <=     O41_N0_S2  +  O41_N2_S2 ;
 assign conv_mac_41 = O41_N0_S3;

logic signed [31:0] conv_mac_42;
logic signed [63:0] chainout_0_O42; 
logic signed [63:0] O42_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O42(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd1),.bx(input_fmap_1[7:0]),.by( 9'sd3),.cx(input_fmap_15[7:0]),.cy( 9'sd1),.dx(input_fmap_19[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O42_N0_S1),.chainout(chainout_0_O42));
logic signed [63:0] chainout_2_O42; 
logic signed [63:0] O42_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O42(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_21[7:0]),.ay( 9'sd1),.bx(input_fmap_23[7:0]),.by(-9'sd1),.cx(input_fmap_25[7:0]),.cy(-9'sd1),.dx(input_fmap_27[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O42_N2_S1),.chainout(chainout_2_O42));
logic signed [63:0] chainout_4_O42; 
logic signed [63:0] O42_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O42(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_31[7:0]),.ay(-9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O42_N4_S1),.chainout(chainout_4_O42));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O42_N0_S2;		always @(posedge clk) O42_N0_S2 <=     O42_N0_S1  +  O42_N2_S1 ;
 logic signed [21:0] O42_N2_S2;		always @(posedge clk) O42_N2_S2 <=     O42_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O42_N0_S3;		always @(posedge clk) O42_N0_S3 <=     O42_N0_S2  +  O42_N2_S2 ;
 assign conv_mac_42 = O42_N0_S3;

logic signed [31:0] conv_mac_43;
logic signed [63:0] chainout_0_O43; 
logic signed [63:0] O43_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O43(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_4[7:0]),.ay( 9'sd1),.bx(input_fmap_5[7:0]),.by(-9'sd1),.cx(input_fmap_6[7:0]),.cy(-9'sd1),.dx(input_fmap_8[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O43_N0_S1),.chainout(chainout_0_O43));
logic signed [63:0] chainout_2_O43; 
logic signed [63:0] O43_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O43(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_11[7:0]),.ay( 9'sd1),.bx(input_fmap_13[7:0]),.by( 9'sd1),.cx(input_fmap_17[7:0]),.cy( 9'sd2),.dx(input_fmap_18[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O43_N2_S1),.chainout(chainout_2_O43));
logic signed [63:0] chainout_4_O43; 
logic signed [63:0] O43_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O43(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_20[7:0]),.ay(-9'sd1),.bx(input_fmap_26[7:0]),.by(-9'sd1),.cx(input_fmap_29[7:0]),.cy(-9'sd1),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O43_N4_S1),.chainout(chainout_4_O43));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O43_N0_S2;		always @(posedge clk) O43_N0_S2 <=     O43_N0_S1  +  O43_N2_S1 ;
 logic signed [21:0] O43_N2_S2;		always @(posedge clk) O43_N2_S2 <=     O43_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O43_N0_S3;		always @(posedge clk) O43_N0_S3 <=     O43_N0_S2  +  O43_N2_S2 ;
 assign conv_mac_43 = O43_N0_S3;

logic signed [31:0] conv_mac_44;
logic signed [63:0] chainout_0_O44; 
logic signed [63:0] O44_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O44(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd2),.bx(input_fmap_1[7:0]),.by( 9'sd2),.cx(input_fmap_2[7:0]),.cy(-9'sd1),.dx(input_fmap_4[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O44_N0_S1),.chainout(chainout_0_O44));
logic signed [63:0] chainout_2_O44; 
logic signed [63:0] O44_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O44(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_5[7:0]),.ay(-9'sd1),.bx(input_fmap_6[7:0]),.by(-9'sd1),.cx(input_fmap_7[7:0]),.cy(-9'sd3),.dx(input_fmap_8[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O44_N2_S1),.chainout(chainout_2_O44));
logic signed [63:0] chainout_4_O44; 
logic signed [63:0] O44_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O44(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_9[7:0]),.ay(-9'sd1),.bx(input_fmap_10[7:0]),.by( 9'sd1),.cx(input_fmap_11[7:0]),.cy( 9'sd2),.dx(input_fmap_13[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O44_N4_S1),.chainout(chainout_4_O44));
logic signed [63:0] chainout_6_O44; 
logic signed [63:0] O44_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O44(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_14[7:0]),.ay(-9'sd2),.bx(input_fmap_15[7:0]),.by(-9'sd2),.cx(input_fmap_16[7:0]),.cy(-9'sd2),.dx(input_fmap_17[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O44_N6_S1),.chainout(chainout_6_O44));
logic signed [63:0] chainout_8_O44; 
logic signed [63:0] O44_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O44(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_18[7:0]),.ay(-9'sd1),.bx(input_fmap_19[7:0]),.by(-9'sd2),.cx(input_fmap_20[7:0]),.cy(-9'sd3),.dx(input_fmap_21[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O44_N8_S1),.chainout(chainout_8_O44));
logic signed [63:0] chainout_10_O44; 
logic signed [63:0] O44_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O44(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_22[7:0]),.ay(-9'sd1),.bx(input_fmap_25[7:0]),.by(-9'sd5),.cx(input_fmap_26[7:0]),.cy(-9'sd1),.dx(input_fmap_27[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O44_N10_S1),.chainout(chainout_10_O44));
logic signed [63:0] chainout_12_O44; 
logic signed [63:0] O44_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O44(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_28[7:0]),.ay( 9'sd4),.bx(input_fmap_30[7:0]),.by(-9'sd2),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O44_N12_S1),.chainout(chainout_12_O44));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O44_N0_S2;		always @(posedge clk) O44_N0_S2 <=     O44_N0_S1  +  O44_N2_S1 ;
 logic signed [21:0] O44_N2_S2;		always @(posedge clk) O44_N2_S2 <=     O44_N4_S1  +  O44_N6_S1 ;
 logic signed [21:0] O44_N4_S2;		always @(posedge clk) O44_N4_S2 <=     O44_N8_S1  +  O44_N10_S1 ;
 logic signed [21:0] O44_N6_S2;		always @(posedge clk) O44_N6_S2 <=     O44_N12_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O44_N0_S3;		always @(posedge clk) O44_N0_S3 <=     O44_N0_S2  +  O44_N2_S2 ;
 logic signed [22:0] O44_N2_S3;		always @(posedge clk) O44_N2_S3 <=     O44_N4_S2  +  O44_N6_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O44_N0_S4;		always @(posedge clk) O44_N0_S4 <=     O44_N0_S3  +  O44_N2_S3 ;
 assign conv_mac_44 = O44_N0_S4;

logic signed [31:0] conv_mac_45;
logic signed [63:0] chainout_0_O45; 
logic signed [63:0] O45_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O45(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay( 9'sd1),.bx(input_fmap_3[7:0]),.by( 9'sd1),.cx(input_fmap_7[7:0]),.cy( 9'sd4),.dx(input_fmap_10[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O45_N0_S1),.chainout(chainout_0_O45));
logic signed [63:0] chainout_2_O45; 
logic signed [63:0] O45_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O45(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_11[7:0]),.ay( 9'sd1),.bx(input_fmap_14[7:0]),.by( 9'sd1),.cx(input_fmap_16[7:0]),.cy(-9'sd1),.dx(input_fmap_17[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O45_N2_S1),.chainout(chainout_2_O45));
logic signed [63:0] chainout_4_O45; 
logic signed [63:0] O45_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O45(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_20[7:0]),.ay(-9'sd1),.bx(input_fmap_21[7:0]),.by( 9'sd2),.cx(input_fmap_22[7:0]),.cy( 9'sd1),.dx(input_fmap_23[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O45_N4_S1),.chainout(chainout_4_O45));
logic signed [63:0] chainout_6_O45; 
logic signed [63:0] O45_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O45(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_24[7:0]),.ay( 9'sd1),.bx(input_fmap_27[7:0]),.by(-9'sd1),.cx(input_fmap_28[7:0]),.cy( 9'sd3),.dx(input_fmap_30[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O45_N6_S1),.chainout(chainout_6_O45));
logic signed [63:0] chainout_8_O45; 
logic signed [63:0] O45_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O45(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_31[7:0]),.ay( 9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O45_N8_S1),.chainout(chainout_8_O45));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O45_N0_S2;		always @(posedge clk) O45_N0_S2 <=     O45_N0_S1  +  O45_N2_S1 ;
 logic signed [21:0] O45_N2_S2;		always @(posedge clk) O45_N2_S2 <=     O45_N4_S1  +  O45_N6_S1 ;
 logic signed [21:0] O45_N4_S2;		always @(posedge clk) O45_N4_S2 <=     O45_N8_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O45_N0_S3;		always @(posedge clk) O45_N0_S3 <=     O45_N0_S2  +  O45_N2_S2 ;
 logic signed [22:0] O45_N2_S3;		always @(posedge clk) O45_N2_S3 <=     O45_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O45_N0_S4;		always @(posedge clk) O45_N0_S4 <=     O45_N0_S3  +  O45_N2_S3 ;
 assign conv_mac_45 = O45_N0_S4;

logic signed [31:0] conv_mac_46;
logic signed [63:0] chainout_0_O46; 
logic signed [63:0] O46_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O46(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay( 9'sd1),.bx(input_fmap_17[7:0]),.by( 9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O46_N0_S1),.chainout(chainout_0_O46));
assign conv_mac_46 = O46_N0_S1;

logic signed [31:0] conv_mac_47;
logic signed [63:0] chainout_0_O47; 
logic signed [63:0] O47_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O47(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_2[7:0]),.ay( 9'sd1),.bx(input_fmap_7[7:0]),.by( 9'sd1),.cx(input_fmap_11[7:0]),.cy(-9'sd1),.dx(input_fmap_14[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O47_N0_S1),.chainout(chainout_0_O47));
logic signed [63:0] chainout_2_O47; 
logic signed [63:0] O47_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O47(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_18[7:0]),.ay( 9'sd1),.bx(input_fmap_26[7:0]),.by(-9'sd1),.cx(input_fmap_27[7:0]),.cy( 9'sd1),.dx(input_fmap_28[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O47_N2_S1),.chainout(chainout_2_O47));
logic signed [63:0] chainout_4_O47; 
logic signed [63:0] O47_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O47(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_30[7:0]),.ay( 9'sd1),.bx(input_fmap_31[7:0]),.by(-9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O47_N4_S1),.chainout(chainout_4_O47));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O47_N0_S2;		always @(posedge clk) O47_N0_S2 <=     O47_N0_S1  +  O47_N2_S1 ;
 logic signed [21:0] O47_N2_S2;		always @(posedge clk) O47_N2_S2 <=     O47_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O47_N0_S3;		always @(posedge clk) O47_N0_S3 <=     O47_N0_S2  +  O47_N2_S2 ;
 assign conv_mac_47 = O47_N0_S3;

logic signed [31:0] conv_mac_48;
logic signed [63:0] chainout_0_O48; 
logic signed [63:0] O48_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O48(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay( 9'sd2),.bx(input_fmap_4[7:0]),.by(-9'sd1),.cx(input_fmap_5[7:0]),.cy(-9'sd1),.dx(input_fmap_6[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O48_N0_S1),.chainout(chainout_0_O48));
logic signed [63:0] chainout_2_O48; 
logic signed [63:0] O48_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O48(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_7[7:0]),.ay(-9'sd1),.bx(input_fmap_11[7:0]),.by(-9'sd1),.cx(input_fmap_12[7:0]),.cy(-9'sd1),.dx(input_fmap_13[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O48_N2_S1),.chainout(chainout_2_O48));
logic signed [63:0] chainout_4_O48; 
logic signed [63:0] O48_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O48(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_18[7:0]),.ay(-9'sd2),.bx(input_fmap_19[7:0]),.by(-9'sd1),.cx(input_fmap_20[7:0]),.cy(-9'sd1),.dx(input_fmap_21[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O48_N4_S1),.chainout(chainout_4_O48));
logic signed [63:0] chainout_6_O48; 
logic signed [63:0] O48_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O48(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_22[7:0]),.ay(-9'sd1),.bx(input_fmap_24[7:0]),.by(-9'sd1),.cx(input_fmap_26[7:0]),.cy( 9'sd2),.dx(input_fmap_29[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O48_N6_S1),.chainout(chainout_6_O48));
logic signed [63:0] chainout_8_O48; 
logic signed [63:0] O48_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O48(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_31[7:0]),.ay( 9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O48_N8_S1),.chainout(chainout_8_O48));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O48_N0_S2;		always @(posedge clk) O48_N0_S2 <=     O48_N0_S1  +  O48_N2_S1 ;
 logic signed [21:0] O48_N2_S2;		always @(posedge clk) O48_N2_S2 <=     O48_N4_S1  +  O48_N6_S1 ;
 logic signed [21:0] O48_N4_S2;		always @(posedge clk) O48_N4_S2 <=     O48_N8_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O48_N0_S3;		always @(posedge clk) O48_N0_S3 <=     O48_N0_S2  +  O48_N2_S2 ;
 logic signed [22:0] O48_N2_S3;		always @(posedge clk) O48_N2_S3 <=     O48_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O48_N0_S4;		always @(posedge clk) O48_N0_S4 <=     O48_N0_S3  +  O48_N2_S3 ;
 assign conv_mac_48 = O48_N0_S4;

logic signed [31:0] conv_mac_49;
logic signed [63:0] chainout_0_O49; 
logic signed [63:0] O49_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O49(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay(-9'sd4),.bx(input_fmap_3[7:0]),.by(-9'sd1),.cx(input_fmap_5[7:0]),.cy(-9'sd1),.dx(input_fmap_6[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O49_N0_S1),.chainout(chainout_0_O49));
logic signed [63:0] chainout_2_O49; 
logic signed [63:0] O49_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O49(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_7[7:0]),.ay( 9'sd2),.bx(input_fmap_9[7:0]),.by( 9'sd1),.cx(input_fmap_10[7:0]),.cy(-9'sd1),.dx(input_fmap_11[7:0]),.dy(-9'sd3),.chainin(63'd0),.result(O49_N2_S1),.chainout(chainout_2_O49));
logic signed [63:0] chainout_4_O49; 
logic signed [63:0] O49_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O49(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_12[7:0]),.ay( 9'sd1),.bx(input_fmap_13[7:0]),.by(-9'sd1),.cx(input_fmap_15[7:0]),.cy( 9'sd2),.dx(input_fmap_16[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O49_N4_S1),.chainout(chainout_4_O49));
logic signed [63:0] chainout_6_O49; 
logic signed [63:0] O49_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O49(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_17[7:0]),.ay(-9'sd3),.bx(input_fmap_18[7:0]),.by(-9'sd1),.cx(input_fmap_19[7:0]),.cy( 9'sd2),.dx(input_fmap_21[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O49_N6_S1),.chainout(chainout_6_O49));
logic signed [63:0] chainout_8_O49; 
logic signed [63:0] O49_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O49(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_22[7:0]),.ay(-9'sd1),.bx(input_fmap_24[7:0]),.by(-9'sd2),.cx(input_fmap_25[7:0]),.cy( 9'sd3),.dx(input_fmap_26[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O49_N8_S1),.chainout(chainout_8_O49));
logic signed [63:0] chainout_10_O49; 
logic signed [63:0] O49_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O49(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_28[7:0]),.ay(-9'sd1),.bx(input_fmap_29[7:0]),.by( 9'sd2),.cx(input_fmap_31[7:0]),.cy( 9'sd2),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O49_N10_S1),.chainout(chainout_10_O49));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O49_N0_S2;		always @(posedge clk) O49_N0_S2 <=     O49_N0_S1  +  O49_N2_S1 ;
 logic signed [21:0] O49_N2_S2;		always @(posedge clk) O49_N2_S2 <=     O49_N4_S1  +  O49_N6_S1 ;
 logic signed [21:0] O49_N4_S2;		always @(posedge clk) O49_N4_S2 <=     O49_N8_S1  +  O49_N10_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O49_N0_S3;		always @(posedge clk) O49_N0_S3 <=     O49_N0_S2  +  O49_N2_S2 ;
 logic signed [22:0] O49_N2_S3;		always @(posedge clk) O49_N2_S3 <=     O49_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O49_N0_S4;		always @(posedge clk) O49_N0_S4 <=     O49_N0_S3  +  O49_N2_S3 ;
 assign conv_mac_49 = O49_N0_S4;

logic signed [31:0] conv_mac_50;
logic signed [63:0] chainout_0_O50; 
logic signed [63:0] O50_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O50(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd1),.bx(input_fmap_1[7:0]),.by(-9'sd3),.cx(input_fmap_2[7:0]),.cy(-9'sd1),.dx(input_fmap_5[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O50_N0_S1),.chainout(chainout_0_O50));
logic signed [63:0] chainout_2_O50; 
logic signed [63:0] O50_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O50(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_7[7:0]),.ay(-9'sd1),.bx(input_fmap_11[7:0]),.by(-9'sd3),.cx(input_fmap_12[7:0]),.cy(-9'sd1),.dx(input_fmap_15[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O50_N2_S1),.chainout(chainout_2_O50));
logic signed [63:0] chainout_4_O50; 
logic signed [63:0] O50_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O50(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_22[7:0]),.ay(-9'sd1),.bx(input_fmap_23[7:0]),.by( 9'sd1),.cx(input_fmap_25[7:0]),.cy( 9'sd1),.dx(input_fmap_26[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O50_N4_S1),.chainout(chainout_4_O50));
logic signed [63:0] chainout_6_O50; 
logic signed [63:0] O50_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O50(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_27[7:0]),.ay( 9'sd1),.bx(input_fmap_28[7:0]),.by(-9'sd2),.cx(input_fmap_31[7:0]),.cy(-9'sd1),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O50_N6_S1),.chainout(chainout_6_O50));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O50_N0_S2;		always @(posedge clk) O50_N0_S2 <=     O50_N0_S1  +  O50_N2_S1 ;
 logic signed [21:0] O50_N2_S2;		always @(posedge clk) O50_N2_S2 <=     O50_N4_S1  +  O50_N6_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O50_N0_S3;		always @(posedge clk) O50_N0_S3 <=     O50_N0_S2  +  O50_N2_S2 ;
 assign conv_mac_50 = O50_N0_S3;

logic signed [31:0] conv_mac_51;
logic signed [63:0] chainout_0_O51; 
logic signed [63:0] O51_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O51(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd1),.bx(input_fmap_1[7:0]),.by(-9'sd1),.cx(input_fmap_2[7:0]),.cy( 9'sd1),.dx(input_fmap_4[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O51_N0_S1),.chainout(chainout_0_O51));
logic signed [63:0] chainout_2_O51; 
logic signed [63:0] O51_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O51(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_5[7:0]),.ay( 9'sd1),.bx(input_fmap_7[7:0]),.by(-9'sd1),.cx(input_fmap_8[7:0]),.cy( 9'sd1),.dx(input_fmap_10[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O51_N2_S1),.chainout(chainout_2_O51));
logic signed [63:0] chainout_4_O51; 
logic signed [63:0] O51_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O51(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_13[7:0]),.ay(-9'sd1),.bx(input_fmap_14[7:0]),.by(-9'sd1),.cx(input_fmap_17[7:0]),.cy( 9'sd1),.dx(input_fmap_18[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O51_N4_S1),.chainout(chainout_4_O51));
logic signed [63:0] chainout_6_O51; 
logic signed [63:0] O51_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O51(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_21[7:0]),.ay(-9'sd1),.bx(input_fmap_26[7:0]),.by( 9'sd2),.cx(input_fmap_27[7:0]),.cy(-9'sd2),.dx(input_fmap_29[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O51_N6_S1),.chainout(chainout_6_O51));
logic signed [63:0] chainout_8_O51; 
logic signed [63:0] O51_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O51(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_30[7:0]),.ay(-9'sd1),.bx(input_fmap_31[7:0]),.by( 9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O51_N8_S1),.chainout(chainout_8_O51));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O51_N0_S2;		always @(posedge clk) O51_N0_S2 <=     O51_N0_S1  +  O51_N2_S1 ;
 logic signed [21:0] O51_N2_S2;		always @(posedge clk) O51_N2_S2 <=     O51_N4_S1  +  O51_N6_S1 ;
 logic signed [21:0] O51_N4_S2;		always @(posedge clk) O51_N4_S2 <=     O51_N8_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O51_N0_S3;		always @(posedge clk) O51_N0_S3 <=     O51_N0_S2  +  O51_N2_S2 ;
 logic signed [22:0] O51_N2_S3;		always @(posedge clk) O51_N2_S3 <=     O51_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O51_N0_S4;		always @(posedge clk) O51_N0_S4 <=     O51_N0_S3  +  O51_N2_S3 ;
 assign conv_mac_51 = O51_N0_S4;

logic signed [31:0] conv_mac_52;
logic signed [63:0] chainout_0_O52; 
logic signed [63:0] O52_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O52(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_2[7:0]),.ay(-9'sd1),.bx(input_fmap_5[7:0]),.by(-9'sd1),.cx(input_fmap_7[7:0]),.cy( 9'sd1),.dx(input_fmap_13[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O52_N0_S1),.chainout(chainout_0_O52));
logic signed [63:0] chainout_2_O52; 
logic signed [63:0] O52_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O52(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_16[7:0]),.ay(-9'sd2),.bx(input_fmap_17[7:0]),.by( 9'sd1),.cx(input_fmap_19[7:0]),.cy( 9'sd1),.dx(input_fmap_20[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O52_N2_S1),.chainout(chainout_2_O52));
logic signed [63:0] chainout_4_O52; 
logic signed [63:0] O52_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O52(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_21[7:0]),.ay(-9'sd2),.bx(input_fmap_23[7:0]),.by( 9'sd2),.cx(input_fmap_25[7:0]),.cy( 9'sd1),.dx(input_fmap_26[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O52_N4_S1),.chainout(chainout_4_O52));
logic signed [63:0] chainout_6_O52; 
logic signed [63:0] O52_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O52(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_27[7:0]),.ay(-9'sd1),.bx(input_fmap_28[7:0]),.by( 9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O52_N6_S1),.chainout(chainout_6_O52));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O52_N0_S2;		always @(posedge clk) O52_N0_S2 <=     O52_N0_S1  +  O52_N2_S1 ;
 logic signed [21:0] O52_N2_S2;		always @(posedge clk) O52_N2_S2 <=     O52_N4_S1  +  O52_N6_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O52_N0_S3;		always @(posedge clk) O52_N0_S3 <=     O52_N0_S2  +  O52_N2_S2 ;
 assign conv_mac_52 = O52_N0_S3;

logic signed [31:0] conv_mac_53;
logic signed [63:0] chainout_0_O53; 
logic signed [63:0] O53_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O53(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_6[7:0]),.ay( 9'sd2),.bx(input_fmap_12[7:0]),.by(-9'sd1),.cx(input_fmap_13[7:0]),.cy(-9'sd1),.dx(input_fmap_20[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O53_N0_S1),.chainout(chainout_0_O53));
logic signed [63:0] chainout_2_O53; 
logic signed [63:0] O53_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O53(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_23[7:0]),.ay(-9'sd1),.bx(input_fmap_25[7:0]),.by(-9'sd1),.cx(input_fmap_26[7:0]),.cy(-9'sd1),.dx(input_fmap_30[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O53_N2_S1),.chainout(chainout_2_O53));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O53_N0_S2;		always @(posedge clk) O53_N0_S2 <=     O53_N0_S1  +  O53_N2_S1 ;
 assign conv_mac_53 = O53_N0_S2;

logic signed [31:0] conv_mac_54;
logic signed [63:0] chainout_0_O54; 
logic signed [63:0] O54_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O54(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd2),.bx(input_fmap_1[7:0]),.by( 9'sd2),.cx(input_fmap_2[7:0]),.cy( 9'sd1),.dx(input_fmap_5[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O54_N0_S1),.chainout(chainout_0_O54));
logic signed [63:0] chainout_2_O54; 
logic signed [63:0] O54_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O54(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_6[7:0]),.ay( 9'sd2),.bx(input_fmap_12[7:0]),.by(-9'sd1),.cx(input_fmap_14[7:0]),.cy( 9'sd2),.dx(input_fmap_15[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O54_N2_S1),.chainout(chainout_2_O54));
logic signed [63:0] chainout_4_O54; 
logic signed [63:0] O54_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O54(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_16[7:0]),.ay(-9'sd1),.bx(input_fmap_18[7:0]),.by(-9'sd1),.cx(input_fmap_19[7:0]),.cy(-9'sd1),.dx(input_fmap_21[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O54_N4_S1),.chainout(chainout_4_O54));
logic signed [63:0] chainout_6_O54; 
logic signed [63:0] O54_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O54(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_23[7:0]),.ay( 9'sd1),.bx(input_fmap_24[7:0]),.by( 9'sd1),.cx(input_fmap_25[7:0]),.cy( 9'sd1),.dx(input_fmap_26[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O54_N6_S1),.chainout(chainout_6_O54));
logic signed [63:0] chainout_8_O54; 
logic signed [63:0] O54_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O54(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_27[7:0]),.ay(-9'sd1),.bx(input_fmap_31[7:0]),.by( 9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O54_N8_S1),.chainout(chainout_8_O54));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O54_N0_S2;		always @(posedge clk) O54_N0_S2 <=     O54_N0_S1  +  O54_N2_S1 ;
 logic signed [21:0] O54_N2_S2;		always @(posedge clk) O54_N2_S2 <=     O54_N4_S1  +  O54_N6_S1 ;
 logic signed [21:0] O54_N4_S2;		always @(posedge clk) O54_N4_S2 <=     O54_N8_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O54_N0_S3;		always @(posedge clk) O54_N0_S3 <=     O54_N0_S2  +  O54_N2_S2 ;
 logic signed [22:0] O54_N2_S3;		always @(posedge clk) O54_N2_S3 <=     O54_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O54_N0_S4;		always @(posedge clk) O54_N0_S4 <=     O54_N0_S3  +  O54_N2_S3 ;
 assign conv_mac_54 = O54_N0_S4;

logic signed [31:0] conv_mac_55;
logic signed [63:0] chainout_0_O55; 
logic signed [63:0] O55_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O55(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_2[7:0]),.ay( 9'sd3),.bx(input_fmap_3[7:0]),.by(-9'sd2),.cx(input_fmap_5[7:0]),.cy(-9'sd1),.dx(input_fmap_6[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O55_N0_S1),.chainout(chainout_0_O55));
logic signed [63:0] chainout_2_O55; 
logic signed [63:0] O55_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O55(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_7[7:0]),.ay(-9'sd2),.bx(input_fmap_8[7:0]),.by( 9'sd1),.cx(input_fmap_10[7:0]),.cy(-9'sd1),.dx(input_fmap_11[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O55_N2_S1),.chainout(chainout_2_O55));
logic signed [63:0] chainout_4_O55; 
logic signed [63:0] O55_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O55(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_13[7:0]),.ay(-9'sd1),.bx(input_fmap_14[7:0]),.by(-9'sd1),.cx(input_fmap_16[7:0]),.cy( 9'sd1),.dx(input_fmap_19[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O55_N4_S1),.chainout(chainout_4_O55));
logic signed [63:0] chainout_6_O55; 
logic signed [63:0] O55_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O55(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_21[7:0]),.ay(-9'sd1),.bx(input_fmap_26[7:0]),.by(-9'sd1),.cx(input_fmap_27[7:0]),.cy( 9'sd1),.dx(input_fmap_30[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O55_N6_S1),.chainout(chainout_6_O55));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O55_N0_S2;		always @(posedge clk) O55_N0_S2 <=     O55_N0_S1  +  O55_N2_S1 ;
 logic signed [21:0] O55_N2_S2;		always @(posedge clk) O55_N2_S2 <=     O55_N4_S1  +  O55_N6_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O55_N0_S3;		always @(posedge clk) O55_N0_S3 <=     O55_N0_S2  +  O55_N2_S2 ;
 assign conv_mac_55 = O55_N0_S3;

logic signed [31:0] conv_mac_56;
logic signed [63:0] chainout_0_O56; 
logic signed [63:0] O56_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O56(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_2[7:0]),.ay( 9'sd2),.bx(input_fmap_6[7:0]),.by(-9'sd1),.cx(input_fmap_7[7:0]),.cy( 9'sd3),.dx(input_fmap_13[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O56_N0_S1),.chainout(chainout_0_O56));
logic signed [63:0] chainout_2_O56; 
logic signed [63:0] O56_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O56(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_14[7:0]),.ay(-9'sd1),.bx(input_fmap_16[7:0]),.by(-9'sd1),.cx(input_fmap_17[7:0]),.cy(-9'sd2),.dx(input_fmap_20[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O56_N2_S1),.chainout(chainout_2_O56));
logic signed [63:0] chainout_4_O56; 
logic signed [63:0] O56_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O56(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_21[7:0]),.ay( 9'sd1),.bx(input_fmap_23[7:0]),.by(-9'sd1),.cx(input_fmap_27[7:0]),.cy(-9'sd1),.dx(input_fmap_28[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O56_N4_S1),.chainout(chainout_4_O56));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O56_N0_S2;		always @(posedge clk) O56_N0_S2 <=     O56_N0_S1  +  O56_N2_S1 ;
 logic signed [21:0] O56_N2_S2;		always @(posedge clk) O56_N2_S2 <=     O56_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O56_N0_S3;		always @(posedge clk) O56_N0_S3 <=     O56_N0_S2  +  O56_N2_S2 ;
 assign conv_mac_56 = O56_N0_S3;

logic signed [31:0] conv_mac_57;
logic signed [63:0] chainout_0_O57; 
logic signed [63:0] O57_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O57(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay(-9'sd1),.bx(input_fmap_2[7:0]),.by(-9'sd3),.cx(input_fmap_3[7:0]),.cy(-9'sd2),.dx(input_fmap_7[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O57_N0_S1),.chainout(chainout_0_O57));
logic signed [63:0] chainout_2_O57; 
logic signed [63:0] O57_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O57(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_10[7:0]),.ay(-9'sd1),.bx(input_fmap_11[7:0]),.by(-9'sd1),.cx(input_fmap_16[7:0]),.cy(-9'sd1),.dx(input_fmap_17[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O57_N2_S1),.chainout(chainout_2_O57));
logic signed [63:0] chainout_4_O57; 
logic signed [63:0] O57_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O57(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_19[7:0]),.ay( 9'sd1),.bx(input_fmap_20[7:0]),.by( 9'sd1),.cx(input_fmap_21[7:0]),.cy(-9'sd1),.dx(input_fmap_22[7:0]),.dy(-9'sd3),.chainin(63'd0),.result(O57_N4_S1),.chainout(chainout_4_O57));
logic signed [63:0] chainout_6_O57; 
logic signed [63:0] O57_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O57(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_23[7:0]),.ay( 9'sd4),.bx(input_fmap_27[7:0]),.by( 9'sd1),.cx(input_fmap_28[7:0]),.cy(-9'sd1),.dx(input_fmap_29[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O57_N6_S1),.chainout(chainout_6_O57));
logic signed [63:0] chainout_8_O57; 
logic signed [63:0] O57_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O57(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_30[7:0]),.ay( 9'sd2),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O57_N8_S1),.chainout(chainout_8_O57));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O57_N0_S2;		always @(posedge clk) O57_N0_S2 <=     O57_N0_S1  +  O57_N2_S1 ;
 logic signed [21:0] O57_N2_S2;		always @(posedge clk) O57_N2_S2 <=     O57_N4_S1  +  O57_N6_S1 ;
 logic signed [21:0] O57_N4_S2;		always @(posedge clk) O57_N4_S2 <=     O57_N8_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O57_N0_S3;		always @(posedge clk) O57_N0_S3 <=     O57_N0_S2  +  O57_N2_S2 ;
 logic signed [22:0] O57_N2_S3;		always @(posedge clk) O57_N2_S3 <=     O57_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O57_N0_S4;		always @(posedge clk) O57_N0_S4 <=     O57_N0_S3  +  O57_N2_S3 ;
 assign conv_mac_57 = O57_N0_S4;

logic signed [31:0] conv_mac_58;
logic signed [63:0] chainout_0_O58; 
logic signed [63:0] O58_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O58(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay(-9'sd1),.bx(input_fmap_2[7:0]),.by(-9'sd1),.cx(input_fmap_5[7:0]),.cy( 9'sd1),.dx(input_fmap_6[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O58_N0_S1),.chainout(chainout_0_O58));
logic signed [63:0] chainout_2_O58; 
logic signed [63:0] O58_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O58(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_11[7:0]),.ay( 9'sd1),.bx(input_fmap_12[7:0]),.by(-9'sd1),.cx(input_fmap_13[7:0]),.cy(-9'sd1),.dx(input_fmap_15[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O58_N2_S1),.chainout(chainout_2_O58));
logic signed [63:0] chainout_4_O58; 
logic signed [63:0] O58_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O58(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_19[7:0]),.ay( 9'sd1),.bx(input_fmap_20[7:0]),.by( 9'sd1),.cx(input_fmap_23[7:0]),.cy(-9'sd1),.dx(input_fmap_24[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O58_N4_S1),.chainout(chainout_4_O58));
logic signed [63:0] chainout_6_O58; 
logic signed [63:0] O58_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O58(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_27[7:0]),.ay(-9'sd1),.bx(input_fmap_28[7:0]),.by( 9'sd1),.cx(input_fmap_29[7:0]),.cy( 9'sd1),.dx(input_fmap_30[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O58_N6_S1),.chainout(chainout_6_O58));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O58_N0_S2;		always @(posedge clk) O58_N0_S2 <=     O58_N0_S1  +  O58_N2_S1 ;
 logic signed [21:0] O58_N2_S2;		always @(posedge clk) O58_N2_S2 <=     O58_N4_S1  +  O58_N6_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O58_N0_S3;		always @(posedge clk) O58_N0_S3 <=     O58_N0_S2  +  O58_N2_S2 ;
 assign conv_mac_58 = O58_N0_S3;

logic signed [31:0] conv_mac_59;
logic signed [63:0] chainout_0_O59; 
logic signed [63:0] O59_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O59(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay(-9'sd1),.bx(input_fmap_2[7:0]),.by( 9'sd1),.cx(input_fmap_3[7:0]),.cy(-9'sd1),.dx(input_fmap_4[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O59_N0_S1),.chainout(chainout_0_O59));
logic signed [63:0] chainout_2_O59; 
logic signed [63:0] O59_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O59(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_5[7:0]),.ay(-9'sd2),.bx(input_fmap_6[7:0]),.by( 9'sd4),.cx(input_fmap_10[7:0]),.cy(-9'sd1),.dx(input_fmap_11[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O59_N2_S1),.chainout(chainout_2_O59));
logic signed [63:0] chainout_4_O59; 
logic signed [63:0] O59_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O59(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_12[7:0]),.ay(-9'sd1),.bx(input_fmap_14[7:0]),.by( 9'sd1),.cx(input_fmap_16[7:0]),.cy(-9'sd1),.dx(input_fmap_18[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O59_N4_S1),.chainout(chainout_4_O59));
logic signed [63:0] chainout_6_O59; 
logic signed [63:0] O59_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O59(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_19[7:0]),.ay( 9'sd1),.bx(input_fmap_21[7:0]),.by(-9'sd1),.cx(input_fmap_23[7:0]),.cy(-9'sd1),.dx(input_fmap_24[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O59_N6_S1),.chainout(chainout_6_O59));
logic signed [63:0] chainout_8_O59; 
logic signed [63:0] O59_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O59(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_25[7:0]),.ay(-9'sd1),.bx(input_fmap_27[7:0]),.by( 9'sd2),.cx(input_fmap_28[7:0]),.cy( 9'sd2),.dx(input_fmap_29[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O59_N8_S1),.chainout(chainout_8_O59));
logic signed [63:0] chainout_10_O59; 
logic signed [63:0] O59_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O59(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_31[7:0]),.ay(-9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O59_N10_S1),.chainout(chainout_10_O59));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O59_N0_S2;		always @(posedge clk) O59_N0_S2 <=     O59_N0_S1  +  O59_N2_S1 ;
 logic signed [21:0] O59_N2_S2;		always @(posedge clk) O59_N2_S2 <=     O59_N4_S1  +  O59_N6_S1 ;
 logic signed [21:0] O59_N4_S2;		always @(posedge clk) O59_N4_S2 <=     O59_N8_S1  +  O59_N10_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O59_N0_S3;		always @(posedge clk) O59_N0_S3 <=     O59_N0_S2  +  O59_N2_S2 ;
 logic signed [22:0] O59_N2_S3;		always @(posedge clk) O59_N2_S3 <=     O59_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O59_N0_S4;		always @(posedge clk) O59_N0_S4 <=     O59_N0_S3  +  O59_N2_S3 ;
 assign conv_mac_59 = O59_N0_S4;

logic signed [31:0] conv_mac_60;
logic signed [63:0] chainout_0_O60; 
logic signed [63:0] O60_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O60(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_6[7:0]),.ay( 9'sd1),.bx(input_fmap_7[7:0]),.by( 9'sd1),.cx(input_fmap_9[7:0]),.cy(-9'sd1),.dx(input_fmap_12[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O60_N0_S1),.chainout(chainout_0_O60));
logic signed [63:0] chainout_2_O60; 
logic signed [63:0] O60_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O60(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_16[7:0]),.ay( 9'sd1),.bx(input_fmap_19[7:0]),.by( 9'sd1),.cx(input_fmap_20[7:0]),.cy(-9'sd1),.dx(input_fmap_21[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O60_N2_S1),.chainout(chainout_2_O60));
logic signed [63:0] chainout_4_O60; 
logic signed [63:0] O60_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O60(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_27[7:0]),.ay(-9'sd1),.bx(input_fmap_30[7:0]),.by( 9'sd3),.cx(input_fmap_31[7:0]),.cy( 9'sd2),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O60_N4_S1),.chainout(chainout_4_O60));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O60_N0_S2;		always @(posedge clk) O60_N0_S2 <=     O60_N0_S1  +  O60_N2_S1 ;
 logic signed [21:0] O60_N2_S2;		always @(posedge clk) O60_N2_S2 <=     O60_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O60_N0_S3;		always @(posedge clk) O60_N0_S3 <=     O60_N0_S2  +  O60_N2_S2 ;
 assign conv_mac_60 = O60_N0_S3;

logic signed [31:0] conv_mac_61;
logic signed [63:0] chainout_0_O61; 
logic signed [63:0] O61_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O61(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay(-9'sd1),.bx(input_fmap_10[7:0]),.by( 9'sd1),.cx(input_fmap_26[7:0]),.cy(-9'sd1),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O61_N0_S1),.chainout(chainout_0_O61));
assign conv_mac_61 = O61_N0_S1;

logic signed [31:0] conv_mac_62;
logic signed [63:0] chainout_0_O62; 
logic signed [63:0] O62_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O62(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd1),.bx(input_fmap_1[7:0]),.by( 9'sd1),.cx(input_fmap_4[7:0]),.cy(-9'sd2),.dx(input_fmap_6[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O62_N0_S1),.chainout(chainout_0_O62));
logic signed [63:0] chainout_2_O62; 
logic signed [63:0] O62_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O62(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_7[7:0]),.ay( 9'sd1),.bx(input_fmap_9[7:0]),.by( 9'sd4),.cx(input_fmap_10[7:0]),.cy(-9'sd2),.dx(input_fmap_11[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O62_N2_S1),.chainout(chainout_2_O62));
logic signed [63:0] chainout_4_O62; 
logic signed [63:0] O62_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O62(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_12[7:0]),.ay(-9'sd2),.bx(input_fmap_13[7:0]),.by( 9'sd1),.cx(input_fmap_14[7:0]),.cy( 9'sd1),.dx(input_fmap_16[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O62_N4_S1),.chainout(chainout_4_O62));
logic signed [63:0] chainout_6_O62; 
logic signed [63:0] O62_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O62(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_17[7:0]),.ay(-9'sd3),.bx(input_fmap_20[7:0]),.by( 9'sd1),.cx(input_fmap_22[7:0]),.cy(-9'sd1),.dx(input_fmap_24[7:0]),.dy(-9'sd3),.chainin(63'd0),.result(O62_N6_S1),.chainout(chainout_6_O62));
logic signed [63:0] chainout_8_O62; 
logic signed [63:0] O62_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O62(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_25[7:0]),.ay(-9'sd2),.bx(input_fmap_28[7:0]),.by(-9'sd1),.cx(input_fmap_31[7:0]),.cy( 9'sd5),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O62_N8_S1),.chainout(chainout_8_O62));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O62_N0_S2;		always @(posedge clk) O62_N0_S2 <=     O62_N0_S1  +  O62_N2_S1 ;
 logic signed [21:0] O62_N2_S2;		always @(posedge clk) O62_N2_S2 <=     O62_N4_S1  +  O62_N6_S1 ;
 logic signed [21:0] O62_N4_S2;		always @(posedge clk) O62_N4_S2 <=     O62_N8_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O62_N0_S3;		always @(posedge clk) O62_N0_S3 <=     O62_N0_S2  +  O62_N2_S2 ;
 logic signed [22:0] O62_N2_S3;		always @(posedge clk) O62_N2_S3 <=     O62_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O62_N0_S4;		always @(posedge clk) O62_N0_S4 <=     O62_N0_S3  +  O62_N2_S3 ;
 assign conv_mac_62 = O62_N0_S4;

logic signed [31:0] conv_mac_63;
logic signed [63:0] chainout_0_O63; 
logic signed [63:0] O63_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O63(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_12[7:0]),.ay(-9'sd1),.bx(input_fmap_13[7:0]),.by( 9'sd2),.cx(input_fmap_25[7:0]),.cy( 9'sd1),.dx(input_fmap_30[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O63_N0_S1),.chainout(chainout_0_O63));
assign conv_mac_63 = O63_N0_S1;

logic valid_D1;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D1<= 0 ;
	else valid_D1<=valid;
end
logic valid_D2;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D2<= 0 ;
	else valid_D2<=valid_D1;
end
logic valid_D3;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D3<= 0 ;
	else valid_D3<=valid_D2;
end
logic valid_D4;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D4<= 0 ;
	else valid_D4<=valid_D3;
end
logic valid_D5;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D5<= 0 ;
	else valid_D5<=valid_D4;
end
always_ff @(posedge clk) begin
	if (rstn == 0) ready <= 0 ;
	else ready <=valid_D5;
end
logic [31:0] bias_add_0;
assign bias_add_0 = conv_mac_0 + 6'd18;
logic [31:0] bias_add_1;
assign bias_add_1 = conv_mac_1 + 5'd8;
logic [31:0] bias_add_2;
assign bias_add_2 = conv_mac_2 + 6'd18;
logic [31:0] bias_add_3;
assign bias_add_3 = conv_mac_3 + 5'd11;
logic [31:0] bias_add_4;
assign bias_add_4 = conv_mac_4 + 5'd14;
logic [31:0] bias_add_5;
assign bias_add_5 = conv_mac_5 + 5'd14;
logic [31:0] bias_add_6;
assign bias_add_6 = conv_mac_6 + 6'd30;
logic [31:0] bias_add_7;
assign bias_add_7 = conv_mac_7 + 5'd14;
logic [31:0] bias_add_8;
assign bias_add_8 = conv_mac_8 + 6'd26;
logic [31:0] bias_add_9;
assign bias_add_9 = conv_mac_9 + 5'd13;
logic [31:0] bias_add_10;
assign bias_add_10 = conv_mac_10;
logic [31:0] bias_add_11;
assign bias_add_11 = conv_mac_11 + 4'd7;
logic [31:0] bias_add_12;
assign bias_add_12 = conv_mac_12 + 4'd4;
logic [31:0] bias_add_13;
assign bias_add_13 = conv_mac_13 + 5'd12;
logic [31:0] bias_add_14;
assign bias_add_14 = conv_mac_14 - 4'd4;
logic [31:0] bias_add_15;
assign bias_add_15 = conv_mac_15 - 3'd2;
logic [31:0] bias_add_16;
assign bias_add_16 = conv_mac_16 + 5'd8;
logic [31:0] bias_add_17;
assign bias_add_17 = conv_mac_17 + 6'd19;
logic [31:0] bias_add_18;
assign bias_add_18 = conv_mac_18 + 5'd13;
logic [31:0] bias_add_19;
assign bias_add_19 = conv_mac_19 + 5'd9;
logic [31:0] bias_add_20;
assign bias_add_20 = conv_mac_20 + 5'd11;
logic [31:0] bias_add_21;
assign bias_add_21 = conv_mac_21 + 6'd30;
logic [31:0] bias_add_22;
assign bias_add_22 = conv_mac_22 + 6'd17;
logic [31:0] bias_add_23;
assign bias_add_23 = conv_mac_23 + 2'd1;
logic [31:0] bias_add_24;
assign bias_add_24 = conv_mac_24 + 6'd17;
logic [31:0] bias_add_25;
assign bias_add_25 = conv_mac_25 + 6'd17;
logic [31:0] bias_add_26;
assign bias_add_26 = conv_mac_26 + 5'd14;
logic [31:0] bias_add_27;
assign bias_add_27 = conv_mac_27 + 5'd11;
logic [31:0] bias_add_28;
assign bias_add_28 = conv_mac_28 - 4'd6;
logic [31:0] bias_add_29;
assign bias_add_29 = conv_mac_29 + 6'd22;
logic [31:0] bias_add_30;
assign bias_add_30 = conv_mac_30 + 4'd6;
logic [31:0] bias_add_31;
assign bias_add_31 = conv_mac_31 + 6'd18;
logic [31:0] bias_add_32;
assign bias_add_32 = conv_mac_32 + 5'd12;
logic [31:0] bias_add_33;
assign bias_add_33 = conv_mac_33 + 6'd16;
logic [31:0] bias_add_34;
assign bias_add_34 = conv_mac_34 - 4'd5;
logic [31:0] bias_add_35;
assign bias_add_35 = conv_mac_35 + 6'd17;
logic [31:0] bias_add_36;
assign bias_add_36 = conv_mac_36 + 5'd14;
logic [31:0] bias_add_37;
assign bias_add_37 = conv_mac_37 + 5'd8;
logic [31:0] bias_add_38;
assign bias_add_38 = conv_mac_38 + 6'd18;
logic [31:0] bias_add_39;
assign bias_add_39 = conv_mac_39 + 4'd7;
logic [31:0] bias_add_40;
assign bias_add_40 = conv_mac_40 + 5'd10;
logic [31:0] bias_add_41;
assign bias_add_41 = conv_mac_41 + 6'd19;
logic [31:0] bias_add_42;
assign bias_add_42 = conv_mac_42 + 6'd16;
logic [31:0] bias_add_43;
assign bias_add_43 = conv_mac_43 + 6'd16;
logic [31:0] bias_add_44;
assign bias_add_44 = conv_mac_44 + 6'd24;
logic [31:0] bias_add_45;
assign bias_add_45 = conv_mac_45;
logic [31:0] bias_add_46;
assign bias_add_46 = conv_mac_46 + 5'd15;
logic [31:0] bias_add_47;
assign bias_add_47 = conv_mac_47 + 6'd16;
logic [31:0] bias_add_48;
assign bias_add_48 = conv_mac_48 + 5'd10;
logic [31:0] bias_add_49;
assign bias_add_49 = conv_mac_49 + 6'd22;
logic [31:0] bias_add_50;
assign bias_add_50 = conv_mac_50 + 7'd33;
logic [31:0] bias_add_51;
assign bias_add_51 = conv_mac_51 + 5'd10;
logic [31:0] bias_add_52;
assign bias_add_52 = conv_mac_52 + 5'd15;
logic [31:0] bias_add_53;
assign bias_add_53 = conv_mac_53 + 6'd22;
logic [31:0] bias_add_54;
assign bias_add_54 = conv_mac_54 - 4'd5;
logic [31:0] bias_add_55;
assign bias_add_55 = conv_mac_55 + 6'd17;
logic [31:0] bias_add_56;
assign bias_add_56 = conv_mac_56 + 5'd13;
logic [31:0] bias_add_57;
assign bias_add_57 = conv_mac_57 + 5'd10;
logic [31:0] bias_add_58;
assign bias_add_58 = conv_mac_58 + 5'd11;
logic [31:0] bias_add_59;
assign bias_add_59 = conv_mac_59 + 6'd16;
logic [31:0] bias_add_60;
assign bias_add_60 = conv_mac_60 + 4'd6;
logic [31:0] bias_add_61;
assign bias_add_61 = conv_mac_61 + 6'd20;
logic [31:0] bias_add_62;
assign bias_add_62 = conv_mac_62 + 2'd1;
logic [31:0] bias_add_63;
assign bias_add_63 = conv_mac_63 + 6'd19;

logic [7:0] relu_0;
assign relu_0[7:0] = (bias_add_0[31]==0) ? ((bias_add_0<3'd6) ? {{bias_add_0[31],bias_add_0[10:4]}} :'d6) : '0;
logic [7:0] relu_1;
assign relu_1[7:0] = (bias_add_1[31]==0) ? ((bias_add_1<3'd6) ? {{bias_add_1[31],bias_add_1[10:4]}} :'d6) : '0;
logic [7:0] relu_2;
assign relu_2[7:0] = (bias_add_2[31]==0) ? ((bias_add_2<3'd6) ? {{bias_add_2[31],bias_add_2[10:4]}} :'d6) : '0;
logic [7:0] relu_3;
assign relu_3[7:0] = (bias_add_3[31]==0) ? ((bias_add_3<3'd6) ? {{bias_add_3[31],bias_add_3[10:4]}} :'d6) : '0;
logic [7:0] relu_4;
assign relu_4[7:0] = (bias_add_4[31]==0) ? ((bias_add_4<3'd6) ? {{bias_add_4[31],bias_add_4[10:4]}} :'d6) : '0;
logic [7:0] relu_5;
assign relu_5[7:0] = (bias_add_5[31]==0) ? ((bias_add_5<3'd6) ? {{bias_add_5[31],bias_add_5[10:4]}} :'d6) : '0;
logic [7:0] relu_6;
assign relu_6[7:0] = (bias_add_6[31]==0) ? ((bias_add_6<3'd6) ? {{bias_add_6[31],bias_add_6[10:4]}} :'d6) : '0;
logic [7:0] relu_7;
assign relu_7[7:0] = (bias_add_7[31]==0) ? ((bias_add_7<3'd6) ? {{bias_add_7[31],bias_add_7[10:4]}} :'d6) : '0;
logic [7:0] relu_8;
assign relu_8[7:0] = (bias_add_8[31]==0) ? ((bias_add_8<3'd6) ? {{bias_add_8[31],bias_add_8[10:4]}} :'d6) : '0;
logic [7:0] relu_9;
assign relu_9[7:0] = (bias_add_9[31]==0) ? ((bias_add_9<3'd6) ? {{bias_add_9[31],bias_add_9[10:4]}} :'d6) : '0;
logic [7:0] relu_10;
assign relu_10[7:0] = (bias_add_10[31]==0) ? ((bias_add_10<3'd6) ? {{bias_add_10[31],bias_add_10[10:4]}} :'d6) : '0;
logic [7:0] relu_11;
assign relu_11[7:0] = (bias_add_11[31]==0) ? ((bias_add_11<3'd6) ? {{bias_add_11[31],bias_add_11[10:4]}} :'d6) : '0;
logic [7:0] relu_12;
assign relu_12[7:0] = (bias_add_12[31]==0) ? ((bias_add_12<3'd6) ? {{bias_add_12[31],bias_add_12[10:4]}} :'d6) : '0;
logic [7:0] relu_13;
assign relu_13[7:0] = (bias_add_13[31]==0) ? ((bias_add_13<3'd6) ? {{bias_add_13[31],bias_add_13[10:4]}} :'d6) : '0;
logic [7:0] relu_14;
assign relu_14[7:0] = (bias_add_14[31]==0) ? ((bias_add_14<3'd6) ? {{bias_add_14[31],bias_add_14[10:4]}} :'d6) : '0;
logic [7:0] relu_15;
assign relu_15[7:0] = (bias_add_15[31]==0) ? ((bias_add_15<3'd6) ? {{bias_add_15[31],bias_add_15[10:4]}} :'d6) : '0;
logic [7:0] relu_16;
assign relu_16[7:0] = (bias_add_16[31]==0) ? ((bias_add_16<3'd6) ? {{bias_add_16[31],bias_add_16[10:4]}} :'d6) : '0;
logic [7:0] relu_17;
assign relu_17[7:0] = (bias_add_17[31]==0) ? ((bias_add_17<3'd6) ? {{bias_add_17[31],bias_add_17[10:4]}} :'d6) : '0;
logic [7:0] relu_18;
assign relu_18[7:0] = (bias_add_18[31]==0) ? ((bias_add_18<3'd6) ? {{bias_add_18[31],bias_add_18[10:4]}} :'d6) : '0;
logic [7:0] relu_19;
assign relu_19[7:0] = (bias_add_19[31]==0) ? ((bias_add_19<3'd6) ? {{bias_add_19[31],bias_add_19[10:4]}} :'d6) : '0;
logic [7:0] relu_20;
assign relu_20[7:0] = (bias_add_20[31]==0) ? ((bias_add_20<3'd6) ? {{bias_add_20[31],bias_add_20[10:4]}} :'d6) : '0;
logic [7:0] relu_21;
assign relu_21[7:0] = (bias_add_21[31]==0) ? ((bias_add_21<3'd6) ? {{bias_add_21[31],bias_add_21[10:4]}} :'d6) : '0;
logic [7:0] relu_22;
assign relu_22[7:0] = (bias_add_22[31]==0) ? ((bias_add_22<3'd6) ? {{bias_add_22[31],bias_add_22[10:4]}} :'d6) : '0;
logic [7:0] relu_23;
assign relu_23[7:0] = (bias_add_23[31]==0) ? ((bias_add_23<3'd6) ? {{bias_add_23[31],bias_add_23[10:4]}} :'d6) : '0;
logic [7:0] relu_24;
assign relu_24[7:0] = (bias_add_24[31]==0) ? ((bias_add_24<3'd6) ? {{bias_add_24[31],bias_add_24[10:4]}} :'d6) : '0;
logic [7:0] relu_25;
assign relu_25[7:0] = (bias_add_25[31]==0) ? ((bias_add_25<3'd6) ? {{bias_add_25[31],bias_add_25[10:4]}} :'d6) : '0;
logic [7:0] relu_26;
assign relu_26[7:0] = (bias_add_26[31]==0) ? ((bias_add_26<3'd6) ? {{bias_add_26[31],bias_add_26[10:4]}} :'d6) : '0;
logic [7:0] relu_27;
assign relu_27[7:0] = (bias_add_27[31]==0) ? ((bias_add_27<3'd6) ? {{bias_add_27[31],bias_add_27[10:4]}} :'d6) : '0;
logic [7:0] relu_28;
assign relu_28[7:0] = (bias_add_28[31]==0) ? ((bias_add_28<3'd6) ? {{bias_add_28[31],bias_add_28[10:4]}} :'d6) : '0;
logic [7:0] relu_29;
assign relu_29[7:0] = (bias_add_29[31]==0) ? ((bias_add_29<3'd6) ? {{bias_add_29[31],bias_add_29[10:4]}} :'d6) : '0;
logic [7:0] relu_30;
assign relu_30[7:0] = (bias_add_30[31]==0) ? ((bias_add_30<3'd6) ? {{bias_add_30[31],bias_add_30[10:4]}} :'d6) : '0;
logic [7:0] relu_31;
assign relu_31[7:0] = (bias_add_31[31]==0) ? ((bias_add_31<3'd6) ? {{bias_add_31[31],bias_add_31[10:4]}} :'d6) : '0;
logic [7:0] relu_32;
assign relu_32[7:0] = (bias_add_32[31]==0) ? ((bias_add_32<3'd6) ? {{bias_add_32[31],bias_add_32[10:4]}} :'d6) : '0;
logic [7:0] relu_33;
assign relu_33[7:0] = (bias_add_33[31]==0) ? ((bias_add_33<3'd6) ? {{bias_add_33[31],bias_add_33[10:4]}} :'d6) : '0;
logic [7:0] relu_34;
assign relu_34[7:0] = (bias_add_34[31]==0) ? ((bias_add_34<3'd6) ? {{bias_add_34[31],bias_add_34[10:4]}} :'d6) : '0;
logic [7:0] relu_35;
assign relu_35[7:0] = (bias_add_35[31]==0) ? ((bias_add_35<3'd6) ? {{bias_add_35[31],bias_add_35[10:4]}} :'d6) : '0;
logic [7:0] relu_36;
assign relu_36[7:0] = (bias_add_36[31]==0) ? ((bias_add_36<3'd6) ? {{bias_add_36[31],bias_add_36[10:4]}} :'d6) : '0;
logic [7:0] relu_37;
assign relu_37[7:0] = (bias_add_37[31]==0) ? ((bias_add_37<3'd6) ? {{bias_add_37[31],bias_add_37[10:4]}} :'d6) : '0;
logic [7:0] relu_38;
assign relu_38[7:0] = (bias_add_38[31]==0) ? ((bias_add_38<3'd6) ? {{bias_add_38[31],bias_add_38[10:4]}} :'d6) : '0;
logic [7:0] relu_39;
assign relu_39[7:0] = (bias_add_39[31]==0) ? ((bias_add_39<3'd6) ? {{bias_add_39[31],bias_add_39[10:4]}} :'d6) : '0;
logic [7:0] relu_40;
assign relu_40[7:0] = (bias_add_40[31]==0) ? ((bias_add_40<3'd6) ? {{bias_add_40[31],bias_add_40[10:4]}} :'d6) : '0;
logic [7:0] relu_41;
assign relu_41[7:0] = (bias_add_41[31]==0) ? ((bias_add_41<3'd6) ? {{bias_add_41[31],bias_add_41[10:4]}} :'d6) : '0;
logic [7:0] relu_42;
assign relu_42[7:0] = (bias_add_42[31]==0) ? ((bias_add_42<3'd6) ? {{bias_add_42[31],bias_add_42[10:4]}} :'d6) : '0;
logic [7:0] relu_43;
assign relu_43[7:0] = (bias_add_43[31]==0) ? ((bias_add_43<3'd6) ? {{bias_add_43[31],bias_add_43[10:4]}} :'d6) : '0;
logic [7:0] relu_44;
assign relu_44[7:0] = (bias_add_44[31]==0) ? ((bias_add_44<3'd6) ? {{bias_add_44[31],bias_add_44[10:4]}} :'d6) : '0;
logic [7:0] relu_45;
assign relu_45[7:0] = (bias_add_45[31]==0) ? ((bias_add_45<3'd6) ? {{bias_add_45[31],bias_add_45[10:4]}} :'d6) : '0;
logic [7:0] relu_46;
assign relu_46[7:0] = (bias_add_46[31]==0) ? ((bias_add_46<3'd6) ? {{bias_add_46[31],bias_add_46[10:4]}} :'d6) : '0;
logic [7:0] relu_47;
assign relu_47[7:0] = (bias_add_47[31]==0) ? ((bias_add_47<3'd6) ? {{bias_add_47[31],bias_add_47[10:4]}} :'d6) : '0;
logic [7:0] relu_48;
assign relu_48[7:0] = (bias_add_48[31]==0) ? ((bias_add_48<3'd6) ? {{bias_add_48[31],bias_add_48[10:4]}} :'d6) : '0;
logic [7:0] relu_49;
assign relu_49[7:0] = (bias_add_49[31]==0) ? ((bias_add_49<3'd6) ? {{bias_add_49[31],bias_add_49[10:4]}} :'d6) : '0;
logic [7:0] relu_50;
assign relu_50[7:0] = (bias_add_50[31]==0) ? ((bias_add_50<3'd6) ? {{bias_add_50[31],bias_add_50[10:4]}} :'d6) : '0;
logic [7:0] relu_51;
assign relu_51[7:0] = (bias_add_51[31]==0) ? ((bias_add_51<3'd6) ? {{bias_add_51[31],bias_add_51[10:4]}} :'d6) : '0;
logic [7:0] relu_52;
assign relu_52[7:0] = (bias_add_52[31]==0) ? ((bias_add_52<3'd6) ? {{bias_add_52[31],bias_add_52[10:4]}} :'d6) : '0;
logic [7:0] relu_53;
assign relu_53[7:0] = (bias_add_53[31]==0) ? ((bias_add_53<3'd6) ? {{bias_add_53[31],bias_add_53[10:4]}} :'d6) : '0;
logic [7:0] relu_54;
assign relu_54[7:0] = (bias_add_54[31]==0) ? ((bias_add_54<3'd6) ? {{bias_add_54[31],bias_add_54[10:4]}} :'d6) : '0;
logic [7:0] relu_55;
assign relu_55[7:0] = (bias_add_55[31]==0) ? ((bias_add_55<3'd6) ? {{bias_add_55[31],bias_add_55[10:4]}} :'d6) : '0;
logic [7:0] relu_56;
assign relu_56[7:0] = (bias_add_56[31]==0) ? ((bias_add_56<3'd6) ? {{bias_add_56[31],bias_add_56[10:4]}} :'d6) : '0;
logic [7:0] relu_57;
assign relu_57[7:0] = (bias_add_57[31]==0) ? ((bias_add_57<3'd6) ? {{bias_add_57[31],bias_add_57[10:4]}} :'d6) : '0;
logic [7:0] relu_58;
assign relu_58[7:0] = (bias_add_58[31]==0) ? ((bias_add_58<3'd6) ? {{bias_add_58[31],bias_add_58[10:4]}} :'d6) : '0;
logic [7:0] relu_59;
assign relu_59[7:0] = (bias_add_59[31]==0) ? ((bias_add_59<3'd6) ? {{bias_add_59[31],bias_add_59[10:4]}} :'d6) : '0;
logic [7:0] relu_60;
assign relu_60[7:0] = (bias_add_60[31]==0) ? ((bias_add_60<3'd6) ? {{bias_add_60[31],bias_add_60[10:4]}} :'d6) : '0;
logic [7:0] relu_61;
assign relu_61[7:0] = (bias_add_61[31]==0) ? ((bias_add_61<3'd6) ? {{bias_add_61[31],bias_add_61[10:4]}} :'d6) : '0;
logic [7:0] relu_62;
assign relu_62[7:0] = (bias_add_62[31]==0) ? ((bias_add_62<3'd6) ? {{bias_add_62[31],bias_add_62[10:4]}} :'d6) : '0;
logic [7:0] relu_63;
assign relu_63[7:0] = (bias_add_63[31]==0) ? ((bias_add_63<3'd6) ? {{bias_add_63[31],bias_add_63[10:4]}} :'d6) : '0;

assign output_act = {
	relu_63,
	relu_62,
	relu_61,
	relu_60,
	relu_59,
	relu_58,
	relu_57,
	relu_56,
	relu_55,
	relu_54,
	relu_53,
	relu_52,
	relu_51,
	relu_50,
	relu_49,
	relu_48,
	relu_47,
	relu_46,
	relu_45,
	relu_44,
	relu_43,
	relu_42,
	relu_41,
	relu_40,
	relu_39,
	relu_38,
	relu_37,
	relu_36,
	relu_35,
	relu_34,
	relu_33,
	relu_32,
	relu_31,
	relu_30,
	relu_29,
	relu_28,
	relu_27,
	relu_26,
	relu_25,
	relu_24,
	relu_23,
	relu_22,
	relu_21,
	relu_20,
	relu_19,
	relu_18,
	relu_17,
	relu_16,
	relu_15,
	relu_14,
	relu_13,
	relu_12,
	relu_11,
	relu_10,
	relu_9,
	relu_8,
	relu_7,
	relu_6,
	relu_5,
	relu_4,
	relu_3,
	relu_2,
	relu_1,
	relu_0
};

endmodule
module conv7_pw (
    input logic clk,
    input logic rstn,
    input logic valid,
    input logic [512-1:0] input_act,
    output logic [512-1:0] output_act,
    output logic ready
);
logic we;
logic [8:0] zero_number; 
assign zero_number = 9'd0; 
//1
logic [512-1:0] input_act_ff ;
always_ff @(posedge clk) begin
    if (rstn == 0) begin
        input_act_ff <= '0;
      //  ready <= '0;
    end
    else begin
        input_act_ff <= input_act;
     //   ready <= valid;
    end
end
logic [7:0] input_fmap_0;
assign input_fmap_0 = input_act_ff[7:0];
logic [7:0] input_fmap_1;
assign input_fmap_1 = input_act_ff[15:8];
logic [7:0] input_fmap_2;
assign input_fmap_2 = input_act_ff[23:16];
logic [7:0] input_fmap_3;
assign input_fmap_3 = input_act_ff[31:24];
logic [7:0] input_fmap_4;
assign input_fmap_4 = input_act_ff[39:32];
logic [7:0] input_fmap_5;
assign input_fmap_5 = input_act_ff[47:40];
logic [7:0] input_fmap_6;
assign input_fmap_6 = input_act_ff[55:48];
logic [7:0] input_fmap_7;
assign input_fmap_7 = input_act_ff[63:56];
logic [7:0] input_fmap_8;
assign input_fmap_8 = input_act_ff[71:64];
logic [7:0] input_fmap_9;
assign input_fmap_9 = input_act_ff[79:72];
logic [7:0] input_fmap_10;
assign input_fmap_10 = input_act_ff[87:80];
logic [7:0] input_fmap_11;
assign input_fmap_11 = input_act_ff[95:88];
logic [7:0] input_fmap_12;
assign input_fmap_12 = input_act_ff[103:96];
logic [7:0] input_fmap_13;
assign input_fmap_13 = input_act_ff[111:104];
logic [7:0] input_fmap_14;
assign input_fmap_14 = input_act_ff[119:112];
logic [7:0] input_fmap_15;
assign input_fmap_15 = input_act_ff[127:120];
logic [7:0] input_fmap_16;
assign input_fmap_16 = input_act_ff[135:128];
logic [7:0] input_fmap_17;
assign input_fmap_17 = input_act_ff[143:136];
logic [7:0] input_fmap_18;
assign input_fmap_18 = input_act_ff[151:144];
logic [7:0] input_fmap_19;
assign input_fmap_19 = input_act_ff[159:152];
logic [7:0] input_fmap_20;
assign input_fmap_20 = input_act_ff[167:160];
logic [7:0] input_fmap_21;
assign input_fmap_21 = input_act_ff[175:168];
logic [7:0] input_fmap_22;
assign input_fmap_22 = input_act_ff[183:176];
logic [7:0] input_fmap_23;
assign input_fmap_23 = input_act_ff[191:184];
logic [7:0] input_fmap_24;
assign input_fmap_24 = input_act_ff[199:192];
logic [7:0] input_fmap_25;
assign input_fmap_25 = input_act_ff[207:200];
logic [7:0] input_fmap_26;
assign input_fmap_26 = input_act_ff[215:208];
logic [7:0] input_fmap_27;
assign input_fmap_27 = input_act_ff[223:216];
logic [7:0] input_fmap_28;
assign input_fmap_28 = input_act_ff[231:224];
logic [7:0] input_fmap_29;
assign input_fmap_29 = input_act_ff[239:232];
logic [7:0] input_fmap_30;
assign input_fmap_30 = input_act_ff[247:240];
logic [7:0] input_fmap_31;
assign input_fmap_31 = input_act_ff[255:248];
logic [7:0] input_fmap_32;
assign input_fmap_32 = input_act_ff[263:256];
logic [7:0] input_fmap_33;
assign input_fmap_33 = input_act_ff[271:264];
logic [7:0] input_fmap_34;
assign input_fmap_34 = input_act_ff[279:272];
logic [7:0] input_fmap_35;
assign input_fmap_35 = input_act_ff[287:280];
logic [7:0] input_fmap_36;
assign input_fmap_36 = input_act_ff[295:288];
logic [7:0] input_fmap_37;
assign input_fmap_37 = input_act_ff[303:296];
logic [7:0] input_fmap_38;
assign input_fmap_38 = input_act_ff[311:304];
logic [7:0] input_fmap_39;
assign input_fmap_39 = input_act_ff[319:312];
logic [7:0] input_fmap_40;
assign input_fmap_40 = input_act_ff[327:320];
logic [7:0] input_fmap_41;
assign input_fmap_41 = input_act_ff[335:328];
logic [7:0] input_fmap_42;
assign input_fmap_42 = input_act_ff[343:336];
logic [7:0] input_fmap_43;
assign input_fmap_43 = input_act_ff[351:344];
logic [7:0] input_fmap_44;
assign input_fmap_44 = input_act_ff[359:352];
logic [7:0] input_fmap_45;
assign input_fmap_45 = input_act_ff[367:360];
logic [7:0] input_fmap_46;
assign input_fmap_46 = input_act_ff[375:368];
logic [7:0] input_fmap_47;
assign input_fmap_47 = input_act_ff[383:376];
logic [7:0] input_fmap_48;
assign input_fmap_48 = input_act_ff[391:384];
logic [7:0] input_fmap_49;
assign input_fmap_49 = input_act_ff[399:392];
logic [7:0] input_fmap_50;
assign input_fmap_50 = input_act_ff[407:400];
logic [7:0] input_fmap_51;
assign input_fmap_51 = input_act_ff[415:408];
logic [7:0] input_fmap_52;
assign input_fmap_52 = input_act_ff[423:416];
logic [7:0] input_fmap_53;
assign input_fmap_53 = input_act_ff[431:424];
logic [7:0] input_fmap_54;
assign input_fmap_54 = input_act_ff[439:432];
logic [7:0] input_fmap_55;
assign input_fmap_55 = input_act_ff[447:440];
logic [7:0] input_fmap_56;
assign input_fmap_56 = input_act_ff[455:448];
logic [7:0] input_fmap_57;
assign input_fmap_57 = input_act_ff[463:456];
logic [7:0] input_fmap_58;
assign input_fmap_58 = input_act_ff[471:464];
logic [7:0] input_fmap_59;
assign input_fmap_59 = input_act_ff[479:472];
logic [7:0] input_fmap_60;
assign input_fmap_60 = input_act_ff[487:480];
logic [7:0] input_fmap_61;
assign input_fmap_61 = input_act_ff[495:488];
logic [7:0] input_fmap_62;
assign input_fmap_62 = input_act_ff[503:496];
logic [7:0] input_fmap_63;
assign input_fmap_63 = input_act_ff[511:504];

logic signed [31:0] conv_mac_0;
logic signed [63:0] chainout_0_O0; 
logic signed [63:0] O0_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O0(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd1),.bx(input_fmap_2[7:0]),.by(-9'sd1),.cx(input_fmap_4[7:0]),.cy(-9'sd1),.dx(input_fmap_5[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O0_N0_S1),.chainout(chainout_0_O0));
logic signed [63:0] chainout_2_O0; 
logic signed [63:0] O0_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O0(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_6[7:0]),.ay(-9'sd1),.bx(input_fmap_7[7:0]),.by( 9'sd1),.cx(input_fmap_10[7:0]),.cy(-9'sd1),.dx(input_fmap_11[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O0_N2_S1),.chainout(chainout_2_O0));
logic signed [63:0] chainout_4_O0; 
logic signed [63:0] O0_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O0(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_12[7:0]),.ay( 9'sd1),.bx(input_fmap_13[7:0]),.by(-9'sd1),.cx(input_fmap_14[7:0]),.cy( 9'sd1),.dx(input_fmap_15[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O0_N4_S1),.chainout(chainout_4_O0));
logic signed [63:0] chainout_6_O0; 
logic signed [63:0] O0_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O0(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_16[7:0]),.ay( 9'sd1),.bx(input_fmap_17[7:0]),.by(-9'sd1),.cx(input_fmap_19[7:0]),.cy( 9'sd1),.dx(input_fmap_22[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O0_N6_S1),.chainout(chainout_6_O0));
logic signed [63:0] chainout_8_O0; 
logic signed [63:0] O0_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O0(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_23[7:0]),.ay(-9'sd1),.bx(input_fmap_24[7:0]),.by(-9'sd1),.cx(input_fmap_25[7:0]),.cy(-9'sd2),.dx(input_fmap_27[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O0_N8_S1),.chainout(chainout_8_O0));
logic signed [63:0] chainout_10_O0; 
logic signed [63:0] O0_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O0(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_30[7:0]),.ay(-9'sd1),.bx(input_fmap_31[7:0]),.by( 9'sd1),.cx(input_fmap_33[7:0]),.cy(-9'sd1),.dx(input_fmap_34[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O0_N10_S1),.chainout(chainout_10_O0));
logic signed [63:0] chainout_12_O0; 
logic signed [63:0] O0_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O0(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_39[7:0]),.ay(-9'sd1),.bx(input_fmap_40[7:0]),.by(-9'sd1),.cx(input_fmap_42[7:0]),.cy( 9'sd1),.dx(input_fmap_43[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O0_N12_S1),.chainout(chainout_12_O0));
logic signed [63:0] chainout_14_O0; 
logic signed [63:0] O0_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O0(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_44[7:0]),.ay(-9'sd2),.bx(input_fmap_45[7:0]),.by(-9'sd1),.cx(input_fmap_46[7:0]),.cy( 9'sd4),.dx(input_fmap_47[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O0_N14_S1),.chainout(chainout_14_O0));
logic signed [63:0] chainout_16_O0; 
logic signed [63:0] O0_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O0(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_49[7:0]),.ay( 9'sd1),.bx(input_fmap_50[7:0]),.by( 9'sd1),.cx(input_fmap_51[7:0]),.cy(-9'sd1),.dx(input_fmap_52[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O0_N16_S1),.chainout(chainout_16_O0));
logic signed [63:0] chainout_18_O0; 
logic signed [63:0] O0_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O0(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_55[7:0]),.ay(-9'sd1),.bx(input_fmap_56[7:0]),.by(-9'sd1),.cx(input_fmap_58[7:0]),.cy( 9'sd1),.dx(input_fmap_60[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O0_N18_S1),.chainout(chainout_18_O0));
logic signed [63:0] chainout_20_O0; 
logic signed [63:0] O0_N20_S1; 
 int_sop_4_wrapper int_sop_4_inst_20_O0(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_61[7:0]),.ay( 9'sd1),.bx(input_fmap_62[7:0]),.by( 9'sd2),.cx(input_fmap_63[7:0]),.cy(-9'sd2),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O0_N20_S1),.chainout(chainout_20_O0));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O0_N0_S2;		always @(posedge clk) O0_N0_S2 <=     O0_N0_S1  +  O0_N2_S1 ;
 logic signed [21:0] O0_N2_S2;		always @(posedge clk) O0_N2_S2 <=     O0_N4_S1  +  O0_N6_S1 ;
 logic signed [21:0] O0_N4_S2;		always @(posedge clk) O0_N4_S2 <=     O0_N8_S1  +  O0_N10_S1 ;
 logic signed [21:0] O0_N6_S2;		always @(posedge clk) O0_N6_S2 <=     O0_N12_S1  +  O0_N14_S1 ;
 logic signed [21:0] O0_N8_S2;		always @(posedge clk) O0_N8_S2 <=     O0_N16_S1  +  O0_N18_S1 ;
 logic signed [21:0] O0_N10_S2;		always @(posedge clk) O0_N10_S2 <=     O0_N20_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O0_N0_S3;		always @(posedge clk) O0_N0_S3 <=     O0_N0_S2  +  O0_N2_S2 ;
 logic signed [22:0] O0_N2_S3;		always @(posedge clk) O0_N2_S3 <=     O0_N4_S2  +  O0_N6_S2 ;
 logic signed [22:0] O0_N4_S3;		always @(posedge clk) O0_N4_S3 <=     O0_N8_S2  +  O0_N10_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O0_N0_S4;		always @(posedge clk) O0_N0_S4 <=     O0_N0_S3  +  O0_N2_S3 ;
 logic signed [23:0] O0_N2_S4;		always @(posedge clk) O0_N2_S4 <=     O0_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O0_N0_S5;		always @(posedge clk) O0_N0_S5 <=     O0_N0_S4  +  O0_N2_S4 ;
 assign conv_mac_0 = O0_N0_S5;

logic signed [31:0] conv_mac_1;
logic signed [63:0] chainout_0_O1; 
logic signed [63:0] O1_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O1(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_3[7:0]),.ay( 9'sd1),.bx(input_fmap_4[7:0]),.by( 9'sd1),.cx(input_fmap_7[7:0]),.cy( 9'sd1),.dx(input_fmap_12[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O1_N0_S1),.chainout(chainout_0_O1));
logic signed [63:0] chainout_2_O1; 
logic signed [63:0] O1_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O1(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_13[7:0]),.ay(-9'sd1),.bx(input_fmap_16[7:0]),.by(-9'sd1),.cx(input_fmap_17[7:0]),.cy(-9'sd1),.dx(input_fmap_18[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O1_N2_S1),.chainout(chainout_2_O1));
logic signed [63:0] chainout_4_O1; 
logic signed [63:0] O1_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O1(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_19[7:0]),.ay(-9'sd1),.bx(input_fmap_20[7:0]),.by( 9'sd1),.cx(input_fmap_21[7:0]),.cy(-9'sd1),.dx(input_fmap_22[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O1_N4_S1),.chainout(chainout_4_O1));
logic signed [63:0] chainout_6_O1; 
logic signed [63:0] O1_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O1(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_23[7:0]),.ay(-9'sd1),.bx(input_fmap_25[7:0]),.by(-9'sd1),.cx(input_fmap_26[7:0]),.cy( 9'sd1),.dx(input_fmap_27[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O1_N6_S1),.chainout(chainout_6_O1));
logic signed [63:0] chainout_8_O1; 
logic signed [63:0] O1_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O1(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_28[7:0]),.ay( 9'sd1),.bx(input_fmap_29[7:0]),.by(-9'sd1),.cx(input_fmap_31[7:0]),.cy(-9'sd1),.dx(input_fmap_33[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O1_N8_S1),.chainout(chainout_8_O1));
logic signed [63:0] chainout_10_O1; 
logic signed [63:0] O1_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O1(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_34[7:0]),.ay(-9'sd1),.bx(input_fmap_35[7:0]),.by( 9'sd1),.cx(input_fmap_39[7:0]),.cy(-9'sd1),.dx(input_fmap_41[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O1_N10_S1),.chainout(chainout_10_O1));
logic signed [63:0] chainout_12_O1; 
logic signed [63:0] O1_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O1(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_43[7:0]),.ay( 9'sd1),.bx(input_fmap_45[7:0]),.by(-9'sd1),.cx(input_fmap_46[7:0]),.cy(-9'sd2),.dx(input_fmap_47[7:0]),.dy( 9'sd3),.chainin(63'd0),.result(O1_N12_S1),.chainout(chainout_12_O1));
logic signed [63:0] chainout_14_O1; 
logic signed [63:0] O1_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O1(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_48[7:0]),.ay(-9'sd1),.bx(input_fmap_49[7:0]),.by( 9'sd1),.cx(input_fmap_50[7:0]),.cy(-9'sd1),.dx(input_fmap_51[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O1_N14_S1),.chainout(chainout_14_O1));
logic signed [63:0] chainout_16_O1; 
logic signed [63:0] O1_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O1(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_52[7:0]),.ay(-9'sd1),.bx(input_fmap_54[7:0]),.by(-9'sd1),.cx(input_fmap_56[7:0]),.cy(-9'sd1),.dx(input_fmap_57[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O1_N16_S1),.chainout(chainout_16_O1));
logic signed [63:0] chainout_18_O1; 
logic signed [63:0] O1_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O1(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_59[7:0]),.ay(-9'sd1),.bx(input_fmap_61[7:0]),.by( 9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O1_N18_S1),.chainout(chainout_18_O1));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O1_N0_S2;		always @(posedge clk) O1_N0_S2 <=     O1_N0_S1  +  O1_N2_S1 ;
 logic signed [21:0] O1_N2_S2;		always @(posedge clk) O1_N2_S2 <=     O1_N4_S1  +  O1_N6_S1 ;
 logic signed [21:0] O1_N4_S2;		always @(posedge clk) O1_N4_S2 <=     O1_N8_S1  +  O1_N10_S1 ;
 logic signed [21:0] O1_N6_S2;		always @(posedge clk) O1_N6_S2 <=     O1_N12_S1  +  O1_N14_S1 ;
 logic signed [21:0] O1_N8_S2;		always @(posedge clk) O1_N8_S2 <=     O1_N16_S1  +  O1_N18_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O1_N0_S3;		always @(posedge clk) O1_N0_S3 <=     O1_N0_S2  +  O1_N2_S2 ;
 logic signed [22:0] O1_N2_S3;		always @(posedge clk) O1_N2_S3 <=     O1_N4_S2  +  O1_N6_S2 ;
 logic signed [22:0] O1_N4_S3;		always @(posedge clk) O1_N4_S3 <=     O1_N8_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O1_N0_S4;		always @(posedge clk) O1_N0_S4 <=     O1_N0_S3  +  O1_N2_S3 ;
 logic signed [23:0] O1_N2_S4;		always @(posedge clk) O1_N2_S4 <=     O1_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O1_N0_S5;		always @(posedge clk) O1_N0_S5 <=     O1_N0_S4  +  O1_N2_S4 ;
 assign conv_mac_1 = O1_N0_S5;

logic signed [31:0] conv_mac_2;
logic signed [63:0] chainout_0_O2; 
logic signed [63:0] O2_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O2(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_9[7:0]),.ay( 9'sd1),.bx(input_fmap_16[7:0]),.by( 9'sd1),.cx(input_fmap_25[7:0]),.cy( 9'sd1),.dx(input_fmap_26[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O2_N0_S1),.chainout(chainout_0_O2));
logic signed [63:0] chainout_2_O2; 
logic signed [63:0] O2_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O2(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_33[7:0]),.ay( 9'sd1),.bx(input_fmap_39[7:0]),.by( 9'sd1),.cx(input_fmap_40[7:0]),.cy( 9'sd1),.dx(input_fmap_45[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O2_N2_S1),.chainout(chainout_2_O2));
logic signed [63:0] chainout_4_O2; 
logic signed [63:0] O2_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O2(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_50[7:0]),.ay( 9'sd1),.bx(input_fmap_54[7:0]),.by( 9'sd1),.cx(input_fmap_60[7:0]),.cy( 9'sd1),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O2_N4_S1),.chainout(chainout_4_O2));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O2_N0_S2;		always @(posedge clk) O2_N0_S2 <=     O2_N0_S1  +  O2_N2_S1 ;
 logic signed [21:0] O2_N2_S2;		always @(posedge clk) O2_N2_S2 <=     O2_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O2_N0_S3;		always @(posedge clk) O2_N0_S3 <=     O2_N0_S2  +  O2_N2_S2 ;
 assign conv_mac_2 = O2_N0_S3;

logic signed [31:0] conv_mac_3;
logic signed [63:0] chainout_0_O3; 
logic signed [63:0] O3_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O3(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_4[7:0]),.ay(-9'sd1),.bx(input_fmap_5[7:0]),.by( 9'sd1),.cx(input_fmap_7[7:0]),.cy(-9'sd1),.dx(input_fmap_9[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O3_N0_S1),.chainout(chainout_0_O3));
logic signed [63:0] chainout_2_O3; 
logic signed [63:0] O3_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O3(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_10[7:0]),.ay(-9'sd1),.bx(input_fmap_12[7:0]),.by( 9'sd1),.cx(input_fmap_13[7:0]),.cy( 9'sd2),.dx(input_fmap_14[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O3_N2_S1),.chainout(chainout_2_O3));
logic signed [63:0] chainout_4_O3; 
logic signed [63:0] O3_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O3(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_16[7:0]),.ay( 9'sd2),.bx(input_fmap_17[7:0]),.by(-9'sd2),.cx(input_fmap_20[7:0]),.cy(-9'sd1),.dx(input_fmap_21[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O3_N4_S1),.chainout(chainout_4_O3));
logic signed [63:0] chainout_6_O3; 
logic signed [63:0] O3_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O3(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_22[7:0]),.ay( 9'sd1),.bx(input_fmap_30[7:0]),.by(-9'sd1),.cx(input_fmap_31[7:0]),.cy(-9'sd1),.dx(input_fmap_32[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O3_N6_S1),.chainout(chainout_6_O3));
logic signed [63:0] chainout_8_O3; 
logic signed [63:0] O3_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O3(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_34[7:0]),.ay(-9'sd1),.bx(input_fmap_35[7:0]),.by( 9'sd1),.cx(input_fmap_36[7:0]),.cy(-9'sd1),.dx(input_fmap_37[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O3_N8_S1),.chainout(chainout_8_O3));
logic signed [63:0] chainout_10_O3; 
logic signed [63:0] O3_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O3(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_38[7:0]),.ay(-9'sd1),.bx(input_fmap_40[7:0]),.by( 9'sd1),.cx(input_fmap_41[7:0]),.cy(-9'sd1),.dx(input_fmap_42[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O3_N10_S1),.chainout(chainout_10_O3));
logic signed [63:0] chainout_12_O3; 
logic signed [63:0] O3_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O3(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_44[7:0]),.ay( 9'sd1),.bx(input_fmap_46[7:0]),.by( 9'sd4),.cx(input_fmap_50[7:0]),.cy( 9'sd1),.dx(input_fmap_51[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O3_N12_S1),.chainout(chainout_12_O3));
logic signed [63:0] chainout_14_O3; 
logic signed [63:0] O3_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O3(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_55[7:0]),.ay( 9'sd1),.bx(input_fmap_57[7:0]),.by( 9'sd1),.cx(input_fmap_59[7:0]),.cy( 9'sd1),.dx(input_fmap_60[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O3_N14_S1),.chainout(chainout_14_O3));
logic signed [63:0] chainout_16_O3; 
logic signed [63:0] O3_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O3(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_61[7:0]),.ay(-9'sd2),.bx(input_fmap_62[7:0]),.by(-9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O3_N16_S1),.chainout(chainout_16_O3));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O3_N0_S2;		always @(posedge clk) O3_N0_S2 <=     O3_N0_S1  +  O3_N2_S1 ;
 logic signed [21:0] O3_N2_S2;		always @(posedge clk) O3_N2_S2 <=     O3_N4_S1  +  O3_N6_S1 ;
 logic signed [21:0] O3_N4_S2;		always @(posedge clk) O3_N4_S2 <=     O3_N8_S1  +  O3_N10_S1 ;
 logic signed [21:0] O3_N6_S2;		always @(posedge clk) O3_N6_S2 <=     O3_N12_S1  +  O3_N14_S1 ;
 logic signed [21:0] O3_N8_S2;		always @(posedge clk) O3_N8_S2 <=     O3_N16_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O3_N0_S3;		always @(posedge clk) O3_N0_S3 <=     O3_N0_S2  +  O3_N2_S2 ;
 logic signed [22:0] O3_N2_S3;		always @(posedge clk) O3_N2_S3 <=     O3_N4_S2  +  O3_N6_S2 ;
 logic signed [22:0] O3_N4_S3;		always @(posedge clk) O3_N4_S3 <=     O3_N8_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O3_N0_S4;		always @(posedge clk) O3_N0_S4 <=     O3_N0_S3  +  O3_N2_S3 ;
 logic signed [23:0] O3_N2_S4;		always @(posedge clk) O3_N2_S4 <=     O3_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O3_N0_S5;		always @(posedge clk) O3_N0_S5 <=     O3_N0_S4  +  O3_N2_S4 ;
 assign conv_mac_3 = O3_N0_S5;

logic signed [31:0] conv_mac_4;
logic signed [63:0] chainout_0_O4; 
logic signed [63:0] O4_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O4(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay( 9'sd1),.bx(input_fmap_2[7:0]),.by( 9'sd1),.cx(input_fmap_3[7:0]),.cy( 9'sd1),.dx(input_fmap_4[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O4_N0_S1),.chainout(chainout_0_O4));
logic signed [63:0] chainout_2_O4; 
logic signed [63:0] O4_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O4(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_6[7:0]),.ay( 9'sd1),.bx(input_fmap_9[7:0]),.by( 9'sd1),.cx(input_fmap_10[7:0]),.cy(-9'sd1),.dx(input_fmap_11[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O4_N2_S1),.chainout(chainout_2_O4));
logic signed [63:0] chainout_4_O4; 
logic signed [63:0] O4_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O4(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_12[7:0]),.ay( 9'sd1),.bx(input_fmap_13[7:0]),.by( 9'sd1),.cx(input_fmap_14[7:0]),.cy( 9'sd1),.dx(input_fmap_16[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O4_N4_S1),.chainout(chainout_4_O4));
logic signed [63:0] chainout_6_O4; 
logic signed [63:0] O4_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O4(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_17[7:0]),.ay(-9'sd1),.bx(input_fmap_24[7:0]),.by( 9'sd1),.cx(input_fmap_25[7:0]),.cy( 9'sd1),.dx(input_fmap_29[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O4_N6_S1),.chainout(chainout_6_O4));
logic signed [63:0] chainout_8_O4; 
logic signed [63:0] O4_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O4(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_30[7:0]),.ay( 9'sd1),.bx(input_fmap_31[7:0]),.by( 9'sd2),.cx(input_fmap_32[7:0]),.cy(-9'sd1),.dx(input_fmap_33[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O4_N8_S1),.chainout(chainout_8_O4));
logic signed [63:0] chainout_10_O4; 
logic signed [63:0] O4_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O4(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_34[7:0]),.ay(-9'sd1),.bx(input_fmap_38[7:0]),.by( 9'sd1),.cx(input_fmap_40[7:0]),.cy( 9'sd1),.dx(input_fmap_41[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O4_N10_S1),.chainout(chainout_10_O4));
logic signed [63:0] chainout_12_O4; 
logic signed [63:0] O4_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O4(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_42[7:0]),.ay( 9'sd2),.bx(input_fmap_47[7:0]),.by( 9'sd1),.cx(input_fmap_49[7:0]),.cy(-9'sd1),.dx(input_fmap_54[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O4_N12_S1),.chainout(chainout_12_O4));
logic signed [63:0] chainout_14_O4; 
logic signed [63:0] O4_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O4(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_55[7:0]),.ay(-9'sd1),.bx(input_fmap_56[7:0]),.by(-9'sd1),.cx(input_fmap_57[7:0]),.cy(-9'sd1),.dx(input_fmap_60[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O4_N14_S1),.chainout(chainout_14_O4));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O4_N0_S2;		always @(posedge clk) O4_N0_S2 <=     O4_N0_S1  +  O4_N2_S1 ;
 logic signed [21:0] O4_N2_S2;		always @(posedge clk) O4_N2_S2 <=     O4_N4_S1  +  O4_N6_S1 ;
 logic signed [21:0] O4_N4_S2;		always @(posedge clk) O4_N4_S2 <=     O4_N8_S1  +  O4_N10_S1 ;
 logic signed [21:0] O4_N6_S2;		always @(posedge clk) O4_N6_S2 <=     O4_N12_S1  +  O4_N14_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O4_N0_S3;		always @(posedge clk) O4_N0_S3 <=     O4_N0_S2  +  O4_N2_S2 ;
 logic signed [22:0] O4_N2_S3;		always @(posedge clk) O4_N2_S3 <=     O4_N4_S2  +  O4_N6_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O4_N0_S4;		always @(posedge clk) O4_N0_S4 <=     O4_N0_S3  +  O4_N2_S3 ;
 assign conv_mac_4 = O4_N0_S4;

logic signed [31:0] conv_mac_5;
logic signed [63:0] chainout_0_O5; 
logic signed [63:0] O5_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O5(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd1),.bx(input_fmap_2[7:0]),.by(-9'sd1),.cx(input_fmap_4[7:0]),.cy( 9'sd1),.dx(input_fmap_6[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O5_N0_S1),.chainout(chainout_0_O5));
logic signed [63:0] chainout_2_O5; 
logic signed [63:0] O5_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O5(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_11[7:0]),.ay( 9'sd1),.bx(input_fmap_13[7:0]),.by(-9'sd1),.cx(input_fmap_14[7:0]),.cy(-9'sd1),.dx(input_fmap_16[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O5_N2_S1),.chainout(chainout_2_O5));
logic signed [63:0] chainout_4_O5; 
logic signed [63:0] O5_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O5(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_17[7:0]),.ay( 9'sd1),.bx(input_fmap_18[7:0]),.by( 9'sd1),.cx(input_fmap_25[7:0]),.cy(-9'sd1),.dx(input_fmap_26[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O5_N4_S1),.chainout(chainout_4_O5));
logic signed [63:0] chainout_6_O5; 
logic signed [63:0] O5_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O5(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_29[7:0]),.ay(-9'sd2),.bx(input_fmap_32[7:0]),.by( 9'sd1),.cx(input_fmap_33[7:0]),.cy(-9'sd1),.dx(input_fmap_39[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O5_N6_S1),.chainout(chainout_6_O5));
logic signed [63:0] chainout_8_O5; 
logic signed [63:0] O5_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O5(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_41[7:0]),.ay(-9'sd1),.bx(input_fmap_42[7:0]),.by( 9'sd2),.cx(input_fmap_46[7:0]),.cy(-9'sd1),.dx(input_fmap_47[7:0]),.dy( 9'sd3),.chainin(63'd0),.result(O5_N8_S1),.chainout(chainout_8_O5));
logic signed [63:0] chainout_10_O5; 
logic signed [63:0] O5_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O5(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_50[7:0]),.ay(-9'sd1),.bx(input_fmap_54[7:0]),.by(-9'sd1),.cx(input_fmap_55[7:0]),.cy(-9'sd1),.dx(input_fmap_56[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O5_N10_S1),.chainout(chainout_10_O5));
logic signed [63:0] chainout_12_O5; 
logic signed [63:0] O5_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O5(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_60[7:0]),.ay(-9'sd1),.bx(input_fmap_63[7:0]),.by( 9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O5_N12_S1),.chainout(chainout_12_O5));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O5_N0_S2;		always @(posedge clk) O5_N0_S2 <=     O5_N0_S1  +  O5_N2_S1 ;
 logic signed [21:0] O5_N2_S2;		always @(posedge clk) O5_N2_S2 <=     O5_N4_S1  +  O5_N6_S1 ;
 logic signed [21:0] O5_N4_S2;		always @(posedge clk) O5_N4_S2 <=     O5_N8_S1  +  O5_N10_S1 ;
 logic signed [21:0] O5_N6_S2;		always @(posedge clk) O5_N6_S2 <=     O5_N12_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O5_N0_S3;		always @(posedge clk) O5_N0_S3 <=     O5_N0_S2  +  O5_N2_S2 ;
 logic signed [22:0] O5_N2_S3;		always @(posedge clk) O5_N2_S3 <=     O5_N4_S2  +  O5_N6_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O5_N0_S4;		always @(posedge clk) O5_N0_S4 <=     O5_N0_S3  +  O5_N2_S3 ;
 assign conv_mac_5 = O5_N0_S4;

logic signed [31:0] conv_mac_6;
logic signed [63:0] chainout_0_O6; 
logic signed [63:0] O6_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O6(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay( 9'sd1),.bx(input_fmap_2[7:0]),.by( 9'sd3),.cx(input_fmap_3[7:0]),.cy(-9'sd2),.dx(input_fmap_4[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O6_N0_S1),.chainout(chainout_0_O6));
logic signed [63:0] chainout_2_O6; 
logic signed [63:0] O6_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O6(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_6[7:0]),.ay( 9'sd2),.bx(input_fmap_7[7:0]),.by( 9'sd1),.cx(input_fmap_10[7:0]),.cy( 9'sd1),.dx(input_fmap_11[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O6_N2_S1),.chainout(chainout_2_O6));
logic signed [63:0] chainout_4_O6; 
logic signed [63:0] O6_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O6(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_12[7:0]),.ay(-9'sd1),.bx(input_fmap_13[7:0]),.by(-9'sd1),.cx(input_fmap_14[7:0]),.cy( 9'sd2),.dx(input_fmap_15[7:0]),.dy(-9'sd3),.chainin(63'd0),.result(O6_N4_S1),.chainout(chainout_4_O6));
logic signed [63:0] chainout_6_O6; 
logic signed [63:0] O6_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O6(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_17[7:0]),.ay( 9'sd2),.bx(input_fmap_18[7:0]),.by(-9'sd3),.cx(input_fmap_19[7:0]),.cy(-9'sd1),.dx(input_fmap_20[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O6_N6_S1),.chainout(chainout_6_O6));
logic signed [63:0] chainout_8_O6; 
logic signed [63:0] O6_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O6(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_22[7:0]),.ay( 9'sd2),.bx(input_fmap_23[7:0]),.by(-9'sd1),.cx(input_fmap_25[7:0]),.cy( 9'sd1),.dx(input_fmap_26[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O6_N8_S1),.chainout(chainout_8_O6));
logic signed [63:0] chainout_10_O6; 
logic signed [63:0] O6_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O6(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_27[7:0]),.ay( 9'sd1),.bx(input_fmap_28[7:0]),.by( 9'sd1),.cx(input_fmap_30[7:0]),.cy( 9'sd1),.dx(input_fmap_31[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O6_N10_S1),.chainout(chainout_10_O6));
logic signed [63:0] chainout_12_O6; 
logic signed [63:0] O6_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O6(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_33[7:0]),.ay(-9'sd2),.bx(input_fmap_34[7:0]),.by(-9'sd1),.cx(input_fmap_35[7:0]),.cy(-9'sd2),.dx(input_fmap_36[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O6_N12_S1),.chainout(chainout_12_O6));
logic signed [63:0] chainout_14_O6; 
logic signed [63:0] O6_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O6(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_37[7:0]),.ay(-9'sd2),.bx(input_fmap_38[7:0]),.by(-9'sd1),.cx(input_fmap_40[7:0]),.cy( 9'sd1),.dx(input_fmap_42[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O6_N14_S1),.chainout(chainout_14_O6));
logic signed [63:0] chainout_16_O6; 
logic signed [63:0] O6_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O6(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_43[7:0]),.ay(-9'sd2),.bx(input_fmap_45[7:0]),.by( 9'sd2),.cx(input_fmap_46[7:0]),.cy( 9'sd1),.dx(input_fmap_47[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O6_N16_S1),.chainout(chainout_16_O6));
logic signed [63:0] chainout_18_O6; 
logic signed [63:0] O6_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O6(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_48[7:0]),.ay( 9'sd2),.bx(input_fmap_50[7:0]),.by( 9'sd1),.cx(input_fmap_52[7:0]),.cy(-9'sd1),.dx(input_fmap_53[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O6_N18_S1),.chainout(chainout_18_O6));
logic signed [63:0] chainout_20_O6; 
logic signed [63:0] O6_N20_S1; 
 int_sop_4_wrapper int_sop_4_inst_20_O6(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_55[7:0]),.ay(-9'sd2),.bx(input_fmap_57[7:0]),.by( 9'sd1),.cx(input_fmap_59[7:0]),.cy( 9'sd4),.dx(input_fmap_60[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O6_N20_S1),.chainout(chainout_20_O6));
logic signed [63:0] chainout_22_O6; 
logic signed [63:0] O6_N22_S1; 
 int_sop_4_wrapper int_sop_4_inst_22_O6(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_61[7:0]),.ay(-9'sd1),.bx(input_fmap_62[7:0]),.by(-9'sd1),.cx(input_fmap_63[7:0]),.cy(-9'sd1),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O6_N22_S1),.chainout(chainout_22_O6));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O6_N0_S2;		always @(posedge clk) O6_N0_S2 <=     O6_N0_S1  +  O6_N2_S1 ;
 logic signed [21:0] O6_N2_S2;		always @(posedge clk) O6_N2_S2 <=     O6_N4_S1  +  O6_N6_S1 ;
 logic signed [21:0] O6_N4_S2;		always @(posedge clk) O6_N4_S2 <=     O6_N8_S1  +  O6_N10_S1 ;
 logic signed [21:0] O6_N6_S2;		always @(posedge clk) O6_N6_S2 <=     O6_N12_S1  +  O6_N14_S1 ;
 logic signed [21:0] O6_N8_S2;		always @(posedge clk) O6_N8_S2 <=     O6_N16_S1  +  O6_N18_S1 ;
 logic signed [21:0] O6_N10_S2;		always @(posedge clk) O6_N10_S2 <=     O6_N20_S1  +  O6_N22_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O6_N0_S3;		always @(posedge clk) O6_N0_S3 <=     O6_N0_S2  +  O6_N2_S2 ;
 logic signed [22:0] O6_N2_S3;		always @(posedge clk) O6_N2_S3 <=     O6_N4_S2  +  O6_N6_S2 ;
 logic signed [22:0] O6_N4_S3;		always @(posedge clk) O6_N4_S3 <=     O6_N8_S2  +  O6_N10_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O6_N0_S4;		always @(posedge clk) O6_N0_S4 <=     O6_N0_S3  +  O6_N2_S3 ;
 logic signed [23:0] O6_N2_S4;		always @(posedge clk) O6_N2_S4 <=     O6_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O6_N0_S5;		always @(posedge clk) O6_N0_S5 <=     O6_N0_S4  +  O6_N2_S4 ;
 assign conv_mac_6 = O6_N0_S5;

logic signed [31:0] conv_mac_7;
logic signed [63:0] chainout_0_O7; 
logic signed [63:0] O7_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O7(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay( 9'sd1),.bx(input_fmap_5[7:0]),.by(-9'sd1),.cx(input_fmap_10[7:0]),.cy(-9'sd2),.dx(input_fmap_11[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O7_N0_S1),.chainout(chainout_0_O7));
logic signed [63:0] chainout_2_O7; 
logic signed [63:0] O7_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O7(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_16[7:0]),.ay(-9'sd1),.bx(input_fmap_17[7:0]),.by(-9'sd3),.cx(input_fmap_19[7:0]),.cy(-9'sd1),.dx(input_fmap_25[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O7_N2_S1),.chainout(chainout_2_O7));
logic signed [63:0] chainout_4_O7; 
logic signed [63:0] O7_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O7(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_26[7:0]),.ay(-9'sd1),.bx(input_fmap_27[7:0]),.by(-9'sd2),.cx(input_fmap_28[7:0]),.cy(-9'sd1),.dx(input_fmap_30[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O7_N4_S1),.chainout(chainout_4_O7));
logic signed [63:0] chainout_6_O7; 
logic signed [63:0] O7_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O7(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_31[7:0]),.ay(-9'sd1),.bx(input_fmap_33[7:0]),.by(-9'sd1),.cx(input_fmap_38[7:0]),.cy(-9'sd1),.dx(input_fmap_40[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O7_N6_S1),.chainout(chainout_6_O7));
logic signed [63:0] chainout_8_O7; 
logic signed [63:0] O7_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O7(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_45[7:0]),.ay(-9'sd1),.bx(input_fmap_46[7:0]),.by(-9'sd1),.cx(input_fmap_47[7:0]),.cy( 9'sd1),.dx(input_fmap_48[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O7_N8_S1),.chainout(chainout_8_O7));
logic signed [63:0] chainout_10_O7; 
logic signed [63:0] O7_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O7(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_50[7:0]),.ay(-9'sd1),.bx(input_fmap_52[7:0]),.by(-9'sd1),.cx(input_fmap_53[7:0]),.cy( 9'sd1),.dx(input_fmap_58[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O7_N10_S1),.chainout(chainout_10_O7));
logic signed [63:0] chainout_12_O7; 
logic signed [63:0] O7_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O7(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_60[7:0]),.ay(-9'sd1),.bx(input_fmap_62[7:0]),.by( 9'sd2),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O7_N12_S1),.chainout(chainout_12_O7));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O7_N0_S2;		always @(posedge clk) O7_N0_S2 <=     O7_N0_S1  +  O7_N2_S1 ;
 logic signed [21:0] O7_N2_S2;		always @(posedge clk) O7_N2_S2 <=     O7_N4_S1  +  O7_N6_S1 ;
 logic signed [21:0] O7_N4_S2;		always @(posedge clk) O7_N4_S2 <=     O7_N8_S1  +  O7_N10_S1 ;
 logic signed [21:0] O7_N6_S2;		always @(posedge clk) O7_N6_S2 <=     O7_N12_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O7_N0_S3;		always @(posedge clk) O7_N0_S3 <=     O7_N0_S2  +  O7_N2_S2 ;
 logic signed [22:0] O7_N2_S3;		always @(posedge clk) O7_N2_S3 <=     O7_N4_S2  +  O7_N6_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O7_N0_S4;		always @(posedge clk) O7_N0_S4 <=     O7_N0_S3  +  O7_N2_S3 ;
 assign conv_mac_7 = O7_N0_S4;

logic signed [31:0] conv_mac_8;
logic signed [63:0] chainout_0_O8; 
logic signed [63:0] O8_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O8(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_11[7:0]),.ay( 9'sd1),.bx(input_fmap_12[7:0]),.by( 9'sd1),.cx(input_fmap_16[7:0]),.cy( 9'sd1),.dx(input_fmap_25[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O8_N0_S1),.chainout(chainout_0_O8));
logic signed [63:0] chainout_2_O8; 
logic signed [63:0] O8_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O8(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_26[7:0]),.ay( 9'sd2),.bx(input_fmap_31[7:0]),.by( 9'sd1),.cx(input_fmap_33[7:0]),.cy( 9'sd1),.dx(input_fmap_35[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O8_N2_S1),.chainout(chainout_2_O8));
logic signed [63:0] chainout_4_O8; 
logic signed [63:0] O8_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O8(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_39[7:0]),.ay( 9'sd1),.bx(input_fmap_40[7:0]),.by( 9'sd2),.cx(input_fmap_42[7:0]),.cy(-9'sd1),.dx(input_fmap_60[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O8_N4_S1),.chainout(chainout_4_O8));
logic signed [63:0] chainout_6_O8; 
logic signed [63:0] O8_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O8(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_62[7:0]),.ay( 9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O8_N6_S1),.chainout(chainout_6_O8));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O8_N0_S2;		always @(posedge clk) O8_N0_S2 <=     O8_N0_S1  +  O8_N2_S1 ;
 logic signed [21:0] O8_N2_S2;		always @(posedge clk) O8_N2_S2 <=     O8_N4_S1  +  O8_N6_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O8_N0_S3;		always @(posedge clk) O8_N0_S3 <=     O8_N0_S2  +  O8_N2_S2 ;
 assign conv_mac_8 = O8_N0_S3;

logic signed [31:0] conv_mac_9;
logic signed [63:0] chainout_0_O9; 
logic signed [63:0] O9_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O9(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay( 9'sd4),.bx(input_fmap_5[7:0]),.by(-9'sd1),.cx(input_fmap_6[7:0]),.cy(-9'sd1),.dx(input_fmap_8[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O9_N0_S1),.chainout(chainout_0_O9));
logic signed [63:0] chainout_2_O9; 
logic signed [63:0] O9_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O9(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_10[7:0]),.ay( 9'sd1),.bx(input_fmap_11[7:0]),.by(-9'sd1),.cx(input_fmap_15[7:0]),.cy(-9'sd1),.dx(input_fmap_16[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O9_N2_S1),.chainout(chainout_2_O9));
logic signed [63:0] chainout_4_O9; 
logic signed [63:0] O9_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O9(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_19[7:0]),.ay( 9'sd1),.bx(input_fmap_20[7:0]),.by(-9'sd1),.cx(input_fmap_29[7:0]),.cy( 9'sd1),.dx(input_fmap_32[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O9_N4_S1),.chainout(chainout_4_O9));
logic signed [63:0] chainout_6_O9; 
logic signed [63:0] O9_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O9(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_41[7:0]),.ay( 9'sd1),.bx(input_fmap_42[7:0]),.by( 9'sd1),.cx(input_fmap_45[7:0]),.cy(-9'sd2),.dx(input_fmap_46[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O9_N6_S1),.chainout(chainout_6_O9));
logic signed [63:0] chainout_8_O9; 
logic signed [63:0] O9_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O9(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_47[7:0]),.ay( 9'sd1),.bx(input_fmap_52[7:0]),.by( 9'sd1),.cx(input_fmap_55[7:0]),.cy(-9'sd1),.dx(input_fmap_56[7:0]),.dy(-9'sd4),.chainin(63'd0),.result(O9_N8_S1),.chainout(chainout_8_O9));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O9_N0_S2;		always @(posedge clk) O9_N0_S2 <=     O9_N0_S1  +  O9_N2_S1 ;
 logic signed [21:0] O9_N2_S2;		always @(posedge clk) O9_N2_S2 <=     O9_N4_S1  +  O9_N6_S1 ;
 logic signed [21:0] O9_N4_S2;		always @(posedge clk) O9_N4_S2 <=     O9_N8_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O9_N0_S3;		always @(posedge clk) O9_N0_S3 <=     O9_N0_S2  +  O9_N2_S2 ;
 logic signed [22:0] O9_N2_S3;		always @(posedge clk) O9_N2_S3 <=     O9_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O9_N0_S4;		always @(posedge clk) O9_N0_S4 <=     O9_N0_S3  +  O9_N2_S3 ;
 assign conv_mac_9 = O9_N0_S4;

logic signed [31:0] conv_mac_10;
logic signed [63:0] chainout_0_O10; 
logic signed [63:0] O10_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O10(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_4[7:0]),.ay( 9'sd1),.bx(input_fmap_5[7:0]),.by( 9'sd4),.cx(input_fmap_6[7:0]),.cy( 9'sd1),.dx(input_fmap_7[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O10_N0_S1),.chainout(chainout_0_O10));
logic signed [63:0] chainout_2_O10; 
logic signed [63:0] O10_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O10(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_8[7:0]),.ay(-9'sd1),.bx(input_fmap_13[7:0]),.by( 9'sd1),.cx(input_fmap_17[7:0]),.cy(-9'sd1),.dx(input_fmap_18[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O10_N2_S1),.chainout(chainout_2_O10));
logic signed [63:0] chainout_4_O10; 
logic signed [63:0] O10_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O10(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_19[7:0]),.ay( 9'sd1),.bx(input_fmap_22[7:0]),.by(-9'sd1),.cx(input_fmap_23[7:0]),.cy( 9'sd2),.dx(input_fmap_24[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O10_N4_S1),.chainout(chainout_4_O10));
logic signed [63:0] chainout_6_O10; 
logic signed [63:0] O10_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O10(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_25[7:0]),.ay( 9'sd1),.bx(input_fmap_27[7:0]),.by( 9'sd2),.cx(input_fmap_28[7:0]),.cy( 9'sd1),.dx(input_fmap_29[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O10_N6_S1),.chainout(chainout_6_O10));
logic signed [63:0] chainout_8_O10; 
logic signed [63:0] O10_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O10(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_30[7:0]),.ay(-9'sd1),.bx(input_fmap_31[7:0]),.by(-9'sd1),.cx(input_fmap_32[7:0]),.cy(-9'sd1),.dx(input_fmap_33[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O10_N8_S1),.chainout(chainout_8_O10));
logic signed [63:0] chainout_10_O10; 
logic signed [63:0] O10_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O10(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_35[7:0]),.ay( 9'sd1),.bx(input_fmap_36[7:0]),.by( 9'sd1),.cx(input_fmap_37[7:0]),.cy( 9'sd1),.dx(input_fmap_39[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O10_N10_S1),.chainout(chainout_10_O10));
logic signed [63:0] chainout_12_O10; 
logic signed [63:0] O10_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O10(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_40[7:0]),.ay( 9'sd1),.bx(input_fmap_41[7:0]),.by(-9'sd1),.cx(input_fmap_42[7:0]),.cy( 9'sd1),.dx(input_fmap_43[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O10_N12_S1),.chainout(chainout_12_O10));
logic signed [63:0] chainout_14_O10; 
logic signed [63:0] O10_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O10(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_44[7:0]),.ay(-9'sd2),.bx(input_fmap_45[7:0]),.by( 9'sd1),.cx(input_fmap_46[7:0]),.cy(-9'sd2),.dx(input_fmap_51[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O10_N14_S1),.chainout(chainout_14_O10));
logic signed [63:0] chainout_16_O10; 
logic signed [63:0] O10_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O10(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_52[7:0]),.ay(-9'sd1),.bx(input_fmap_62[7:0]),.by(-9'sd1),.cx(input_fmap_63[7:0]),.cy( 9'sd1),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O10_N16_S1),.chainout(chainout_16_O10));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O10_N0_S2;		always @(posedge clk) O10_N0_S2 <=     O10_N0_S1  +  O10_N2_S1 ;
 logic signed [21:0] O10_N2_S2;		always @(posedge clk) O10_N2_S2 <=     O10_N4_S1  +  O10_N6_S1 ;
 logic signed [21:0] O10_N4_S2;		always @(posedge clk) O10_N4_S2 <=     O10_N8_S1  +  O10_N10_S1 ;
 logic signed [21:0] O10_N6_S2;		always @(posedge clk) O10_N6_S2 <=     O10_N12_S1  +  O10_N14_S1 ;
 logic signed [21:0] O10_N8_S2;		always @(posedge clk) O10_N8_S2 <=     O10_N16_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O10_N0_S3;		always @(posedge clk) O10_N0_S3 <=     O10_N0_S2  +  O10_N2_S2 ;
 logic signed [22:0] O10_N2_S3;		always @(posedge clk) O10_N2_S3 <=     O10_N4_S2  +  O10_N6_S2 ;
 logic signed [22:0] O10_N4_S3;		always @(posedge clk) O10_N4_S3 <=     O10_N8_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O10_N0_S4;		always @(posedge clk) O10_N0_S4 <=     O10_N0_S3  +  O10_N2_S3 ;
 logic signed [23:0] O10_N2_S4;		always @(posedge clk) O10_N2_S4 <=     O10_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O10_N0_S5;		always @(posedge clk) O10_N0_S5 <=     O10_N0_S4  +  O10_N2_S4 ;
 assign conv_mac_10 = O10_N0_S5;

logic signed [31:0] conv_mac_11;
logic signed [63:0] chainout_0_O11; 
logic signed [63:0] O11_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O11(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd2),.bx(input_fmap_4[7:0]),.by(-9'sd1),.cx(input_fmap_9[7:0]),.cy( 9'sd1),.dx(input_fmap_10[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O11_N0_S1),.chainout(chainout_0_O11));
logic signed [63:0] chainout_2_O11; 
logic signed [63:0] O11_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O11(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_11[7:0]),.ay(-9'sd1),.bx(input_fmap_14[7:0]),.by(-9'sd2),.cx(input_fmap_16[7:0]),.cy( 9'sd1),.dx(input_fmap_18[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O11_N2_S1),.chainout(chainout_2_O11));
logic signed [63:0] chainout_4_O11; 
logic signed [63:0] O11_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O11(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_19[7:0]),.ay(-9'sd1),.bx(input_fmap_20[7:0]),.by( 9'sd1),.cx(input_fmap_21[7:0]),.cy( 9'sd2),.dx(input_fmap_22[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O11_N4_S1),.chainout(chainout_4_O11));
logic signed [63:0] chainout_6_O11; 
logic signed [63:0] O11_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O11(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_23[7:0]),.ay( 9'sd1),.bx(input_fmap_25[7:0]),.by( 9'sd1),.cx(input_fmap_30[7:0]),.cy( 9'sd1),.dx(input_fmap_31[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O11_N6_S1),.chainout(chainout_6_O11));
logic signed [63:0] chainout_8_O11; 
logic signed [63:0] O11_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O11(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_32[7:0]),.ay( 9'sd1),.bx(input_fmap_33[7:0]),.by( 9'sd1),.cx(input_fmap_37[7:0]),.cy( 9'sd1),.dx(input_fmap_40[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O11_N8_S1),.chainout(chainout_8_O11));
logic signed [63:0] chainout_10_O11; 
logic signed [63:0] O11_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O11(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_42[7:0]),.ay( 9'sd1),.bx(input_fmap_43[7:0]),.by( 9'sd1),.cx(input_fmap_46[7:0]),.cy( 9'sd1),.dx(input_fmap_47[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O11_N10_S1),.chainout(chainout_10_O11));
logic signed [63:0] chainout_12_O11; 
logic signed [63:0] O11_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O11(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_50[7:0]),.ay( 9'sd1),.bx(input_fmap_51[7:0]),.by(-9'sd2),.cx(input_fmap_52[7:0]),.cy(-9'sd1),.dx(input_fmap_54[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O11_N12_S1),.chainout(chainout_12_O11));
logic signed [63:0] chainout_14_O11; 
logic signed [63:0] O11_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O11(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_56[7:0]),.ay( 9'sd1),.bx(input_fmap_58[7:0]),.by( 9'sd1),.cx(input_fmap_59[7:0]),.cy( 9'sd1),.dx(input_fmap_60[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O11_N14_S1),.chainout(chainout_14_O11));
logic signed [63:0] chainout_16_O11; 
logic signed [63:0] O11_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O11(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_63[7:0]),.ay( 9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O11_N16_S1),.chainout(chainout_16_O11));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O11_N0_S2;		always @(posedge clk) O11_N0_S2 <=     O11_N0_S1  +  O11_N2_S1 ;
 logic signed [21:0] O11_N2_S2;		always @(posedge clk) O11_N2_S2 <=     O11_N4_S1  +  O11_N6_S1 ;
 logic signed [21:0] O11_N4_S2;		always @(posedge clk) O11_N4_S2 <=     O11_N8_S1  +  O11_N10_S1 ;
 logic signed [21:0] O11_N6_S2;		always @(posedge clk) O11_N6_S2 <=     O11_N12_S1  +  O11_N14_S1 ;
 logic signed [21:0] O11_N8_S2;		always @(posedge clk) O11_N8_S2 <=     O11_N16_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O11_N0_S3;		always @(posedge clk) O11_N0_S3 <=     O11_N0_S2  +  O11_N2_S2 ;
 logic signed [22:0] O11_N2_S3;		always @(posedge clk) O11_N2_S3 <=     O11_N4_S2  +  O11_N6_S2 ;
 logic signed [22:0] O11_N4_S3;		always @(posedge clk) O11_N4_S3 <=     O11_N8_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O11_N0_S4;		always @(posedge clk) O11_N0_S4 <=     O11_N0_S3  +  O11_N2_S3 ;
 logic signed [23:0] O11_N2_S4;		always @(posedge clk) O11_N2_S4 <=     O11_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O11_N0_S5;		always @(posedge clk) O11_N0_S5 <=     O11_N0_S4  +  O11_N2_S4 ;
 assign conv_mac_11 = O11_N0_S5;

logic signed [31:0] conv_mac_12;
logic signed [63:0] chainout_0_O12; 
logic signed [63:0] O12_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O12(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_4[7:0]),.ay( 9'sd1),.bx(input_fmap_5[7:0]),.by(-9'sd1),.cx(input_fmap_7[7:0]),.cy( 9'sd1),.dx(input_fmap_11[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O12_N0_S1),.chainout(chainout_0_O12));
logic signed [63:0] chainout_2_O12; 
logic signed [63:0] O12_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O12(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_17[7:0]),.ay( 9'sd1),.bx(input_fmap_18[7:0]),.by( 9'sd1),.cx(input_fmap_19[7:0]),.cy( 9'sd1),.dx(input_fmap_23[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O12_N2_S1),.chainout(chainout_2_O12));
logic signed [63:0] chainout_4_O12; 
logic signed [63:0] O12_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O12(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_28[7:0]),.ay( 9'sd1),.bx(input_fmap_30[7:0]),.by(-9'sd1),.cx(input_fmap_31[7:0]),.cy( 9'sd2),.dx(input_fmap_35[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O12_N4_S1),.chainout(chainout_4_O12));
logic signed [63:0] chainout_6_O12; 
logic signed [63:0] O12_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O12(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_43[7:0]),.ay( 9'sd2),.bx(input_fmap_46[7:0]),.by( 9'sd1),.cx(input_fmap_52[7:0]),.cy( 9'sd1),.dx(input_fmap_53[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O12_N6_S1),.chainout(chainout_6_O12));
logic signed [63:0] chainout_8_O12; 
logic signed [63:0] O12_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O12(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_54[7:0]),.ay( 9'sd1),.bx(input_fmap_58[7:0]),.by( 9'sd1),.cx(input_fmap_59[7:0]),.cy( 9'sd1),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O12_N8_S1),.chainout(chainout_8_O12));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O12_N0_S2;		always @(posedge clk) O12_N0_S2 <=     O12_N0_S1  +  O12_N2_S1 ;
 logic signed [21:0] O12_N2_S2;		always @(posedge clk) O12_N2_S2 <=     O12_N4_S1  +  O12_N6_S1 ;
 logic signed [21:0] O12_N4_S2;		always @(posedge clk) O12_N4_S2 <=     O12_N8_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O12_N0_S3;		always @(posedge clk) O12_N0_S3 <=     O12_N0_S2  +  O12_N2_S2 ;
 logic signed [22:0] O12_N2_S3;		always @(posedge clk) O12_N2_S3 <=     O12_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O12_N0_S4;		always @(posedge clk) O12_N0_S4 <=     O12_N0_S3  +  O12_N2_S3 ;
 assign conv_mac_12 = O12_N0_S4;

logic signed [31:0] conv_mac_13;
logic signed [63:0] chainout_0_O13; 
logic signed [63:0] O13_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O13(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_3[7:0]),.ay(-9'sd4),.bx(input_fmap_5[7:0]),.by(-9'sd3),.cx(input_fmap_6[7:0]),.cy( 9'sd1),.dx(input_fmap_7[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O13_N0_S1),.chainout(chainout_0_O13));
logic signed [63:0] chainout_2_O13; 
logic signed [63:0] O13_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O13(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_9[7:0]),.ay(-9'sd1),.bx(input_fmap_10[7:0]),.by(-9'sd2),.cx(input_fmap_12[7:0]),.cy(-9'sd3),.dx(input_fmap_13[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O13_N2_S1),.chainout(chainout_2_O13));
logic signed [63:0] chainout_4_O13; 
logic signed [63:0] O13_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O13(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_14[7:0]),.ay(-9'sd1),.bx(input_fmap_17[7:0]),.by(-9'sd1),.cx(input_fmap_19[7:0]),.cy(-9'sd4),.dx(input_fmap_20[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O13_N4_S1),.chainout(chainout_4_O13));
logic signed [63:0] chainout_6_O13; 
logic signed [63:0] O13_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O13(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_21[7:0]),.ay( 9'sd2),.bx(input_fmap_22[7:0]),.by( 9'sd1),.cx(input_fmap_23[7:0]),.cy( 9'sd2),.dx(input_fmap_24[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O13_N6_S1),.chainout(chainout_6_O13));
logic signed [63:0] chainout_8_O13; 
logic signed [63:0] O13_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O13(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_25[7:0]),.ay(-9'sd1),.bx(input_fmap_26[7:0]),.by(-9'sd2),.cx(input_fmap_27[7:0]),.cy( 9'sd1),.dx(input_fmap_28[7:0]),.dy(-9'sd3),.chainin(63'd0),.result(O13_N8_S1),.chainout(chainout_8_O13));
logic signed [63:0] chainout_10_O13; 
logic signed [63:0] O13_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O13(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_29[7:0]),.ay( 9'sd3),.bx(input_fmap_31[7:0]),.by( 9'sd1),.cx(input_fmap_32[7:0]),.cy( 9'sd2),.dx(input_fmap_33[7:0]),.dy( 9'sd3),.chainin(63'd0),.result(O13_N10_S1),.chainout(chainout_10_O13));
logic signed [63:0] chainout_12_O13; 
logic signed [63:0] O13_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O13(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_34[7:0]),.ay(-9'sd2),.bx(input_fmap_35[7:0]),.by( 9'sd2),.cx(input_fmap_36[7:0]),.cy(-9'sd1),.dx(input_fmap_37[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O13_N12_S1),.chainout(chainout_12_O13));
logic signed [63:0] chainout_14_O13; 
logic signed [63:0] O13_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O13(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_38[7:0]),.ay( 9'sd4),.bx(input_fmap_39[7:0]),.by(-9'sd2),.cx(input_fmap_41[7:0]),.cy(-9'sd1),.dx(input_fmap_43[7:0]),.dy( 9'sd3),.chainin(63'd0),.result(O13_N14_S1),.chainout(chainout_14_O13));
logic signed [63:0] chainout_16_O13; 
logic signed [63:0] O13_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O13(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_45[7:0]),.ay(-9'sd1),.bx(input_fmap_46[7:0]),.by(-9'sd3),.cx(input_fmap_47[7:0]),.cy(-9'sd3),.dx(input_fmap_48[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O13_N16_S1),.chainout(chainout_16_O13));
logic signed [63:0] chainout_18_O13; 
logic signed [63:0] O13_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O13(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_49[7:0]),.ay(-9'sd2),.bx(input_fmap_50[7:0]),.by( 9'sd1),.cx(input_fmap_51[7:0]),.cy(-9'sd3),.dx(input_fmap_52[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O13_N18_S1),.chainout(chainout_18_O13));
logic signed [63:0] chainout_20_O13; 
logic signed [63:0] O13_N20_S1; 
 int_sop_4_wrapper int_sop_4_inst_20_O13(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_53[7:0]),.ay( 9'sd1),.bx(input_fmap_55[7:0]),.by(-9'sd2),.cx(input_fmap_56[7:0]),.cy( 9'sd2),.dx(input_fmap_58[7:0]),.dy( 9'sd5),.chainin(63'd0),.result(O13_N20_S1),.chainout(chainout_20_O13));
logic signed [63:0] chainout_22_O13; 
logic signed [63:0] O13_N22_S1; 
 int_sop_4_wrapper int_sop_4_inst_22_O13(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_59[7:0]),.ay(-9'sd1),.bx(input_fmap_60[7:0]),.by(-9'sd1),.cx(input_fmap_61[7:0]),.cy(-9'sd1),.dx(input_fmap_62[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O13_N22_S1),.chainout(chainout_22_O13));
logic signed [63:0] chainout_24_O13; 
logic signed [63:0] O13_N24_S1; 
 int_sop_4_wrapper int_sop_4_inst_24_O13(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_63[7:0]),.ay( 9'sd3),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O13_N24_S1),.chainout(chainout_24_O13));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O13_N0_S2;		always @(posedge clk) O13_N0_S2 <=     O13_N0_S1  +  O13_N2_S1 ;
 logic signed [21:0] O13_N2_S2;		always @(posedge clk) O13_N2_S2 <=     O13_N4_S1  +  O13_N6_S1 ;
 logic signed [21:0] O13_N4_S2;		always @(posedge clk) O13_N4_S2 <=     O13_N8_S1  +  O13_N10_S1 ;
 logic signed [21:0] O13_N6_S2;		always @(posedge clk) O13_N6_S2 <=     O13_N12_S1  +  O13_N14_S1 ;
 logic signed [21:0] O13_N8_S2;		always @(posedge clk) O13_N8_S2 <=     O13_N16_S1  +  O13_N18_S1 ;
 logic signed [21:0] O13_N10_S2;		always @(posedge clk) O13_N10_S2 <=     O13_N20_S1  +  O13_N22_S1 ;
 logic signed [21:0] O13_N12_S2;		always @(posedge clk) O13_N12_S2 <=     O13_N24_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O13_N0_S3;		always @(posedge clk) O13_N0_S3 <=     O13_N0_S2  +  O13_N2_S2 ;
 logic signed [22:0] O13_N2_S3;		always @(posedge clk) O13_N2_S3 <=     O13_N4_S2  +  O13_N6_S2 ;
 logic signed [22:0] O13_N4_S3;		always @(posedge clk) O13_N4_S3 <=     O13_N8_S2  +  O13_N10_S2 ;
 logic signed [22:0] O13_N6_S3;		always @(posedge clk) O13_N6_S3 <=     O13_N12_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O13_N0_S4;		always @(posedge clk) O13_N0_S4 <=     O13_N0_S3  +  O13_N2_S3 ;
 logic signed [23:0] O13_N2_S4;		always @(posedge clk) O13_N2_S4 <=     O13_N4_S3  +  O13_N6_S3 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O13_N0_S5;		always @(posedge clk) O13_N0_S5 <=     O13_N0_S4  +  O13_N2_S4 ;
 assign conv_mac_13 = O13_N0_S5;

logic signed [31:0] conv_mac_14;
logic signed [63:0] chainout_0_O14; 
logic signed [63:0] O14_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O14(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd1),.bx(input_fmap_1[7:0]),.by(-9'sd1),.cx(input_fmap_3[7:0]),.cy( 9'sd1),.dx(input_fmap_4[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O14_N0_S1),.chainout(chainout_0_O14));
logic signed [63:0] chainout_2_O14; 
logic signed [63:0] O14_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O14(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_5[7:0]),.ay(-9'sd3),.bx(input_fmap_6[7:0]),.by(-9'sd1),.cx(input_fmap_7[7:0]),.cy(-9'sd1),.dx(input_fmap_9[7:0]),.dy( 9'sd4),.chainin(63'd0),.result(O14_N2_S1),.chainout(chainout_2_O14));
logic signed [63:0] chainout_4_O14; 
logic signed [63:0] O14_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O14(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_10[7:0]),.ay( 9'sd2),.bx(input_fmap_11[7:0]),.by(-9'sd1),.cx(input_fmap_12[7:0]),.cy( 9'sd2),.dx(input_fmap_14[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O14_N4_S1),.chainout(chainout_4_O14));
logic signed [63:0] chainout_6_O14; 
logic signed [63:0] O14_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O14(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_15[7:0]),.ay(-9'sd2),.bx(input_fmap_16[7:0]),.by(-9'sd2),.cx(input_fmap_17[7:0]),.cy( 9'sd4),.dx(input_fmap_19[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O14_N6_S1),.chainout(chainout_6_O14));
logic signed [63:0] chainout_8_O14; 
logic signed [63:0] O14_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O14(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_25[7:0]),.ay( 9'sd1),.bx(input_fmap_26[7:0]),.by(-9'sd2),.cx(input_fmap_27[7:0]),.cy(-9'sd1),.dx(input_fmap_30[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O14_N8_S1),.chainout(chainout_8_O14));
logic signed [63:0] chainout_10_O14; 
logic signed [63:0] O14_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O14(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_31[7:0]),.ay(-9'sd2),.bx(input_fmap_34[7:0]),.by(-9'sd1),.cx(input_fmap_37[7:0]),.cy(-9'sd2),.dx(input_fmap_40[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O14_N10_S1),.chainout(chainout_10_O14));
logic signed [63:0] chainout_12_O14; 
logic signed [63:0] O14_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O14(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_42[7:0]),.ay( 9'sd1),.bx(input_fmap_43[7:0]),.by(-9'sd1),.cx(input_fmap_45[7:0]),.cy(-9'sd1),.dx(input_fmap_46[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O14_N12_S1),.chainout(chainout_12_O14));
logic signed [63:0] chainout_14_O14; 
logic signed [63:0] O14_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O14(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_48[7:0]),.ay( 9'sd1),.bx(input_fmap_51[7:0]),.by( 9'sd3),.cx(input_fmap_56[7:0]),.cy(-9'sd1),.dx(input_fmap_57[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O14_N14_S1),.chainout(chainout_14_O14));
logic signed [63:0] chainout_16_O14; 
logic signed [63:0] O14_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O14(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_60[7:0]),.ay(-9'sd2),.bx(input_fmap_61[7:0]),.by(-9'sd1),.cx(input_fmap_62[7:0]),.cy(-9'sd2),.dx(input_fmap_63[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O14_N16_S1),.chainout(chainout_16_O14));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O14_N0_S2;		always @(posedge clk) O14_N0_S2 <=     O14_N0_S1  +  O14_N2_S1 ;
 logic signed [21:0] O14_N2_S2;		always @(posedge clk) O14_N2_S2 <=     O14_N4_S1  +  O14_N6_S1 ;
 logic signed [21:0] O14_N4_S2;		always @(posedge clk) O14_N4_S2 <=     O14_N8_S1  +  O14_N10_S1 ;
 logic signed [21:0] O14_N6_S2;		always @(posedge clk) O14_N6_S2 <=     O14_N12_S1  +  O14_N14_S1 ;
 logic signed [21:0] O14_N8_S2;		always @(posedge clk) O14_N8_S2 <=     O14_N16_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O14_N0_S3;		always @(posedge clk) O14_N0_S3 <=     O14_N0_S2  +  O14_N2_S2 ;
 logic signed [22:0] O14_N2_S3;		always @(posedge clk) O14_N2_S3 <=     O14_N4_S2  +  O14_N6_S2 ;
 logic signed [22:0] O14_N4_S3;		always @(posedge clk) O14_N4_S3 <=     O14_N8_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O14_N0_S4;		always @(posedge clk) O14_N0_S4 <=     O14_N0_S3  +  O14_N2_S3 ;
 logic signed [23:0] O14_N2_S4;		always @(posedge clk) O14_N2_S4 <=     O14_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O14_N0_S5;		always @(posedge clk) O14_N0_S5 <=     O14_N0_S4  +  O14_N2_S4 ;
 assign conv_mac_14 = O14_N0_S5;

logic signed [31:0] conv_mac_15;
logic signed [63:0] chainout_0_O15; 
logic signed [63:0] O15_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O15(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_4[7:0]),.ay(-9'sd2),.bx(input_fmap_5[7:0]),.by(-9'sd1),.cx(input_fmap_7[7:0]),.cy(-9'sd1),.dx(input_fmap_21[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O15_N0_S1),.chainout(chainout_0_O15));
logic signed [63:0] chainout_2_O15; 
logic signed [63:0] O15_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O15(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_23[7:0]),.ay(-9'sd1),.bx(input_fmap_31[7:0]),.by(-9'sd1),.cx(input_fmap_35[7:0]),.cy( 9'sd1),.dx(input_fmap_36[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O15_N2_S1),.chainout(chainout_2_O15));
logic signed [63:0] chainout_4_O15; 
logic signed [63:0] O15_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O15(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_47[7:0]),.ay(-9'sd1),.bx(input_fmap_48[7:0]),.by( 9'sd1),.cx(input_fmap_51[7:0]),.cy( 9'sd1),.dx(input_fmap_54[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O15_N4_S1),.chainout(chainout_4_O15));
logic signed [63:0] chainout_6_O15; 
logic signed [63:0] O15_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O15(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_61[7:0]),.ay( 9'sd3),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O15_N6_S1),.chainout(chainout_6_O15));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O15_N0_S2;		always @(posedge clk) O15_N0_S2 <=     O15_N0_S1  +  O15_N2_S1 ;
 logic signed [21:0] O15_N2_S2;		always @(posedge clk) O15_N2_S2 <=     O15_N4_S1  +  O15_N6_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O15_N0_S3;		always @(posedge clk) O15_N0_S3 <=     O15_N0_S2  +  O15_N2_S2 ;
 assign conv_mac_15 = O15_N0_S3;

logic signed [31:0] conv_mac_16;
logic signed [63:0] chainout_0_O16; 
logic signed [63:0] O16_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O16(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd1),.bx(input_fmap_1[7:0]),.by(-9'sd1),.cx(input_fmap_5[7:0]),.cy(-9'sd1),.dx(input_fmap_6[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O16_N0_S1),.chainout(chainout_0_O16));
logic signed [63:0] chainout_2_O16; 
logic signed [63:0] O16_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O16(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_7[7:0]),.ay(-9'sd2),.bx(input_fmap_9[7:0]),.by(-9'sd1),.cx(input_fmap_10[7:0]),.cy( 9'sd1),.dx(input_fmap_11[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O16_N2_S1),.chainout(chainout_2_O16));
logic signed [63:0] chainout_4_O16; 
logic signed [63:0] O16_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O16(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_12[7:0]),.ay( 9'sd1),.bx(input_fmap_13[7:0]),.by(-9'sd1),.cx(input_fmap_15[7:0]),.cy( 9'sd1),.dx(input_fmap_16[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O16_N4_S1),.chainout(chainout_4_O16));
logic signed [63:0] chainout_6_O16; 
logic signed [63:0] O16_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O16(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_17[7:0]),.ay( 9'sd1),.bx(input_fmap_18[7:0]),.by(-9'sd1),.cx(input_fmap_21[7:0]),.cy( 9'sd1),.dx(input_fmap_23[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O16_N6_S1),.chainout(chainout_6_O16));
logic signed [63:0] chainout_8_O16; 
logic signed [63:0] O16_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O16(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_26[7:0]),.ay(-9'sd1),.bx(input_fmap_27[7:0]),.by( 9'sd1),.cx(input_fmap_28[7:0]),.cy(-9'sd1),.dx(input_fmap_31[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O16_N8_S1),.chainout(chainout_8_O16));
logic signed [63:0] chainout_10_O16; 
logic signed [63:0] O16_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O16(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_34[7:0]),.ay(-9'sd1),.bx(input_fmap_35[7:0]),.by(-9'sd1),.cx(input_fmap_37[7:0]),.cy( 9'sd1),.dx(input_fmap_38[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O16_N10_S1),.chainout(chainout_10_O16));
logic signed [63:0] chainout_12_O16; 
logic signed [63:0] O16_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O16(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_39[7:0]),.ay(-9'sd1),.bx(input_fmap_41[7:0]),.by(-9'sd1),.cx(input_fmap_42[7:0]),.cy( 9'sd2),.dx(input_fmap_43[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O16_N12_S1),.chainout(chainout_12_O16));
logic signed [63:0] chainout_14_O16; 
logic signed [63:0] O16_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O16(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_44[7:0]),.ay(-9'sd1),.bx(input_fmap_46[7:0]),.by( 9'sd1),.cx(input_fmap_47[7:0]),.cy(-9'sd1),.dx(input_fmap_48[7:0]),.dy( 9'sd3),.chainin(63'd0),.result(O16_N14_S1),.chainout(chainout_14_O16));
logic signed [63:0] chainout_16_O16; 
logic signed [63:0] O16_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O16(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_49[7:0]),.ay( 9'sd1),.bx(input_fmap_52[7:0]),.by( 9'sd1),.cx(input_fmap_59[7:0]),.cy(-9'sd1),.dx(input_fmap_61[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O16_N16_S1),.chainout(chainout_16_O16));
logic signed [63:0] chainout_18_O16; 
logic signed [63:0] O16_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O16(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_63[7:0]),.ay( 9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O16_N18_S1),.chainout(chainout_18_O16));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O16_N0_S2;		always @(posedge clk) O16_N0_S2 <=     O16_N0_S1  +  O16_N2_S1 ;
 logic signed [21:0] O16_N2_S2;		always @(posedge clk) O16_N2_S2 <=     O16_N4_S1  +  O16_N6_S1 ;
 logic signed [21:0] O16_N4_S2;		always @(posedge clk) O16_N4_S2 <=     O16_N8_S1  +  O16_N10_S1 ;
 logic signed [21:0] O16_N6_S2;		always @(posedge clk) O16_N6_S2 <=     O16_N12_S1  +  O16_N14_S1 ;
 logic signed [21:0] O16_N8_S2;		always @(posedge clk) O16_N8_S2 <=     O16_N16_S1  +  O16_N18_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O16_N0_S3;		always @(posedge clk) O16_N0_S3 <=     O16_N0_S2  +  O16_N2_S2 ;
 logic signed [22:0] O16_N2_S3;		always @(posedge clk) O16_N2_S3 <=     O16_N4_S2  +  O16_N6_S2 ;
 logic signed [22:0] O16_N4_S3;		always @(posedge clk) O16_N4_S3 <=     O16_N8_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O16_N0_S4;		always @(posedge clk) O16_N0_S4 <=     O16_N0_S3  +  O16_N2_S3 ;
 logic signed [23:0] O16_N2_S4;		always @(posedge clk) O16_N2_S4 <=     O16_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O16_N0_S5;		always @(posedge clk) O16_N0_S5 <=     O16_N0_S4  +  O16_N2_S4 ;
 assign conv_mac_16 = O16_N0_S5;

logic signed [31:0] conv_mac_17;
logic signed [63:0] chainout_0_O17; 
logic signed [63:0] O17_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O17(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd1),.bx(input_fmap_2[7:0]),.by(-9'sd1),.cx(input_fmap_3[7:0]),.cy(-9'sd2),.dx(input_fmap_5[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O17_N0_S1),.chainout(chainout_0_O17));
logic signed [63:0] chainout_2_O17; 
logic signed [63:0] O17_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O17(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_6[7:0]),.ay(-9'sd1),.bx(input_fmap_7[7:0]),.by( 9'sd1),.cx(input_fmap_8[7:0]),.cy(-9'sd1),.dx(input_fmap_9[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O17_N2_S1),.chainout(chainout_2_O17));
logic signed [63:0] chainout_4_O17; 
logic signed [63:0] O17_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O17(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_10[7:0]),.ay( 9'sd3),.bx(input_fmap_11[7:0]),.by(-9'sd1),.cx(input_fmap_12[7:0]),.cy( 9'sd1),.dx(input_fmap_16[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O17_N4_S1),.chainout(chainout_4_O17));
logic signed [63:0] chainout_6_O17; 
logic signed [63:0] O17_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O17(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_17[7:0]),.ay( 9'sd1),.bx(input_fmap_19[7:0]),.by(-9'sd1),.cx(input_fmap_21[7:0]),.cy( 9'sd2),.dx(input_fmap_22[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O17_N6_S1),.chainout(chainout_6_O17));
logic signed [63:0] chainout_8_O17; 
logic signed [63:0] O17_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O17(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_25[7:0]),.ay(-9'sd2),.bx(input_fmap_27[7:0]),.by(-9'sd1),.cx(input_fmap_28[7:0]),.cy( 9'sd1),.dx(input_fmap_29[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O17_N8_S1),.chainout(chainout_8_O17));
logic signed [63:0] chainout_10_O17; 
logic signed [63:0] O17_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O17(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_30[7:0]),.ay(-9'sd1),.bx(input_fmap_31[7:0]),.by(-9'sd2),.cx(input_fmap_32[7:0]),.cy( 9'sd2),.dx(input_fmap_33[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O17_N10_S1),.chainout(chainout_10_O17));
logic signed [63:0] chainout_12_O17; 
logic signed [63:0] O17_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O17(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_34[7:0]),.ay( 9'sd1),.bx(input_fmap_35[7:0]),.by( 9'sd1),.cx(input_fmap_37[7:0]),.cy(-9'sd2),.dx(input_fmap_38[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O17_N12_S1),.chainout(chainout_12_O17));
logic signed [63:0] chainout_14_O17; 
logic signed [63:0] O17_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O17(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_39[7:0]),.ay( 9'sd1),.bx(input_fmap_42[7:0]),.by(-9'sd1),.cx(input_fmap_43[7:0]),.cy(-9'sd2),.dx(input_fmap_44[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O17_N14_S1),.chainout(chainout_14_O17));
logic signed [63:0] chainout_16_O17; 
logic signed [63:0] O17_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O17(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_45[7:0]),.ay(-9'sd1),.bx(input_fmap_46[7:0]),.by(-9'sd1),.cx(input_fmap_47[7:0]),.cy(-9'sd1),.dx(input_fmap_48[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O17_N16_S1),.chainout(chainout_16_O17));
logic signed [63:0] chainout_18_O17; 
logic signed [63:0] O17_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O17(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_51[7:0]),.ay( 9'sd2),.bx(input_fmap_52[7:0]),.by( 9'sd1),.cx(input_fmap_56[7:0]),.cy(-9'sd1),.dx(input_fmap_57[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O17_N18_S1),.chainout(chainout_18_O17));
logic signed [63:0] chainout_20_O17; 
logic signed [63:0] O17_N20_S1; 
 int_sop_4_wrapper int_sop_4_inst_20_O17(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_63[7:0]),.ay(-9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O17_N20_S1),.chainout(chainout_20_O17));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O17_N0_S2;		always @(posedge clk) O17_N0_S2 <=     O17_N0_S1  +  O17_N2_S1 ;
 logic signed [21:0] O17_N2_S2;		always @(posedge clk) O17_N2_S2 <=     O17_N4_S1  +  O17_N6_S1 ;
 logic signed [21:0] O17_N4_S2;		always @(posedge clk) O17_N4_S2 <=     O17_N8_S1  +  O17_N10_S1 ;
 logic signed [21:0] O17_N6_S2;		always @(posedge clk) O17_N6_S2 <=     O17_N12_S1  +  O17_N14_S1 ;
 logic signed [21:0] O17_N8_S2;		always @(posedge clk) O17_N8_S2 <=     O17_N16_S1  +  O17_N18_S1 ;
 logic signed [21:0] O17_N10_S2;		always @(posedge clk) O17_N10_S2 <=     O17_N20_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O17_N0_S3;		always @(posedge clk) O17_N0_S3 <=     O17_N0_S2  +  O17_N2_S2 ;
 logic signed [22:0] O17_N2_S3;		always @(posedge clk) O17_N2_S3 <=     O17_N4_S2  +  O17_N6_S2 ;
 logic signed [22:0] O17_N4_S3;		always @(posedge clk) O17_N4_S3 <=     O17_N8_S2  +  O17_N10_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O17_N0_S4;		always @(posedge clk) O17_N0_S4 <=     O17_N0_S3  +  O17_N2_S3 ;
 logic signed [23:0] O17_N2_S4;		always @(posedge clk) O17_N2_S4 <=     O17_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O17_N0_S5;		always @(posedge clk) O17_N0_S5 <=     O17_N0_S4  +  O17_N2_S4 ;
 assign conv_mac_17 = O17_N0_S5;

logic signed [31:0] conv_mac_18;
logic signed [63:0] chainout_0_O18; 
logic signed [63:0] O18_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O18(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd1),.bx(input_fmap_7[7:0]),.by(-9'sd2),.cx(input_fmap_10[7:0]),.cy( 9'sd1),.dx(input_fmap_11[7:0]),.dy( 9'sd3),.chainin(63'd0),.result(O18_N0_S1),.chainout(chainout_0_O18));
logic signed [63:0] chainout_2_O18; 
logic signed [63:0] O18_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O18(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_18[7:0]),.ay(-9'sd1),.bx(input_fmap_31[7:0]),.by(-9'sd1),.cx(input_fmap_35[7:0]),.cy(-9'sd1),.dx(input_fmap_42[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O18_N2_S1),.chainout(chainout_2_O18));
logic signed [63:0] chainout_4_O18; 
logic signed [63:0] O18_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O18(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_43[7:0]),.ay(-9'sd1),.bx(input_fmap_44[7:0]),.by(-9'sd1),.cx(input_fmap_47[7:0]),.cy(-9'sd1),.dx(input_fmap_53[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O18_N4_S1),.chainout(chainout_4_O18));
logic signed [63:0] chainout_6_O18; 
logic signed [63:0] O18_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O18(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_56[7:0]),.ay(-9'sd1),.bx(input_fmap_58[7:0]),.by(-9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O18_N6_S1),.chainout(chainout_6_O18));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O18_N0_S2;		always @(posedge clk) O18_N0_S2 <=     O18_N0_S1  +  O18_N2_S1 ;
 logic signed [21:0] O18_N2_S2;		always @(posedge clk) O18_N2_S2 <=     O18_N4_S1  +  O18_N6_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O18_N0_S3;		always @(posedge clk) O18_N0_S3 <=     O18_N0_S2  +  O18_N2_S2 ;
 assign conv_mac_18 = O18_N0_S3;

logic signed [31:0] conv_mac_19;
logic signed [63:0] chainout_0_O19; 
logic signed [63:0] O19_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O19(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd1),.bx(input_fmap_5[7:0]),.by(-9'sd1),.cx(input_fmap_29[7:0]),.cy(-9'sd1),.dx(input_fmap_35[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O19_N0_S1),.chainout(chainout_0_O19));
logic signed [63:0] chainout_2_O19; 
logic signed [63:0] O19_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O19(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_43[7:0]),.ay( 9'sd1),.bx(input_fmap_44[7:0]),.by(-9'sd1),.cx(input_fmap_46[7:0]),.cy( 9'sd2),.dx(input_fmap_47[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O19_N2_S1),.chainout(chainout_2_O19));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O19_N0_S2;		always @(posedge clk) O19_N0_S2 <=     O19_N0_S1  +  O19_N2_S1 ;
 assign conv_mac_19 = O19_N0_S2;

logic signed [31:0] conv_mac_20;
logic signed [63:0] chainout_0_O20; 
logic signed [63:0] O20_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O20(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_2[7:0]),.ay( 9'sd1),.bx(input_fmap_4[7:0]),.by(-9'sd1),.cx(input_fmap_5[7:0]),.cy(-9'sd1),.dx(input_fmap_6[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O20_N0_S1),.chainout(chainout_0_O20));
logic signed [63:0] chainout_2_O20; 
logic signed [63:0] O20_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O20(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_8[7:0]),.ay( 9'sd1),.bx(input_fmap_10[7:0]),.by(-9'sd1),.cx(input_fmap_12[7:0]),.cy( 9'sd1),.dx(input_fmap_13[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O20_N2_S1),.chainout(chainout_2_O20));
logic signed [63:0] chainout_4_O20; 
logic signed [63:0] O20_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O20(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_14[7:0]),.ay(-9'sd1),.bx(input_fmap_15[7:0]),.by(-9'sd1),.cx(input_fmap_18[7:0]),.cy( 9'sd1),.dx(input_fmap_19[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O20_N4_S1),.chainout(chainout_4_O20));
logic signed [63:0] chainout_6_O20; 
logic signed [63:0] O20_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O20(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_20[7:0]),.ay(-9'sd1),.bx(input_fmap_22[7:0]),.by( 9'sd1),.cx(input_fmap_24[7:0]),.cy(-9'sd6),.dx(input_fmap_28[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O20_N6_S1),.chainout(chainout_6_O20));
logic signed [63:0] chainout_8_O20; 
logic signed [63:0] O20_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O20(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_30[7:0]),.ay( 9'sd2),.bx(input_fmap_31[7:0]),.by( 9'sd1),.cx(input_fmap_33[7:0]),.cy( 9'sd1),.dx(input_fmap_35[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O20_N8_S1),.chainout(chainout_8_O20));
logic signed [63:0] chainout_10_O20; 
logic signed [63:0] O20_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O20(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_36[7:0]),.ay( 9'sd1),.bx(input_fmap_37[7:0]),.by( 9'sd3),.cx(input_fmap_38[7:0]),.cy( 9'sd1),.dx(input_fmap_39[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O20_N10_S1),.chainout(chainout_10_O20));
logic signed [63:0] chainout_12_O20; 
logic signed [63:0] O20_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O20(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_40[7:0]),.ay( 9'sd1),.bx(input_fmap_42[7:0]),.by(-9'sd1),.cx(input_fmap_44[7:0]),.cy(-9'sd1),.dx(input_fmap_45[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O20_N12_S1),.chainout(chainout_12_O20));
logic signed [63:0] chainout_14_O20; 
logic signed [63:0] O20_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O20(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_46[7:0]),.ay(-9'sd1),.bx(input_fmap_51[7:0]),.by( 9'sd1),.cx(input_fmap_55[7:0]),.cy( 9'sd1),.dx(input_fmap_56[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O20_N14_S1),.chainout(chainout_14_O20));
logic signed [63:0] chainout_16_O20; 
logic signed [63:0] O20_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O20(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_57[7:0]),.ay(-9'sd4),.bx(input_fmap_63[7:0]),.by( 9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O20_N16_S1),.chainout(chainout_16_O20));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O20_N0_S2;		always @(posedge clk) O20_N0_S2 <=     O20_N0_S1  +  O20_N2_S1 ;
 logic signed [21:0] O20_N2_S2;		always @(posedge clk) O20_N2_S2 <=     O20_N4_S1  +  O20_N6_S1 ;
 logic signed [21:0] O20_N4_S2;		always @(posedge clk) O20_N4_S2 <=     O20_N8_S1  +  O20_N10_S1 ;
 logic signed [21:0] O20_N6_S2;		always @(posedge clk) O20_N6_S2 <=     O20_N12_S1  +  O20_N14_S1 ;
 logic signed [21:0] O20_N8_S2;		always @(posedge clk) O20_N8_S2 <=     O20_N16_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O20_N0_S3;		always @(posedge clk) O20_N0_S3 <=     O20_N0_S2  +  O20_N2_S2 ;
 logic signed [22:0] O20_N2_S3;		always @(posedge clk) O20_N2_S3 <=     O20_N4_S2  +  O20_N6_S2 ;
 logic signed [22:0] O20_N4_S3;		always @(posedge clk) O20_N4_S3 <=     O20_N8_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O20_N0_S4;		always @(posedge clk) O20_N0_S4 <=     O20_N0_S3  +  O20_N2_S3 ;
 logic signed [23:0] O20_N2_S4;		always @(posedge clk) O20_N2_S4 <=     O20_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O20_N0_S5;		always @(posedge clk) O20_N0_S5 <=     O20_N0_S4  +  O20_N2_S4 ;
 assign conv_mac_20 = O20_N0_S5;

logic signed [31:0] conv_mac_21;
logic signed [63:0] chainout_0_O21; 
logic signed [63:0] O21_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O21(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_7[7:0]),.ay(-9'sd1),.bx(input_fmap_18[7:0]),.by(-9'sd1),.cx(input_fmap_61[7:0]),.cy( 9'sd2),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O21_N0_S1),.chainout(chainout_0_O21));
assign conv_mac_21 = O21_N0_S1;

logic signed [31:0] conv_mac_22;
logic signed [63:0] chainout_0_O22; 
logic signed [63:0] O22_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O22(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd1),.bx(input_fmap_1[7:0]),.by( 9'sd1),.cx(input_fmap_2[7:0]),.cy(-9'sd2),.dx(input_fmap_3[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O22_N0_S1),.chainout(chainout_0_O22));
logic signed [63:0] chainout_2_O22; 
logic signed [63:0] O22_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O22(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_4[7:0]),.ay(-9'sd1),.bx(input_fmap_5[7:0]),.by(-9'sd1),.cx(input_fmap_6[7:0]),.cy( 9'sd1),.dx(input_fmap_8[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O22_N2_S1),.chainout(chainout_2_O22));
logic signed [63:0] chainout_4_O22; 
logic signed [63:0] O22_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O22(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_10[7:0]),.ay(-9'sd2),.bx(input_fmap_12[7:0]),.by(-9'sd1),.cx(input_fmap_13[7:0]),.cy( 9'sd1),.dx(input_fmap_14[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O22_N4_S1),.chainout(chainout_4_O22));
logic signed [63:0] chainout_6_O22; 
logic signed [63:0] O22_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O22(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_15[7:0]),.ay( 9'sd1),.bx(input_fmap_16[7:0]),.by(-9'sd1),.cx(input_fmap_17[7:0]),.cy(-9'sd2),.dx(input_fmap_18[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O22_N6_S1),.chainout(chainout_6_O22));
logic signed [63:0] chainout_8_O22; 
logic signed [63:0] O22_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O22(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_19[7:0]),.ay( 9'sd1),.bx(input_fmap_20[7:0]),.by( 9'sd1),.cx(input_fmap_21[7:0]),.cy( 9'sd3),.dx(input_fmap_22[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O22_N8_S1),.chainout(chainout_8_O22));
logic signed [63:0] chainout_10_O22; 
logic signed [63:0] O22_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O22(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_23[7:0]),.ay( 9'sd1),.bx(input_fmap_26[7:0]),.by( 9'sd1),.cx(input_fmap_27[7:0]),.cy( 9'sd1),.dx(input_fmap_28[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O22_N10_S1),.chainout(chainout_10_O22));
logic signed [63:0] chainout_12_O22; 
logic signed [63:0] O22_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O22(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_29[7:0]),.ay( 9'sd1),.bx(input_fmap_32[7:0]),.by(-9'sd2),.cx(input_fmap_33[7:0]),.cy( 9'sd1),.dx(input_fmap_36[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O22_N12_S1),.chainout(chainout_12_O22));
logic signed [63:0] chainout_14_O22; 
logic signed [63:0] O22_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O22(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_37[7:0]),.ay( 9'sd1),.bx(input_fmap_38[7:0]),.by( 9'sd2),.cx(input_fmap_39[7:0]),.cy(-9'sd1),.dx(input_fmap_43[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O22_N14_S1),.chainout(chainout_14_O22));
logic signed [63:0] chainout_16_O22; 
logic signed [63:0] O22_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O22(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_44[7:0]),.ay( 9'sd1),.bx(input_fmap_45[7:0]),.by(-9'sd1),.cx(input_fmap_46[7:0]),.cy(-9'sd1),.dx(input_fmap_47[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O22_N16_S1),.chainout(chainout_16_O22));
logic signed [63:0] chainout_18_O22; 
logic signed [63:0] O22_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O22(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_50[7:0]),.ay(-9'sd1),.bx(input_fmap_52[7:0]),.by(-9'sd1),.cx(input_fmap_53[7:0]),.cy(-9'sd1),.dx(input_fmap_55[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O22_N18_S1),.chainout(chainout_18_O22));
logic signed [63:0] chainout_20_O22; 
logic signed [63:0] O22_N20_S1; 
 int_sop_4_wrapper int_sop_4_inst_20_O22(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_56[7:0]),.ay( 9'sd1),.bx(input_fmap_57[7:0]),.by( 9'sd1),.cx(input_fmap_58[7:0]),.cy( 9'sd2),.dx(input_fmap_59[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O22_N20_S1),.chainout(chainout_20_O22));
logic signed [63:0] chainout_22_O22; 
logic signed [63:0] O22_N22_S1; 
 int_sop_4_wrapper int_sop_4_inst_22_O22(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_60[7:0]),.ay( 9'sd1),.bx(input_fmap_62[7:0]),.by( 9'sd1),.cx(input_fmap_63[7:0]),.cy( 9'sd3),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O22_N22_S1),.chainout(chainout_22_O22));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O22_N0_S2;		always @(posedge clk) O22_N0_S2 <=     O22_N0_S1  +  O22_N2_S1 ;
 logic signed [21:0] O22_N2_S2;		always @(posedge clk) O22_N2_S2 <=     O22_N4_S1  +  O22_N6_S1 ;
 logic signed [21:0] O22_N4_S2;		always @(posedge clk) O22_N4_S2 <=     O22_N8_S1  +  O22_N10_S1 ;
 logic signed [21:0] O22_N6_S2;		always @(posedge clk) O22_N6_S2 <=     O22_N12_S1  +  O22_N14_S1 ;
 logic signed [21:0] O22_N8_S2;		always @(posedge clk) O22_N8_S2 <=     O22_N16_S1  +  O22_N18_S1 ;
 logic signed [21:0] O22_N10_S2;		always @(posedge clk) O22_N10_S2 <=     O22_N20_S1  +  O22_N22_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O22_N0_S3;		always @(posedge clk) O22_N0_S3 <=     O22_N0_S2  +  O22_N2_S2 ;
 logic signed [22:0] O22_N2_S3;		always @(posedge clk) O22_N2_S3 <=     O22_N4_S2  +  O22_N6_S2 ;
 logic signed [22:0] O22_N4_S3;		always @(posedge clk) O22_N4_S3 <=     O22_N8_S2  +  O22_N10_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O22_N0_S4;		always @(posedge clk) O22_N0_S4 <=     O22_N0_S3  +  O22_N2_S3 ;
 logic signed [23:0] O22_N2_S4;		always @(posedge clk) O22_N2_S4 <=     O22_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O22_N0_S5;		always @(posedge clk) O22_N0_S5 <=     O22_N0_S4  +  O22_N2_S4 ;
 assign conv_mac_22 = O22_N0_S5;

logic signed [31:0] conv_mac_23;
logic signed [63:0] chainout_0_O23; 
logic signed [63:0] O23_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O23(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay( 9'sd1),.bx(input_fmap_2[7:0]),.by(-9'sd2),.cx(input_fmap_5[7:0]),.cy( 9'sd2),.dx(input_fmap_6[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O23_N0_S1),.chainout(chainout_0_O23));
logic signed [63:0] chainout_2_O23; 
logic signed [63:0] O23_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O23(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_7[7:0]),.ay(-9'sd1),.bx(input_fmap_8[7:0]),.by( 9'sd3),.cx(input_fmap_10[7:0]),.cy(-9'sd1),.dx(input_fmap_11[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O23_N2_S1),.chainout(chainout_2_O23));
logic signed [63:0] chainout_4_O23; 
logic signed [63:0] O23_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O23(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_12[7:0]),.ay(-9'sd1),.bx(input_fmap_13[7:0]),.by( 9'sd2),.cx(input_fmap_14[7:0]),.cy(-9'sd2),.dx(input_fmap_15[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O23_N4_S1),.chainout(chainout_4_O23));
logic signed [63:0] chainout_6_O23; 
logic signed [63:0] O23_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O23(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_17[7:0]),.ay(-9'sd2),.bx(input_fmap_18[7:0]),.by( 9'sd1),.cx(input_fmap_19[7:0]),.cy( 9'sd2),.dx(input_fmap_20[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O23_N6_S1),.chainout(chainout_6_O23));
logic signed [63:0] chainout_8_O23; 
logic signed [63:0] O23_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O23(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_22[7:0]),.ay(-9'sd1),.bx(input_fmap_29[7:0]),.by( 9'sd1),.cx(input_fmap_30[7:0]),.cy(-9'sd2),.dx(input_fmap_31[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O23_N8_S1),.chainout(chainout_8_O23));
logic signed [63:0] chainout_10_O23; 
logic signed [63:0] O23_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O23(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_32[7:0]),.ay(-9'sd2),.bx(input_fmap_33[7:0]),.by( 9'sd1),.cx(input_fmap_34[7:0]),.cy(-9'sd1),.dx(input_fmap_35[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O23_N10_S1),.chainout(chainout_10_O23));
logic signed [63:0] chainout_12_O23; 
logic signed [63:0] O23_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O23(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_36[7:0]),.ay(-9'sd2),.bx(input_fmap_40[7:0]),.by(-9'sd1),.cx(input_fmap_41[7:0]),.cy(-9'sd3),.dx(input_fmap_42[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O23_N12_S1),.chainout(chainout_12_O23));
logic signed [63:0] chainout_14_O23; 
logic signed [63:0] O23_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O23(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_45[7:0]),.ay( 9'sd1),.bx(input_fmap_46[7:0]),.by( 9'sd2),.cx(input_fmap_47[7:0]),.cy( 9'sd1),.dx(input_fmap_48[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O23_N14_S1),.chainout(chainout_14_O23));
logic signed [63:0] chainout_16_O23; 
logic signed [63:0] O23_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O23(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_49[7:0]),.ay( 9'sd1),.bx(input_fmap_50[7:0]),.by( 9'sd1),.cx(input_fmap_52[7:0]),.cy(-9'sd2),.dx(input_fmap_53[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O23_N16_S1),.chainout(chainout_16_O23));
logic signed [63:0] chainout_18_O23; 
logic signed [63:0] O23_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O23(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_54[7:0]),.ay(-9'sd1),.bx(input_fmap_55[7:0]),.by( 9'sd1),.cx(input_fmap_56[7:0]),.cy(-9'sd1),.dx(input_fmap_59[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O23_N18_S1),.chainout(chainout_18_O23));
logic signed [63:0] chainout_20_O23; 
logic signed [63:0] O23_N20_S1; 
 int_sop_4_wrapper int_sop_4_inst_20_O23(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_60[7:0]),.ay( 9'sd2),.bx(input_fmap_63[7:0]),.by( 9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O23_N20_S1),.chainout(chainout_20_O23));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O23_N0_S2;		always @(posedge clk) O23_N0_S2 <=     O23_N0_S1  +  O23_N2_S1 ;
 logic signed [21:0] O23_N2_S2;		always @(posedge clk) O23_N2_S2 <=     O23_N4_S1  +  O23_N6_S1 ;
 logic signed [21:0] O23_N4_S2;		always @(posedge clk) O23_N4_S2 <=     O23_N8_S1  +  O23_N10_S1 ;
 logic signed [21:0] O23_N6_S2;		always @(posedge clk) O23_N6_S2 <=     O23_N12_S1  +  O23_N14_S1 ;
 logic signed [21:0] O23_N8_S2;		always @(posedge clk) O23_N8_S2 <=     O23_N16_S1  +  O23_N18_S1 ;
 logic signed [21:0] O23_N10_S2;		always @(posedge clk) O23_N10_S2 <=     O23_N20_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O23_N0_S3;		always @(posedge clk) O23_N0_S3 <=     O23_N0_S2  +  O23_N2_S2 ;
 logic signed [22:0] O23_N2_S3;		always @(posedge clk) O23_N2_S3 <=     O23_N4_S2  +  O23_N6_S2 ;
 logic signed [22:0] O23_N4_S3;		always @(posedge clk) O23_N4_S3 <=     O23_N8_S2  +  O23_N10_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O23_N0_S4;		always @(posedge clk) O23_N0_S4 <=     O23_N0_S3  +  O23_N2_S3 ;
 logic signed [23:0] O23_N2_S4;		always @(posedge clk) O23_N2_S4 <=     O23_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O23_N0_S5;		always @(posedge clk) O23_N0_S5 <=     O23_N0_S4  +  O23_N2_S4 ;
 assign conv_mac_23 = O23_N0_S5;

logic signed [31:0] conv_mac_24;
logic signed [63:0] chainout_0_O24; 
logic signed [63:0] O24_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O24(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd3),.bx(input_fmap_2[7:0]),.by( 9'sd3),.cx(input_fmap_3[7:0]),.cy(-9'sd3),.dx(input_fmap_5[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O24_N0_S1),.chainout(chainout_0_O24));
logic signed [63:0] chainout_2_O24; 
logic signed [63:0] O24_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O24(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_6[7:0]),.ay( 9'sd2),.bx(input_fmap_7[7:0]),.by(-9'sd1),.cx(input_fmap_8[7:0]),.cy(-9'sd1),.dx(input_fmap_9[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O24_N2_S1),.chainout(chainout_2_O24));
logic signed [63:0] chainout_4_O24; 
logic signed [63:0] O24_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O24(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_11[7:0]),.ay(-9'sd4),.bx(input_fmap_12[7:0]),.by(-9'sd2),.cx(input_fmap_13[7:0]),.cy(-9'sd3),.dx(input_fmap_14[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O24_N4_S1),.chainout(chainout_4_O24));
logic signed [63:0] chainout_6_O24; 
logic signed [63:0] O24_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O24(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_15[7:0]),.ay(-9'sd3),.bx(input_fmap_16[7:0]),.by(-9'sd1),.cx(input_fmap_18[7:0]),.cy(-9'sd2),.dx(input_fmap_19[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O24_N6_S1),.chainout(chainout_6_O24));
logic signed [63:0] chainout_8_O24; 
logic signed [63:0] O24_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O24(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_20[7:0]),.ay( 9'sd2),.bx(input_fmap_21[7:0]),.by( 9'sd1),.cx(input_fmap_23[7:0]),.cy(-9'sd2),.dx(input_fmap_24[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O24_N8_S1),.chainout(chainout_8_O24));
logic signed [63:0] chainout_10_O24; 
logic signed [63:0] O24_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O24(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_25[7:0]),.ay(-9'sd1),.bx(input_fmap_26[7:0]),.by( 9'sd2),.cx(input_fmap_27[7:0]),.cy(-9'sd2),.dx(input_fmap_28[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O24_N10_S1),.chainout(chainout_10_O24));
logic signed [63:0] chainout_12_O24; 
logic signed [63:0] O24_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O24(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_30[7:0]),.ay( 9'sd1),.bx(input_fmap_31[7:0]),.by( 9'sd2),.cx(input_fmap_32[7:0]),.cy(-9'sd2),.dx(input_fmap_33[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O24_N12_S1),.chainout(chainout_12_O24));
logic signed [63:0] chainout_14_O24; 
logic signed [63:0] O24_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O24(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_34[7:0]),.ay(-9'sd3),.bx(input_fmap_35[7:0]),.by(-9'sd2),.cx(input_fmap_36[7:0]),.cy( 9'sd2),.dx(input_fmap_38[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O24_N14_S1),.chainout(chainout_14_O24));
logic signed [63:0] chainout_16_O24; 
logic signed [63:0] O24_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O24(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_39[7:0]),.ay( 9'sd2),.bx(input_fmap_40[7:0]),.by( 9'sd2),.cx(input_fmap_41[7:0]),.cy(-9'sd1),.dx(input_fmap_42[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O24_N16_S1),.chainout(chainout_16_O24));
logic signed [63:0] chainout_18_O24; 
logic signed [63:0] O24_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O24(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_46[7:0]),.ay(-9'sd3),.bx(input_fmap_47[7:0]),.by( 9'sd1),.cx(input_fmap_48[7:0]),.cy( 9'sd1),.dx(input_fmap_49[7:0]),.dy( 9'sd3),.chainin(63'd0),.result(O24_N18_S1),.chainout(chainout_18_O24));
logic signed [63:0] chainout_20_O24; 
logic signed [63:0] O24_N20_S1; 
 int_sop_4_wrapper int_sop_4_inst_20_O24(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_50[7:0]),.ay(-9'sd3),.bx(input_fmap_51[7:0]),.by( 9'sd1),.cx(input_fmap_52[7:0]),.cy( 9'sd3),.dx(input_fmap_53[7:0]),.dy( 9'sd6),.chainin(63'd0),.result(O24_N20_S1),.chainout(chainout_20_O24));
logic signed [63:0] chainout_22_O24; 
logic signed [63:0] O24_N22_S1; 
 int_sop_4_wrapper int_sop_4_inst_22_O24(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_54[7:0]),.ay(-9'sd1),.bx(input_fmap_56[7:0]),.by( 9'sd2),.cx(input_fmap_58[7:0]),.cy(-9'sd1),.dx(input_fmap_59[7:0]),.dy( 9'sd4),.chainin(63'd0),.result(O24_N22_S1),.chainout(chainout_22_O24));
logic signed [63:0] chainout_24_O24; 
logic signed [63:0] O24_N24_S1; 
 int_sop_4_wrapper int_sop_4_inst_24_O24(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_61[7:0]),.ay(-9'sd2),.bx(input_fmap_62[7:0]),.by( 9'sd1),.cx(input_fmap_63[7:0]),.cy(-9'sd2),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O24_N24_S1),.chainout(chainout_24_O24));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O24_N0_S2;		always @(posedge clk) O24_N0_S2 <=     O24_N0_S1  +  O24_N2_S1 ;
 logic signed [21:0] O24_N2_S2;		always @(posedge clk) O24_N2_S2 <=     O24_N4_S1  +  O24_N6_S1 ;
 logic signed [21:0] O24_N4_S2;		always @(posedge clk) O24_N4_S2 <=     O24_N8_S1  +  O24_N10_S1 ;
 logic signed [21:0] O24_N6_S2;		always @(posedge clk) O24_N6_S2 <=     O24_N12_S1  +  O24_N14_S1 ;
 logic signed [21:0] O24_N8_S2;		always @(posedge clk) O24_N8_S2 <=     O24_N16_S1  +  O24_N18_S1 ;
 logic signed [21:0] O24_N10_S2;		always @(posedge clk) O24_N10_S2 <=     O24_N20_S1  +  O24_N22_S1 ;
 logic signed [21:0] O24_N12_S2;		always @(posedge clk) O24_N12_S2 <=     O24_N24_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O24_N0_S3;		always @(posedge clk) O24_N0_S3 <=     O24_N0_S2  +  O24_N2_S2 ;
 logic signed [22:0] O24_N2_S3;		always @(posedge clk) O24_N2_S3 <=     O24_N4_S2  +  O24_N6_S2 ;
 logic signed [22:0] O24_N4_S3;		always @(posedge clk) O24_N4_S3 <=     O24_N8_S2  +  O24_N10_S2 ;
 logic signed [22:0] O24_N6_S3;		always @(posedge clk) O24_N6_S3 <=     O24_N12_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O24_N0_S4;		always @(posedge clk) O24_N0_S4 <=     O24_N0_S3  +  O24_N2_S3 ;
 logic signed [23:0] O24_N2_S4;		always @(posedge clk) O24_N2_S4 <=     O24_N4_S3  +  O24_N6_S3 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O24_N0_S5;		always @(posedge clk) O24_N0_S5 <=     O24_N0_S4  +  O24_N2_S4 ;
 assign conv_mac_24 = O24_N0_S5;

logic signed [31:0] conv_mac_25;
logic signed [63:0] chainout_0_O25; 
logic signed [63:0] O25_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O25(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd2),.bx(input_fmap_1[7:0]),.by( 9'sd1),.cx(input_fmap_3[7:0]),.cy( 9'sd1),.dx(input_fmap_4[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O25_N0_S1),.chainout(chainout_0_O25));
logic signed [63:0] chainout_2_O25; 
logic signed [63:0] O25_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O25(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_6[7:0]),.ay( 9'sd1),.bx(input_fmap_7[7:0]),.by( 9'sd1),.cx(input_fmap_9[7:0]),.cy( 9'sd1),.dx(input_fmap_10[7:0]),.dy(-9'sd4),.chainin(63'd0),.result(O25_N2_S1),.chainout(chainout_2_O25));
logic signed [63:0] chainout_4_O25; 
logic signed [63:0] O25_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O25(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_11[7:0]),.ay(-9'sd1),.bx(input_fmap_13[7:0]),.by(-9'sd1),.cx(input_fmap_15[7:0]),.cy( 9'sd1),.dx(input_fmap_18[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O25_N4_S1),.chainout(chainout_4_O25));
logic signed [63:0] chainout_6_O25; 
logic signed [63:0] O25_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O25(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_20[7:0]),.ay(-9'sd1),.bx(input_fmap_21[7:0]),.by( 9'sd1),.cx(input_fmap_22[7:0]),.cy(-9'sd1),.dx(input_fmap_23[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O25_N6_S1),.chainout(chainout_6_O25));
logic signed [63:0] chainout_8_O25; 
logic signed [63:0] O25_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O25(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_24[7:0]),.ay(-9'sd1),.bx(input_fmap_27[7:0]),.by( 9'sd1),.cx(input_fmap_28[7:0]),.cy(-9'sd1),.dx(input_fmap_30[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O25_N8_S1),.chainout(chainout_8_O25));
logic signed [63:0] chainout_10_O25; 
logic signed [63:0] O25_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O25(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_31[7:0]),.ay(-9'sd2),.bx(input_fmap_32[7:0]),.by(-9'sd1),.cx(input_fmap_33[7:0]),.cy(-9'sd1),.dx(input_fmap_34[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O25_N10_S1),.chainout(chainout_10_O25));
logic signed [63:0] chainout_12_O25; 
logic signed [63:0] O25_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O25(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_37[7:0]),.ay(-9'sd1),.bx(input_fmap_39[7:0]),.by(-9'sd1),.cx(input_fmap_42[7:0]),.cy( 9'sd2),.dx(input_fmap_43[7:0]),.dy( 9'sd3),.chainin(63'd0),.result(O25_N12_S1),.chainout(chainout_12_O25));
logic signed [63:0] chainout_14_O25; 
logic signed [63:0] O25_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O25(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_44[7:0]),.ay(-9'sd6),.bx(input_fmap_45[7:0]),.by( 9'sd1),.cx(input_fmap_47[7:0]),.cy( 9'sd1),.dx(input_fmap_48[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O25_N14_S1),.chainout(chainout_14_O25));
logic signed [63:0] chainout_16_O25; 
logic signed [63:0] O25_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O25(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_51[7:0]),.ay(-9'sd1),.bx(input_fmap_52[7:0]),.by(-9'sd1),.cx(input_fmap_54[7:0]),.cy(-9'sd1),.dx(input_fmap_55[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O25_N16_S1),.chainout(chainout_16_O25));
logic signed [63:0] chainout_18_O25; 
logic signed [63:0] O25_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O25(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_56[7:0]),.ay(-9'sd1),.bx(input_fmap_58[7:0]),.by( 9'sd3),.cx(input_fmap_60[7:0]),.cy(-9'sd1),.dx(input_fmap_62[7:0]),.dy(-9'sd3),.chainin(63'd0),.result(O25_N18_S1),.chainout(chainout_18_O25));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O25_N0_S2;		always @(posedge clk) O25_N0_S2 <=     O25_N0_S1  +  O25_N2_S1 ;
 logic signed [21:0] O25_N2_S2;		always @(posedge clk) O25_N2_S2 <=     O25_N4_S1  +  O25_N6_S1 ;
 logic signed [21:0] O25_N4_S2;		always @(posedge clk) O25_N4_S2 <=     O25_N8_S1  +  O25_N10_S1 ;
 logic signed [21:0] O25_N6_S2;		always @(posedge clk) O25_N6_S2 <=     O25_N12_S1  +  O25_N14_S1 ;
 logic signed [21:0] O25_N8_S2;		always @(posedge clk) O25_N8_S2 <=     O25_N16_S1  +  O25_N18_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O25_N0_S3;		always @(posedge clk) O25_N0_S3 <=     O25_N0_S2  +  O25_N2_S2 ;
 logic signed [22:0] O25_N2_S3;		always @(posedge clk) O25_N2_S3 <=     O25_N4_S2  +  O25_N6_S2 ;
 logic signed [22:0] O25_N4_S3;		always @(posedge clk) O25_N4_S3 <=     O25_N8_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O25_N0_S4;		always @(posedge clk) O25_N0_S4 <=     O25_N0_S3  +  O25_N2_S3 ;
 logic signed [23:0] O25_N2_S4;		always @(posedge clk) O25_N2_S4 <=     O25_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O25_N0_S5;		always @(posedge clk) O25_N0_S5 <=     O25_N0_S4  +  O25_N2_S4 ;
 assign conv_mac_25 = O25_N0_S5;

logic signed [31:0] conv_mac_26;
logic signed [63:0] chainout_0_O26; 
logic signed [63:0] O26_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O26(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd1),.bx(input_fmap_2[7:0]),.by( 9'sd1),.cx(input_fmap_4[7:0]),.cy(-9'sd1),.dx(input_fmap_6[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O26_N0_S1),.chainout(chainout_0_O26));
logic signed [63:0] chainout_2_O26; 
logic signed [63:0] O26_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O26(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_7[7:0]),.ay( 9'sd1),.bx(input_fmap_8[7:0]),.by( 9'sd1),.cx(input_fmap_10[7:0]),.cy( 9'sd3),.dx(input_fmap_11[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O26_N2_S1),.chainout(chainout_2_O26));
logic signed [63:0] chainout_4_O26; 
logic signed [63:0] O26_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O26(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_13[7:0]),.ay(-9'sd1),.bx(input_fmap_14[7:0]),.by(-9'sd1),.cx(input_fmap_16[7:0]),.cy(-9'sd1),.dx(input_fmap_17[7:0]),.dy(-9'sd3),.chainin(63'd0),.result(O26_N4_S1),.chainout(chainout_4_O26));
logic signed [63:0] chainout_6_O26; 
logic signed [63:0] O26_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O26(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_18[7:0]),.ay(-9'sd1),.bx(input_fmap_19[7:0]),.by( 9'sd2),.cx(input_fmap_20[7:0]),.cy( 9'sd1),.dx(input_fmap_21[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O26_N6_S1),.chainout(chainout_6_O26));
logic signed [63:0] chainout_8_O26; 
logic signed [63:0] O26_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O26(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_22[7:0]),.ay(-9'sd1),.bx(input_fmap_25[7:0]),.by( 9'sd1),.cx(input_fmap_26[7:0]),.cy( 9'sd1),.dx(input_fmap_27[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O26_N8_S1),.chainout(chainout_8_O26));
logic signed [63:0] chainout_10_O26; 
logic signed [63:0] O26_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O26(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_28[7:0]),.ay(-9'sd2),.bx(input_fmap_29[7:0]),.by( 9'sd1),.cx(input_fmap_33[7:0]),.cy( 9'sd1),.dx(input_fmap_34[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O26_N10_S1),.chainout(chainout_10_O26));
logic signed [63:0] chainout_12_O26; 
logic signed [63:0] O26_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O26(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_36[7:0]),.ay(-9'sd1),.bx(input_fmap_37[7:0]),.by(-9'sd1),.cx(input_fmap_40[7:0]),.cy( 9'sd1),.dx(input_fmap_41[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O26_N12_S1),.chainout(chainout_12_O26));
logic signed [63:0] chainout_14_O26; 
logic signed [63:0] O26_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O26(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_42[7:0]),.ay( 9'sd1),.bx(input_fmap_43[7:0]),.by(-9'sd1),.cx(input_fmap_44[7:0]),.cy( 9'sd2),.dx(input_fmap_46[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O26_N14_S1),.chainout(chainout_14_O26));
logic signed [63:0] chainout_16_O26; 
logic signed [63:0] O26_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O26(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_47[7:0]),.ay( 9'sd1),.bx(input_fmap_48[7:0]),.by( 9'sd1),.cx(input_fmap_49[7:0]),.cy(-9'sd1),.dx(input_fmap_54[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O26_N16_S1),.chainout(chainout_16_O26));
logic signed [63:0] chainout_18_O26; 
logic signed [63:0] O26_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O26(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_55[7:0]),.ay( 9'sd1),.bx(input_fmap_57[7:0]),.by(-9'sd1),.cx(input_fmap_59[7:0]),.cy(-9'sd2),.dx(input_fmap_61[7:0]),.dy( 9'sd3),.chainin(63'd0),.result(O26_N18_S1),.chainout(chainout_18_O26));
logic signed [63:0] chainout_20_O26; 
logic signed [63:0] O26_N20_S1; 
 int_sop_4_wrapper int_sop_4_inst_20_O26(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_62[7:0]),.ay( 9'sd4),.bx(input_fmap_63[7:0]),.by(-9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O26_N20_S1),.chainout(chainout_20_O26));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O26_N0_S2;		always @(posedge clk) O26_N0_S2 <=     O26_N0_S1  +  O26_N2_S1 ;
 logic signed [21:0] O26_N2_S2;		always @(posedge clk) O26_N2_S2 <=     O26_N4_S1  +  O26_N6_S1 ;
 logic signed [21:0] O26_N4_S2;		always @(posedge clk) O26_N4_S2 <=     O26_N8_S1  +  O26_N10_S1 ;
 logic signed [21:0] O26_N6_S2;		always @(posedge clk) O26_N6_S2 <=     O26_N12_S1  +  O26_N14_S1 ;
 logic signed [21:0] O26_N8_S2;		always @(posedge clk) O26_N8_S2 <=     O26_N16_S1  +  O26_N18_S1 ;
 logic signed [21:0] O26_N10_S2;		always @(posedge clk) O26_N10_S2 <=     O26_N20_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O26_N0_S3;		always @(posedge clk) O26_N0_S3 <=     O26_N0_S2  +  O26_N2_S2 ;
 logic signed [22:0] O26_N2_S3;		always @(posedge clk) O26_N2_S3 <=     O26_N4_S2  +  O26_N6_S2 ;
 logic signed [22:0] O26_N4_S3;		always @(posedge clk) O26_N4_S3 <=     O26_N8_S2  +  O26_N10_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O26_N0_S4;		always @(posedge clk) O26_N0_S4 <=     O26_N0_S3  +  O26_N2_S3 ;
 logic signed [23:0] O26_N2_S4;		always @(posedge clk) O26_N2_S4 <=     O26_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O26_N0_S5;		always @(posedge clk) O26_N0_S5 <=     O26_N0_S4  +  O26_N2_S4 ;
 assign conv_mac_26 = O26_N0_S5;

logic signed [31:0] conv_mac_27;
logic signed [63:0] chainout_0_O27; 
logic signed [63:0] O27_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O27(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_3[7:0]),.ay(-9'sd3),.bx(input_fmap_4[7:0]),.by( 9'sd1),.cx(input_fmap_5[7:0]),.cy(-9'sd3),.dx(input_fmap_6[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O27_N0_S1),.chainout(chainout_0_O27));
logic signed [63:0] chainout_2_O27; 
logic signed [63:0] O27_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O27(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_10[7:0]),.ay( 9'sd1),.bx(input_fmap_11[7:0]),.by(-9'sd1),.cx(input_fmap_13[7:0]),.cy( 9'sd1),.dx(input_fmap_14[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O27_N2_S1),.chainout(chainout_2_O27));
logic signed [63:0] chainout_4_O27; 
logic signed [63:0] O27_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O27(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_15[7:0]),.ay(-9'sd1),.bx(input_fmap_18[7:0]),.by( 9'sd1),.cx(input_fmap_21[7:0]),.cy( 9'sd1),.dx(input_fmap_25[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O27_N4_S1),.chainout(chainout_4_O27));
logic signed [63:0] chainout_6_O27; 
logic signed [63:0] O27_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O27(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_26[7:0]),.ay( 9'sd3),.bx(input_fmap_27[7:0]),.by(-9'sd1),.cx(input_fmap_28[7:0]),.cy(-9'sd1),.dx(input_fmap_34[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O27_N6_S1),.chainout(chainout_6_O27));
logic signed [63:0] chainout_8_O27; 
logic signed [63:0] O27_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O27(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_35[7:0]),.ay(-9'sd1),.bx(input_fmap_36[7:0]),.by(-9'sd1),.cx(input_fmap_37[7:0]),.cy( 9'sd2),.dx(input_fmap_38[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O27_N8_S1),.chainout(chainout_8_O27));
logic signed [63:0] chainout_10_O27; 
logic signed [63:0] O27_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O27(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_41[7:0]),.ay( 9'sd1),.bx(input_fmap_42[7:0]),.by(-9'sd1),.cx(input_fmap_46[7:0]),.cy(-9'sd2),.dx(input_fmap_48[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O27_N10_S1),.chainout(chainout_10_O27));
logic signed [63:0] chainout_12_O27; 
logic signed [63:0] O27_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O27(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_50[7:0]),.ay(-9'sd2),.bx(input_fmap_51[7:0]),.by(-9'sd1),.cx(input_fmap_52[7:0]),.cy(-9'sd1),.dx(input_fmap_53[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O27_N12_S1),.chainout(chainout_12_O27));
logic signed [63:0] chainout_14_O27; 
logic signed [63:0] O27_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O27(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_55[7:0]),.ay( 9'sd1),.bx(input_fmap_56[7:0]),.by(-9'sd1),.cx(input_fmap_57[7:0]),.cy(-9'sd1),.dx(input_fmap_59[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O27_N14_S1),.chainout(chainout_14_O27));
logic signed [63:0] chainout_16_O27; 
logic signed [63:0] O27_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O27(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_60[7:0]),.ay( 9'sd1),.bx(input_fmap_63[7:0]),.by( 9'sd2),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O27_N16_S1),.chainout(chainout_16_O27));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O27_N0_S2;		always @(posedge clk) O27_N0_S2 <=     O27_N0_S1  +  O27_N2_S1 ;
 logic signed [21:0] O27_N2_S2;		always @(posedge clk) O27_N2_S2 <=     O27_N4_S1  +  O27_N6_S1 ;
 logic signed [21:0] O27_N4_S2;		always @(posedge clk) O27_N4_S2 <=     O27_N8_S1  +  O27_N10_S1 ;
 logic signed [21:0] O27_N6_S2;		always @(posedge clk) O27_N6_S2 <=     O27_N12_S1  +  O27_N14_S1 ;
 logic signed [21:0] O27_N8_S2;		always @(posedge clk) O27_N8_S2 <=     O27_N16_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O27_N0_S3;		always @(posedge clk) O27_N0_S3 <=     O27_N0_S2  +  O27_N2_S2 ;
 logic signed [22:0] O27_N2_S3;		always @(posedge clk) O27_N2_S3 <=     O27_N4_S2  +  O27_N6_S2 ;
 logic signed [22:0] O27_N4_S3;		always @(posedge clk) O27_N4_S3 <=     O27_N8_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O27_N0_S4;		always @(posedge clk) O27_N0_S4 <=     O27_N0_S3  +  O27_N2_S3 ;
 logic signed [23:0] O27_N2_S4;		always @(posedge clk) O27_N2_S4 <=     O27_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O27_N0_S5;		always @(posedge clk) O27_N0_S5 <=     O27_N0_S4  +  O27_N2_S4 ;
 assign conv_mac_27 = O27_N0_S5;

logic signed [31:0] conv_mac_28;
logic signed [63:0] chainout_0_O28; 
logic signed [63:0] O28_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O28(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd4),.bx(input_fmap_1[7:0]),.by(-9'sd3),.cx(input_fmap_2[7:0]),.cy( 9'sd5),.dx(input_fmap_8[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O28_N0_S1),.chainout(chainout_0_O28));
logic signed [63:0] chainout_2_O28; 
logic signed [63:0] O28_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O28(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_10[7:0]),.ay(-9'sd1),.bx(input_fmap_11[7:0]),.by( 9'sd2),.cx(input_fmap_14[7:0]),.cy( 9'sd1),.dx(input_fmap_16[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O28_N2_S1),.chainout(chainout_2_O28));
logic signed [63:0] chainout_4_O28; 
logic signed [63:0] O28_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O28(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_18[7:0]),.ay(-9'sd2),.bx(input_fmap_19[7:0]),.by(-9'sd1),.cx(input_fmap_20[7:0]),.cy( 9'sd1),.dx(input_fmap_21[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O28_N4_S1),.chainout(chainout_4_O28));
logic signed [63:0] chainout_6_O28; 
logic signed [63:0] O28_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O28(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_22[7:0]),.ay( 9'sd2),.bx(input_fmap_24[7:0]),.by(-9'sd1),.cx(input_fmap_25[7:0]),.cy( 9'sd1),.dx(input_fmap_26[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O28_N6_S1),.chainout(chainout_6_O28));
logic signed [63:0] chainout_8_O28; 
logic signed [63:0] O28_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O28(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_27[7:0]),.ay(-9'sd1),.bx(input_fmap_28[7:0]),.by( 9'sd1),.cx(input_fmap_29[7:0]),.cy(-9'sd1),.dx(input_fmap_30[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O28_N8_S1),.chainout(chainout_8_O28));
logic signed [63:0] chainout_10_O28; 
logic signed [63:0] O28_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O28(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_31[7:0]),.ay(-9'sd1),.bx(input_fmap_32[7:0]),.by( 9'sd2),.cx(input_fmap_33[7:0]),.cy( 9'sd1),.dx(input_fmap_34[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O28_N10_S1),.chainout(chainout_10_O28));
logic signed [63:0] chainout_12_O28; 
logic signed [63:0] O28_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O28(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_35[7:0]),.ay(-9'sd1),.bx(input_fmap_36[7:0]),.by( 9'sd1),.cx(input_fmap_37[7:0]),.cy(-9'sd1),.dx(input_fmap_39[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O28_N12_S1),.chainout(chainout_12_O28));
logic signed [63:0] chainout_14_O28; 
logic signed [63:0] O28_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O28(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_41[7:0]),.ay(-9'sd1),.bx(input_fmap_43[7:0]),.by( 9'sd1),.cx(input_fmap_44[7:0]),.cy(-9'sd1),.dx(input_fmap_45[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O28_N14_S1),.chainout(chainout_14_O28));
logic signed [63:0] chainout_16_O28; 
logic signed [63:0] O28_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O28(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_46[7:0]),.ay( 9'sd3),.bx(input_fmap_47[7:0]),.by(-9'sd1),.cx(input_fmap_48[7:0]),.cy( 9'sd1),.dx(input_fmap_50[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O28_N16_S1),.chainout(chainout_16_O28));
logic signed [63:0] chainout_18_O28; 
logic signed [63:0] O28_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O28(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_51[7:0]),.ay( 9'sd3),.bx(input_fmap_52[7:0]),.by(-9'sd2),.cx(input_fmap_53[7:0]),.cy(-9'sd1),.dx(input_fmap_54[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O28_N18_S1),.chainout(chainout_18_O28));
logic signed [63:0] chainout_20_O28; 
logic signed [63:0] O28_N20_S1; 
 int_sop_4_wrapper int_sop_4_inst_20_O28(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_55[7:0]),.ay(-9'sd1),.bx(input_fmap_56[7:0]),.by( 9'sd1),.cx(input_fmap_57[7:0]),.cy(-9'sd1),.dx(input_fmap_58[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O28_N20_S1),.chainout(chainout_20_O28));
logic signed [63:0] chainout_22_O28; 
logic signed [63:0] O28_N22_S1; 
 int_sop_4_wrapper int_sop_4_inst_22_O28(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_59[7:0]),.ay(-9'sd1),.bx(input_fmap_62[7:0]),.by( 9'sd1),.cx(input_fmap_63[7:0]),.cy(-9'sd1),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O28_N22_S1),.chainout(chainout_22_O28));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O28_N0_S2;		always @(posedge clk) O28_N0_S2 <=     O28_N0_S1  +  O28_N2_S1 ;
 logic signed [21:0] O28_N2_S2;		always @(posedge clk) O28_N2_S2 <=     O28_N4_S1  +  O28_N6_S1 ;
 logic signed [21:0] O28_N4_S2;		always @(posedge clk) O28_N4_S2 <=     O28_N8_S1  +  O28_N10_S1 ;
 logic signed [21:0] O28_N6_S2;		always @(posedge clk) O28_N6_S2 <=     O28_N12_S1  +  O28_N14_S1 ;
 logic signed [21:0] O28_N8_S2;		always @(posedge clk) O28_N8_S2 <=     O28_N16_S1  +  O28_N18_S1 ;
 logic signed [21:0] O28_N10_S2;		always @(posedge clk) O28_N10_S2 <=     O28_N20_S1  +  O28_N22_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O28_N0_S3;		always @(posedge clk) O28_N0_S3 <=     O28_N0_S2  +  O28_N2_S2 ;
 logic signed [22:0] O28_N2_S3;		always @(posedge clk) O28_N2_S3 <=     O28_N4_S2  +  O28_N6_S2 ;
 logic signed [22:0] O28_N4_S3;		always @(posedge clk) O28_N4_S3 <=     O28_N8_S2  +  O28_N10_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O28_N0_S4;		always @(posedge clk) O28_N0_S4 <=     O28_N0_S3  +  O28_N2_S3 ;
 logic signed [23:0] O28_N2_S4;		always @(posedge clk) O28_N2_S4 <=     O28_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O28_N0_S5;		always @(posedge clk) O28_N0_S5 <=     O28_N0_S4  +  O28_N2_S4 ;
 assign conv_mac_28 = O28_N0_S5;

logic signed [31:0] conv_mac_29;
logic signed [63:0] chainout_0_O29; 
logic signed [63:0] O29_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O29(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay(-9'sd1),.bx(input_fmap_3[7:0]),.by(-9'sd1),.cx(input_fmap_4[7:0]),.cy(-9'sd1),.dx(input_fmap_5[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O29_N0_S1),.chainout(chainout_0_O29));
logic signed [63:0] chainout_2_O29; 
logic signed [63:0] O29_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O29(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_6[7:0]),.ay(-9'sd1),.bx(input_fmap_9[7:0]),.by( 9'sd1),.cx(input_fmap_10[7:0]),.cy( 9'sd1),.dx(input_fmap_11[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O29_N2_S1),.chainout(chainout_2_O29));
logic signed [63:0] chainout_4_O29; 
logic signed [63:0] O29_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O29(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_12[7:0]),.ay(-9'sd1),.bx(input_fmap_13[7:0]),.by( 9'sd1),.cx(input_fmap_16[7:0]),.cy( 9'sd1),.dx(input_fmap_19[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O29_N4_S1),.chainout(chainout_4_O29));
logic signed [63:0] chainout_6_O29; 
logic signed [63:0] O29_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O29(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_27[7:0]),.ay( 9'sd1),.bx(input_fmap_28[7:0]),.by( 9'sd1),.cx(input_fmap_32[7:0]),.cy( 9'sd1),.dx(input_fmap_34[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O29_N6_S1),.chainout(chainout_6_O29));
logic signed [63:0] chainout_8_O29; 
logic signed [63:0] O29_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O29(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_35[7:0]),.ay( 9'sd1),.bx(input_fmap_37[7:0]),.by(-9'sd1),.cx(input_fmap_39[7:0]),.cy( 9'sd1),.dx(input_fmap_42[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O29_N8_S1),.chainout(chainout_8_O29));
logic signed [63:0] chainout_10_O29; 
logic signed [63:0] O29_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O29(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_43[7:0]),.ay(-9'sd1),.bx(input_fmap_44[7:0]),.by( 9'sd1),.cx(input_fmap_45[7:0]),.cy(-9'sd1),.dx(input_fmap_46[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O29_N10_S1),.chainout(chainout_10_O29));
logic signed [63:0] chainout_12_O29; 
logic signed [63:0] O29_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O29(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_47[7:0]),.ay(-9'sd1),.bx(input_fmap_48[7:0]),.by( 9'sd1),.cx(input_fmap_51[7:0]),.cy( 9'sd2),.dx(input_fmap_52[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O29_N12_S1),.chainout(chainout_12_O29));
logic signed [63:0] chainout_14_O29; 
logic signed [63:0] O29_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O29(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_56[7:0]),.ay(-9'sd1),.bx(input_fmap_58[7:0]),.by(-9'sd2),.cx(input_fmap_59[7:0]),.cy(-9'sd1),.dx(input_fmap_61[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O29_N14_S1),.chainout(chainout_14_O29));
logic signed [63:0] chainout_16_O29; 
logic signed [63:0] O29_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O29(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_62[7:0]),.ay(-9'sd1),.bx(input_fmap_63[7:0]),.by( 9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O29_N16_S1),.chainout(chainout_16_O29));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O29_N0_S2;		always @(posedge clk) O29_N0_S2 <=     O29_N0_S1  +  O29_N2_S1 ;
 logic signed [21:0] O29_N2_S2;		always @(posedge clk) O29_N2_S2 <=     O29_N4_S1  +  O29_N6_S1 ;
 logic signed [21:0] O29_N4_S2;		always @(posedge clk) O29_N4_S2 <=     O29_N8_S1  +  O29_N10_S1 ;
 logic signed [21:0] O29_N6_S2;		always @(posedge clk) O29_N6_S2 <=     O29_N12_S1  +  O29_N14_S1 ;
 logic signed [21:0] O29_N8_S2;		always @(posedge clk) O29_N8_S2 <=     O29_N16_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O29_N0_S3;		always @(posedge clk) O29_N0_S3 <=     O29_N0_S2  +  O29_N2_S2 ;
 logic signed [22:0] O29_N2_S3;		always @(posedge clk) O29_N2_S3 <=     O29_N4_S2  +  O29_N6_S2 ;
 logic signed [22:0] O29_N4_S3;		always @(posedge clk) O29_N4_S3 <=     O29_N8_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O29_N0_S4;		always @(posedge clk) O29_N0_S4 <=     O29_N0_S3  +  O29_N2_S3 ;
 logic signed [23:0] O29_N2_S4;		always @(posedge clk) O29_N2_S4 <=     O29_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O29_N0_S5;		always @(posedge clk) O29_N0_S5 <=     O29_N0_S4  +  O29_N2_S4 ;
 assign conv_mac_29 = O29_N0_S5;

logic signed [31:0] conv_mac_30;
logic signed [63:0] chainout_0_O30; 
logic signed [63:0] O30_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O30(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay( 9'sd1),.bx(input_fmap_2[7:0]),.by(-9'sd1),.cx(input_fmap_4[7:0]),.cy(-9'sd2),.dx(input_fmap_5[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O30_N0_S1),.chainout(chainout_0_O30));
logic signed [63:0] chainout_2_O30; 
logic signed [63:0] O30_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O30(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_6[7:0]),.ay(-9'sd1),.bx(input_fmap_7[7:0]),.by(-9'sd1),.cx(input_fmap_9[7:0]),.cy( 9'sd1),.dx(input_fmap_14[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O30_N2_S1),.chainout(chainout_2_O30));
logic signed [63:0] chainout_4_O30; 
logic signed [63:0] O30_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O30(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_15[7:0]),.ay(-9'sd1),.bx(input_fmap_16[7:0]),.by(-9'sd1),.cx(input_fmap_18[7:0]),.cy(-9'sd1),.dx(input_fmap_19[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O30_N4_S1),.chainout(chainout_4_O30));
logic signed [63:0] chainout_6_O30; 
logic signed [63:0] O30_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O30(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_20[7:0]),.ay(-9'sd2),.bx(input_fmap_21[7:0]),.by(-9'sd3),.cx(input_fmap_22[7:0]),.cy( 9'sd2),.dx(input_fmap_23[7:0]),.dy( 9'sd3),.chainin(63'd0),.result(O30_N6_S1),.chainout(chainout_6_O30));
logic signed [63:0] chainout_8_O30; 
logic signed [63:0] O30_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O30(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_25[7:0]),.ay(-9'sd1),.bx(input_fmap_27[7:0]),.by( 9'sd2),.cx(input_fmap_28[7:0]),.cy( 9'sd1),.dx(input_fmap_30[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O30_N8_S1),.chainout(chainout_8_O30));
logic signed [63:0] chainout_10_O30; 
logic signed [63:0] O30_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O30(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_31[7:0]),.ay(-9'sd1),.bx(input_fmap_32[7:0]),.by(-9'sd1),.cx(input_fmap_34[7:0]),.cy( 9'sd3),.dx(input_fmap_37[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O30_N10_S1),.chainout(chainout_10_O30));
logic signed [63:0] chainout_12_O30; 
logic signed [63:0] O30_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O30(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_38[7:0]),.ay( 9'sd2),.bx(input_fmap_39[7:0]),.by( 9'sd1),.cx(input_fmap_40[7:0]),.cy( 9'sd2),.dx(input_fmap_41[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O30_N12_S1),.chainout(chainout_12_O30));
logic signed [63:0] chainout_14_O30; 
logic signed [63:0] O30_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O30(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_42[7:0]),.ay(-9'sd2),.bx(input_fmap_45[7:0]),.by( 9'sd1),.cx(input_fmap_46[7:0]),.cy( 9'sd2),.dx(input_fmap_48[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O30_N14_S1),.chainout(chainout_14_O30));
logic signed [63:0] chainout_16_O30; 
logic signed [63:0] O30_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O30(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_49[7:0]),.ay( 9'sd1),.bx(input_fmap_50[7:0]),.by(-9'sd2),.cx(input_fmap_52[7:0]),.cy( 9'sd2),.dx(input_fmap_53[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O30_N16_S1),.chainout(chainout_16_O30));
logic signed [63:0] chainout_18_O30; 
logic signed [63:0] O30_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O30(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_55[7:0]),.ay( 9'sd2),.bx(input_fmap_56[7:0]),.by(-9'sd4),.cx(input_fmap_57[7:0]),.cy( 9'sd2),.dx(input_fmap_59[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O30_N18_S1),.chainout(chainout_18_O30));
logic signed [63:0] chainout_20_O30; 
logic signed [63:0] O30_N20_S1; 
 int_sop_4_wrapper int_sop_4_inst_20_O30(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_61[7:0]),.ay(-9'sd3),.bx(input_fmap_63[7:0]),.by( 9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O30_N20_S1),.chainout(chainout_20_O30));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O30_N0_S2;		always @(posedge clk) O30_N0_S2 <=     O30_N0_S1  +  O30_N2_S1 ;
 logic signed [21:0] O30_N2_S2;		always @(posedge clk) O30_N2_S2 <=     O30_N4_S1  +  O30_N6_S1 ;
 logic signed [21:0] O30_N4_S2;		always @(posedge clk) O30_N4_S2 <=     O30_N8_S1  +  O30_N10_S1 ;
 logic signed [21:0] O30_N6_S2;		always @(posedge clk) O30_N6_S2 <=     O30_N12_S1  +  O30_N14_S1 ;
 logic signed [21:0] O30_N8_S2;		always @(posedge clk) O30_N8_S2 <=     O30_N16_S1  +  O30_N18_S1 ;
 logic signed [21:0] O30_N10_S2;		always @(posedge clk) O30_N10_S2 <=     O30_N20_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O30_N0_S3;		always @(posedge clk) O30_N0_S3 <=     O30_N0_S2  +  O30_N2_S2 ;
 logic signed [22:0] O30_N2_S3;		always @(posedge clk) O30_N2_S3 <=     O30_N4_S2  +  O30_N6_S2 ;
 logic signed [22:0] O30_N4_S3;		always @(posedge clk) O30_N4_S3 <=     O30_N8_S2  +  O30_N10_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O30_N0_S4;		always @(posedge clk) O30_N0_S4 <=     O30_N0_S3  +  O30_N2_S3 ;
 logic signed [23:0] O30_N2_S4;		always @(posedge clk) O30_N2_S4 <=     O30_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O30_N0_S5;		always @(posedge clk) O30_N0_S5 <=     O30_N0_S4  +  O30_N2_S4 ;
 assign conv_mac_30 = O30_N0_S5;

logic signed [31:0] conv_mac_31;
logic signed [63:0] chainout_0_O31; 
logic signed [63:0] O31_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O31(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay(-9'sd1),.bx(input_fmap_3[7:0]),.by( 9'sd2),.cx(input_fmap_4[7:0]),.cy(-9'sd1),.dx(input_fmap_5[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O31_N0_S1),.chainout(chainout_0_O31));
logic signed [63:0] chainout_2_O31; 
logic signed [63:0] O31_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O31(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_6[7:0]),.ay(-9'sd1),.bx(input_fmap_9[7:0]),.by( 9'sd1),.cx(input_fmap_10[7:0]),.cy( 9'sd1),.dx(input_fmap_11[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O31_N2_S1),.chainout(chainout_2_O31));
logic signed [63:0] chainout_4_O31; 
logic signed [63:0] O31_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O31(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_13[7:0]),.ay( 9'sd1),.bx(input_fmap_14[7:0]),.by( 9'sd1),.cx(input_fmap_15[7:0]),.cy( 9'sd1),.dx(input_fmap_16[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O31_N4_S1),.chainout(chainout_4_O31));
logic signed [63:0] chainout_6_O31; 
logic signed [63:0] O31_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O31(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_19[7:0]),.ay(-9'sd1),.bx(input_fmap_21[7:0]),.by(-9'sd1),.cx(input_fmap_22[7:0]),.cy(-9'sd1),.dx(input_fmap_27[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O31_N6_S1),.chainout(chainout_6_O31));
logic signed [63:0] chainout_8_O31; 
logic signed [63:0] O31_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O31(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_29[7:0]),.ay( 9'sd1),.bx(input_fmap_31[7:0]),.by(-9'sd1),.cx(input_fmap_34[7:0]),.cy( 9'sd1),.dx(input_fmap_35[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O31_N8_S1),.chainout(chainout_8_O31));
logic signed [63:0] chainout_10_O31; 
logic signed [63:0] O31_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O31(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_36[7:0]),.ay( 9'sd1),.bx(input_fmap_37[7:0]),.by( 9'sd1),.cx(input_fmap_38[7:0]),.cy( 9'sd1),.dx(input_fmap_40[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O31_N10_S1),.chainout(chainout_10_O31));
logic signed [63:0] chainout_12_O31; 
logic signed [63:0] O31_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O31(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_41[7:0]),.ay(-9'sd1),.bx(input_fmap_42[7:0]),.by( 9'sd1),.cx(input_fmap_43[7:0]),.cy( 9'sd2),.dx(input_fmap_45[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O31_N12_S1),.chainout(chainout_12_O31));
logic signed [63:0] chainout_14_O31; 
logic signed [63:0] O31_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O31(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_46[7:0]),.ay( 9'sd1),.bx(input_fmap_48[7:0]),.by( 9'sd1),.cx(input_fmap_51[7:0]),.cy(-9'sd2),.dx(input_fmap_52[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O31_N14_S1),.chainout(chainout_14_O31));
logic signed [63:0] chainout_16_O31; 
logic signed [63:0] O31_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O31(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_53[7:0]),.ay(-9'sd1),.bx(input_fmap_55[7:0]),.by( 9'sd1),.cx(input_fmap_56[7:0]),.cy( 9'sd1),.dx(input_fmap_58[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O31_N16_S1),.chainout(chainout_16_O31));
logic signed [63:0] chainout_18_O31; 
logic signed [63:0] O31_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O31(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_60[7:0]),.ay( 9'sd1),.bx(input_fmap_61[7:0]),.by(-9'sd1),.cx(input_fmap_63[7:0]),.cy( 9'sd1),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O31_N18_S1),.chainout(chainout_18_O31));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O31_N0_S2;		always @(posedge clk) O31_N0_S2 <=     O31_N0_S1  +  O31_N2_S1 ;
 logic signed [21:0] O31_N2_S2;		always @(posedge clk) O31_N2_S2 <=     O31_N4_S1  +  O31_N6_S1 ;
 logic signed [21:0] O31_N4_S2;		always @(posedge clk) O31_N4_S2 <=     O31_N8_S1  +  O31_N10_S1 ;
 logic signed [21:0] O31_N6_S2;		always @(posedge clk) O31_N6_S2 <=     O31_N12_S1  +  O31_N14_S1 ;
 logic signed [21:0] O31_N8_S2;		always @(posedge clk) O31_N8_S2 <=     O31_N16_S1  +  O31_N18_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O31_N0_S3;		always @(posedge clk) O31_N0_S3 <=     O31_N0_S2  +  O31_N2_S2 ;
 logic signed [22:0] O31_N2_S3;		always @(posedge clk) O31_N2_S3 <=     O31_N4_S2  +  O31_N6_S2 ;
 logic signed [22:0] O31_N4_S3;		always @(posedge clk) O31_N4_S3 <=     O31_N8_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O31_N0_S4;		always @(posedge clk) O31_N0_S4 <=     O31_N0_S3  +  O31_N2_S3 ;
 logic signed [23:0] O31_N2_S4;		always @(posedge clk) O31_N2_S4 <=     O31_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O31_N0_S5;		always @(posedge clk) O31_N0_S5 <=     O31_N0_S4  +  O31_N2_S4 ;
 assign conv_mac_31 = O31_N0_S5;

logic signed [31:0] conv_mac_32;
logic signed [63:0] chainout_0_O32; 
logic signed [63:0] O32_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O32(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_2[7:0]),.ay( 9'sd1),.bx(input_fmap_13[7:0]),.by(-9'sd1),.cx(input_fmap_16[7:0]),.cy(-9'sd1),.dx(input_fmap_20[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O32_N0_S1),.chainout(chainout_0_O32));
logic signed [63:0] chainout_2_O32; 
logic signed [63:0] O32_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O32(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_24[7:0]),.ay( 9'sd7),.bx(input_fmap_30[7:0]),.by(-9'sd1),.cx(input_fmap_50[7:0]),.cy(-9'sd1),.dx(input_fmap_63[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O32_N2_S1),.chainout(chainout_2_O32));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O32_N0_S2;		always @(posedge clk) O32_N0_S2 <=     O32_N0_S1  +  O32_N2_S1 ;
 assign conv_mac_32 = O32_N0_S2;

logic signed [31:0] conv_mac_33;
logic signed [63:0] chainout_0_O33; 
logic signed [63:0] O33_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O33(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_2[7:0]),.ay(-9'sd1),.bx(input_fmap_6[7:0]),.by( 9'sd1),.cx(input_fmap_7[7:0]),.cy( 9'sd1),.dx(input_fmap_8[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O33_N0_S1),.chainout(chainout_0_O33));
logic signed [63:0] chainout_2_O33; 
logic signed [63:0] O33_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O33(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_10[7:0]),.ay(-9'sd1),.bx(input_fmap_11[7:0]),.by(-9'sd1),.cx(input_fmap_12[7:0]),.cy( 9'sd2),.dx(input_fmap_13[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O33_N2_S1),.chainout(chainout_2_O33));
logic signed [63:0] chainout_4_O33; 
logic signed [63:0] O33_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O33(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_16[7:0]),.ay(-9'sd1),.bx(input_fmap_18[7:0]),.by(-9'sd1),.cx(input_fmap_20[7:0]),.cy(-9'sd1),.dx(input_fmap_23[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O33_N4_S1),.chainout(chainout_4_O33));
logic signed [63:0] chainout_6_O33; 
logic signed [63:0] O33_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O33(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_26[7:0]),.ay( 9'sd2),.bx(input_fmap_32[7:0]),.by(-9'sd1),.cx(input_fmap_33[7:0]),.cy(-9'sd1),.dx(input_fmap_34[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O33_N6_S1),.chainout(chainout_6_O33));
logic signed [63:0] chainout_8_O33; 
logic signed [63:0] O33_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O33(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_35[7:0]),.ay(-9'sd1),.bx(input_fmap_37[7:0]),.by(-9'sd1),.cx(input_fmap_38[7:0]),.cy(-9'sd1),.dx(input_fmap_40[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O33_N8_S1),.chainout(chainout_8_O33));
logic signed [63:0] chainout_10_O33; 
logic signed [63:0] O33_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O33(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_43[7:0]),.ay(-9'sd1),.bx(input_fmap_44[7:0]),.by(-9'sd1),.cx(input_fmap_45[7:0]),.cy( 9'sd1),.dx(input_fmap_46[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O33_N10_S1),.chainout(chainout_10_O33));
logic signed [63:0] chainout_12_O33; 
logic signed [63:0] O33_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O33(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_47[7:0]),.ay(-9'sd2),.bx(input_fmap_48[7:0]),.by( 9'sd1),.cx(input_fmap_49[7:0]),.cy(-9'sd1),.dx(input_fmap_51[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O33_N12_S1),.chainout(chainout_12_O33));
logic signed [63:0] chainout_14_O33; 
logic signed [63:0] O33_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O33(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_53[7:0]),.ay( 9'sd2),.bx(input_fmap_57[7:0]),.by(-9'sd1),.cx(input_fmap_59[7:0]),.cy( 9'sd1),.dx(input_fmap_60[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O33_N14_S1),.chainout(chainout_14_O33));
logic signed [63:0] chainout_16_O33; 
logic signed [63:0] O33_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O33(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_62[7:0]),.ay(-9'sd1),.bx(input_fmap_63[7:0]),.by( 9'sd3),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O33_N16_S1),.chainout(chainout_16_O33));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O33_N0_S2;		always @(posedge clk) O33_N0_S2 <=     O33_N0_S1  +  O33_N2_S1 ;
 logic signed [21:0] O33_N2_S2;		always @(posedge clk) O33_N2_S2 <=     O33_N4_S1  +  O33_N6_S1 ;
 logic signed [21:0] O33_N4_S2;		always @(posedge clk) O33_N4_S2 <=     O33_N8_S1  +  O33_N10_S1 ;
 logic signed [21:0] O33_N6_S2;		always @(posedge clk) O33_N6_S2 <=     O33_N12_S1  +  O33_N14_S1 ;
 logic signed [21:0] O33_N8_S2;		always @(posedge clk) O33_N8_S2 <=     O33_N16_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O33_N0_S3;		always @(posedge clk) O33_N0_S3 <=     O33_N0_S2  +  O33_N2_S2 ;
 logic signed [22:0] O33_N2_S3;		always @(posedge clk) O33_N2_S3 <=     O33_N4_S2  +  O33_N6_S2 ;
 logic signed [22:0] O33_N4_S3;		always @(posedge clk) O33_N4_S3 <=     O33_N8_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O33_N0_S4;		always @(posedge clk) O33_N0_S4 <=     O33_N0_S3  +  O33_N2_S3 ;
 logic signed [23:0] O33_N2_S4;		always @(posedge clk) O33_N2_S4 <=     O33_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O33_N0_S5;		always @(posedge clk) O33_N0_S5 <=     O33_N0_S4  +  O33_N2_S4 ;
 assign conv_mac_33 = O33_N0_S5;

logic signed [31:0] conv_mac_34;
logic signed [63:0] chainout_0_O34; 
logic signed [63:0] O34_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O34(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd1),.bx(input_fmap_1[7:0]),.by(-9'sd1),.cx(input_fmap_2[7:0]),.cy(-9'sd2),.dx(input_fmap_3[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O34_N0_S1),.chainout(chainout_0_O34));
logic signed [63:0] chainout_2_O34; 
logic signed [63:0] O34_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O34(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_7[7:0]),.ay( 9'sd1),.bx(input_fmap_8[7:0]),.by(-9'sd2),.cx(input_fmap_10[7:0]),.cy( 9'sd2),.dx(input_fmap_12[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O34_N2_S1),.chainout(chainout_2_O34));
logic signed [63:0] chainout_4_O34; 
logic signed [63:0] O34_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O34(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_18[7:0]),.ay( 9'sd2),.bx(input_fmap_19[7:0]),.by(-9'sd1),.cx(input_fmap_21[7:0]),.cy( 9'sd3),.dx(input_fmap_22[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O34_N4_S1),.chainout(chainout_4_O34));
logic signed [63:0] chainout_6_O34; 
logic signed [63:0] O34_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O34(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_23[7:0]),.ay( 9'sd1),.bx(input_fmap_26[7:0]),.by(-9'sd2),.cx(input_fmap_27[7:0]),.cy(-9'sd1),.dx(input_fmap_28[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O34_N6_S1),.chainout(chainout_6_O34));
logic signed [63:0] chainout_8_O34; 
logic signed [63:0] O34_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O34(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_29[7:0]),.ay(-9'sd1),.bx(input_fmap_30[7:0]),.by(-9'sd2),.cx(input_fmap_33[7:0]),.cy(-9'sd1),.dx(input_fmap_35[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O34_N8_S1),.chainout(chainout_8_O34));
logic signed [63:0] chainout_10_O34; 
logic signed [63:0] O34_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O34(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_38[7:0]),.ay(-9'sd2),.bx(input_fmap_40[7:0]),.by(-9'sd1),.cx(input_fmap_43[7:0]),.cy(-9'sd1),.dx(input_fmap_44[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O34_N10_S1),.chainout(chainout_10_O34));
logic signed [63:0] chainout_12_O34; 
logic signed [63:0] O34_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O34(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_46[7:0]),.ay( 9'sd4),.bx(input_fmap_49[7:0]),.by(-9'sd1),.cx(input_fmap_50[7:0]),.cy(-9'sd1),.dx(input_fmap_55[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O34_N12_S1),.chainout(chainout_12_O34));
logic signed [63:0] chainout_14_O34; 
logic signed [63:0] O34_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O34(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_56[7:0]),.ay(-9'sd2),.bx(input_fmap_57[7:0]),.by(-9'sd1),.cx(input_fmap_59[7:0]),.cy(-9'sd1),.dx(input_fmap_60[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O34_N14_S1),.chainout(chainout_14_O34));
logic signed [63:0] chainout_16_O34; 
logic signed [63:0] O34_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O34(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_62[7:0]),.ay( 9'sd1),.bx(input_fmap_63[7:0]),.by(-9'sd3),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O34_N16_S1),.chainout(chainout_16_O34));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O34_N0_S2;		always @(posedge clk) O34_N0_S2 <=     O34_N0_S1  +  O34_N2_S1 ;
 logic signed [21:0] O34_N2_S2;		always @(posedge clk) O34_N2_S2 <=     O34_N4_S1  +  O34_N6_S1 ;
 logic signed [21:0] O34_N4_S2;		always @(posedge clk) O34_N4_S2 <=     O34_N8_S1  +  O34_N10_S1 ;
 logic signed [21:0] O34_N6_S2;		always @(posedge clk) O34_N6_S2 <=     O34_N12_S1  +  O34_N14_S1 ;
 logic signed [21:0] O34_N8_S2;		always @(posedge clk) O34_N8_S2 <=     O34_N16_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O34_N0_S3;		always @(posedge clk) O34_N0_S3 <=     O34_N0_S2  +  O34_N2_S2 ;
 logic signed [22:0] O34_N2_S3;		always @(posedge clk) O34_N2_S3 <=     O34_N4_S2  +  O34_N6_S2 ;
 logic signed [22:0] O34_N4_S3;		always @(posedge clk) O34_N4_S3 <=     O34_N8_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O34_N0_S4;		always @(posedge clk) O34_N0_S4 <=     O34_N0_S3  +  O34_N2_S3 ;
 logic signed [23:0] O34_N2_S4;		always @(posedge clk) O34_N2_S4 <=     O34_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O34_N0_S5;		always @(posedge clk) O34_N0_S5 <=     O34_N0_S4  +  O34_N2_S4 ;
 assign conv_mac_34 = O34_N0_S5;

logic signed [31:0] conv_mac_35;
logic signed [63:0] chainout_0_O35; 
logic signed [63:0] O35_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O35(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_4[7:0]),.ay(-9'sd1),.bx(input_fmap_6[7:0]),.by( 9'sd1),.cx(input_fmap_9[7:0]),.cy( 9'sd1),.dx(input_fmap_10[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O35_N0_S1),.chainout(chainout_0_O35));
logic signed [63:0] chainout_2_O35; 
logic signed [63:0] O35_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O35(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_15[7:0]),.ay(-9'sd1),.bx(input_fmap_17[7:0]),.by(-9'sd1),.cx(input_fmap_19[7:0]),.cy( 9'sd1),.dx(input_fmap_22[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O35_N2_S1),.chainout(chainout_2_O35));
logic signed [63:0] chainout_4_O35; 
logic signed [63:0] O35_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O35(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_27[7:0]),.ay(-9'sd1),.bx(input_fmap_28[7:0]),.by( 9'sd2),.cx(input_fmap_29[7:0]),.cy( 9'sd1),.dx(input_fmap_30[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O35_N4_S1),.chainout(chainout_4_O35));
logic signed [63:0] chainout_6_O35; 
logic signed [63:0] O35_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O35(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_31[7:0]),.ay( 9'sd1),.bx(input_fmap_32[7:0]),.by(-9'sd1),.cx(input_fmap_34[7:0]),.cy( 9'sd2),.dx(input_fmap_35[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O35_N6_S1),.chainout(chainout_6_O35));
logic signed [63:0] chainout_8_O35; 
logic signed [63:0] O35_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O35(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_36[7:0]),.ay( 9'sd1),.bx(input_fmap_42[7:0]),.by(-9'sd1),.cx(input_fmap_43[7:0]),.cy(-9'sd1),.dx(input_fmap_46[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O35_N8_S1),.chainout(chainout_8_O35));
logic signed [63:0] chainout_10_O35; 
logic signed [63:0] O35_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O35(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_48[7:0]),.ay( 9'sd1),.bx(input_fmap_49[7:0]),.by( 9'sd1),.cx(input_fmap_50[7:0]),.cy( 9'sd1),.dx(input_fmap_56[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O35_N10_S1),.chainout(chainout_10_O35));
logic signed [63:0] chainout_12_O35; 
logic signed [63:0] O35_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O35(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_58[7:0]),.ay( 9'sd1),.bx(input_fmap_62[7:0]),.by( 9'sd1),.cx(input_fmap_63[7:0]),.cy( 9'sd1),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O35_N12_S1),.chainout(chainout_12_O35));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O35_N0_S2;		always @(posedge clk) O35_N0_S2 <=     O35_N0_S1  +  O35_N2_S1 ;
 logic signed [21:0] O35_N2_S2;		always @(posedge clk) O35_N2_S2 <=     O35_N4_S1  +  O35_N6_S1 ;
 logic signed [21:0] O35_N4_S2;		always @(posedge clk) O35_N4_S2 <=     O35_N8_S1  +  O35_N10_S1 ;
 logic signed [21:0] O35_N6_S2;		always @(posedge clk) O35_N6_S2 <=     O35_N12_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O35_N0_S3;		always @(posedge clk) O35_N0_S3 <=     O35_N0_S2  +  O35_N2_S2 ;
 logic signed [22:0] O35_N2_S3;		always @(posedge clk) O35_N2_S3 <=     O35_N4_S2  +  O35_N6_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O35_N0_S4;		always @(posedge clk) O35_N0_S4 <=     O35_N0_S3  +  O35_N2_S3 ;
 assign conv_mac_35 = O35_N0_S4;

logic signed [31:0] conv_mac_36;
logic signed [63:0] chainout_0_O36; 
logic signed [63:0] O36_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O36(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd1),.bx(input_fmap_2[7:0]),.by(-9'sd1),.cx(input_fmap_6[7:0]),.cy(-9'sd1),.dx(input_fmap_7[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O36_N0_S1),.chainout(chainout_0_O36));
logic signed [63:0] chainout_2_O36; 
logic signed [63:0] O36_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O36(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_8[7:0]),.ay( 9'sd1),.bx(input_fmap_10[7:0]),.by(-9'sd1),.cx(input_fmap_14[7:0]),.cy(-9'sd2),.dx(input_fmap_15[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O36_N2_S1),.chainout(chainout_2_O36));
logic signed [63:0] chainout_4_O36; 
logic signed [63:0] O36_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O36(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_17[7:0]),.ay(-9'sd2),.bx(input_fmap_18[7:0]),.by(-9'sd1),.cx(input_fmap_20[7:0]),.cy(-9'sd1),.dx(input_fmap_22[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O36_N4_S1),.chainout(chainout_4_O36));
logic signed [63:0] chainout_6_O36; 
logic signed [63:0] O36_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O36(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_24[7:0]),.ay( 9'sd5),.bx(input_fmap_25[7:0]),.by(-9'sd1),.cx(input_fmap_27[7:0]),.cy( 9'sd1),.dx(input_fmap_28[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O36_N6_S1),.chainout(chainout_6_O36));
logic signed [63:0] chainout_8_O36; 
logic signed [63:0] O36_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O36(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_30[7:0]),.ay( 9'sd2),.bx(input_fmap_35[7:0]),.by( 9'sd2),.cx(input_fmap_36[7:0]),.cy( 9'sd1),.dx(input_fmap_37[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O36_N8_S1),.chainout(chainout_8_O36));
logic signed [63:0] chainout_10_O36; 
logic signed [63:0] O36_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O36(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_38[7:0]),.ay( 9'sd4),.bx(input_fmap_39[7:0]),.by(-9'sd1),.cx(input_fmap_41[7:0]),.cy(-9'sd2),.dx(input_fmap_45[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O36_N10_S1),.chainout(chainout_10_O36));
logic signed [63:0] chainout_12_O36; 
logic signed [63:0] O36_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O36(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_46[7:0]),.ay( 9'sd1),.bx(input_fmap_47[7:0]),.by(-9'sd1),.cx(input_fmap_48[7:0]),.cy( 9'sd1),.dx(input_fmap_50[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O36_N12_S1),.chainout(chainout_12_O36));
logic signed [63:0] chainout_14_O36; 
logic signed [63:0] O36_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O36(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_51[7:0]),.ay( 9'sd2),.bx(input_fmap_55[7:0]),.by(-9'sd3),.cx(input_fmap_56[7:0]),.cy( 9'sd2),.dx(input_fmap_58[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O36_N14_S1),.chainout(chainout_14_O36));
logic signed [63:0] chainout_16_O36; 
logic signed [63:0] O36_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O36(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_59[7:0]),.ay( 9'sd1),.bx(input_fmap_60[7:0]),.by( 9'sd1),.cx(input_fmap_61[7:0]),.cy(-9'sd1),.dx(input_fmap_62[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O36_N16_S1),.chainout(chainout_16_O36));
logic signed [63:0] chainout_18_O36; 
logic signed [63:0] O36_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O36(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_63[7:0]),.ay( 9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O36_N18_S1),.chainout(chainout_18_O36));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O36_N0_S2;		always @(posedge clk) O36_N0_S2 <=     O36_N0_S1  +  O36_N2_S1 ;
 logic signed [21:0] O36_N2_S2;		always @(posedge clk) O36_N2_S2 <=     O36_N4_S1  +  O36_N6_S1 ;
 logic signed [21:0] O36_N4_S2;		always @(posedge clk) O36_N4_S2 <=     O36_N8_S1  +  O36_N10_S1 ;
 logic signed [21:0] O36_N6_S2;		always @(posedge clk) O36_N6_S2 <=     O36_N12_S1  +  O36_N14_S1 ;
 logic signed [21:0] O36_N8_S2;		always @(posedge clk) O36_N8_S2 <=     O36_N16_S1  +  O36_N18_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O36_N0_S3;		always @(posedge clk) O36_N0_S3 <=     O36_N0_S2  +  O36_N2_S2 ;
 logic signed [22:0] O36_N2_S3;		always @(posedge clk) O36_N2_S3 <=     O36_N4_S2  +  O36_N6_S2 ;
 logic signed [22:0] O36_N4_S3;		always @(posedge clk) O36_N4_S3 <=     O36_N8_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O36_N0_S4;		always @(posedge clk) O36_N0_S4 <=     O36_N0_S3  +  O36_N2_S3 ;
 logic signed [23:0] O36_N2_S4;		always @(posedge clk) O36_N2_S4 <=     O36_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O36_N0_S5;		always @(posedge clk) O36_N0_S5 <=     O36_N0_S4  +  O36_N2_S4 ;
 assign conv_mac_36 = O36_N0_S5;

logic signed [31:0] conv_mac_37;
logic signed [63:0] chainout_0_O37; 
logic signed [63:0] O37_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O37(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd1),.bx(input_fmap_2[7:0]),.by( 9'sd1),.cx(input_fmap_3[7:0]),.cy( 9'sd1),.dx(input_fmap_4[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O37_N0_S1),.chainout(chainout_0_O37));
logic signed [63:0] chainout_2_O37; 
logic signed [63:0] O37_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O37(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_8[7:0]),.ay( 9'sd1),.bx(input_fmap_11[7:0]),.by( 9'sd1),.cx(input_fmap_14[7:0]),.cy( 9'sd1),.dx(input_fmap_15[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O37_N2_S1),.chainout(chainout_2_O37));
logic signed [63:0] chainout_4_O37; 
logic signed [63:0] O37_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O37(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_17[7:0]),.ay( 9'sd1),.bx(input_fmap_18[7:0]),.by(-9'sd2),.cx(input_fmap_19[7:0]),.cy(-9'sd1),.dx(input_fmap_20[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O37_N4_S1),.chainout(chainout_4_O37));
logic signed [63:0] chainout_6_O37; 
logic signed [63:0] O37_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O37(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_23[7:0]),.ay(-9'sd1),.bx(input_fmap_24[7:0]),.by(-9'sd1),.cx(input_fmap_25[7:0]),.cy( 9'sd1),.dx(input_fmap_26[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O37_N6_S1),.chainout(chainout_6_O37));
logic signed [63:0] chainout_8_O37; 
logic signed [63:0] O37_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O37(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_28[7:0]),.ay( 9'sd1),.bx(input_fmap_30[7:0]),.by( 9'sd2),.cx(input_fmap_32[7:0]),.cy( 9'sd1),.dx(input_fmap_35[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O37_N8_S1),.chainout(chainout_8_O37));
logic signed [63:0] chainout_10_O37; 
logic signed [63:0] O37_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O37(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_38[7:0]),.ay(-9'sd1),.bx(input_fmap_43[7:0]),.by(-9'sd1),.cx(input_fmap_45[7:0]),.cy(-9'sd1),.dx(input_fmap_46[7:0]),.dy(-9'sd3),.chainin(63'd0),.result(O37_N10_S1),.chainout(chainout_10_O37));
logic signed [63:0] chainout_12_O37; 
logic signed [63:0] O37_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O37(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_47[7:0]),.ay( 9'sd3),.bx(input_fmap_48[7:0]),.by( 9'sd1),.cx(input_fmap_50[7:0]),.cy(-9'sd2),.dx(input_fmap_52[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O37_N12_S1),.chainout(chainout_12_O37));
logic signed [63:0] chainout_14_O37; 
logic signed [63:0] O37_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O37(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_53[7:0]),.ay( 9'sd1),.bx(input_fmap_54[7:0]),.by(-9'sd1),.cx(input_fmap_56[7:0]),.cy(-9'sd1),.dx(input_fmap_57[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O37_N14_S1),.chainout(chainout_14_O37));
logic signed [63:0] chainout_16_O37; 
logic signed [63:0] O37_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O37(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_59[7:0]),.ay( 9'sd1),.bx(input_fmap_61[7:0]),.by(-9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O37_N16_S1),.chainout(chainout_16_O37));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O37_N0_S2;		always @(posedge clk) O37_N0_S2 <=     O37_N0_S1  +  O37_N2_S1 ;
 logic signed [21:0] O37_N2_S2;		always @(posedge clk) O37_N2_S2 <=     O37_N4_S1  +  O37_N6_S1 ;
 logic signed [21:0] O37_N4_S2;		always @(posedge clk) O37_N4_S2 <=     O37_N8_S1  +  O37_N10_S1 ;
 logic signed [21:0] O37_N6_S2;		always @(posedge clk) O37_N6_S2 <=     O37_N12_S1  +  O37_N14_S1 ;
 logic signed [21:0] O37_N8_S2;		always @(posedge clk) O37_N8_S2 <=     O37_N16_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O37_N0_S3;		always @(posedge clk) O37_N0_S3 <=     O37_N0_S2  +  O37_N2_S2 ;
 logic signed [22:0] O37_N2_S3;		always @(posedge clk) O37_N2_S3 <=     O37_N4_S2  +  O37_N6_S2 ;
 logic signed [22:0] O37_N4_S3;		always @(posedge clk) O37_N4_S3 <=     O37_N8_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O37_N0_S4;		always @(posedge clk) O37_N0_S4 <=     O37_N0_S3  +  O37_N2_S3 ;
 logic signed [23:0] O37_N2_S4;		always @(posedge clk) O37_N2_S4 <=     O37_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O37_N0_S5;		always @(posedge clk) O37_N0_S5 <=     O37_N0_S4  +  O37_N2_S4 ;
 assign conv_mac_37 = O37_N0_S5;

logic signed [31:0] conv_mac_38;
logic signed [63:0] chainout_0_O38; 
logic signed [63:0] O38_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O38(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_15[7:0]),.ay( 9'sd1),.bx(input_fmap_17[7:0]),.by(-9'sd1),.cx(input_fmap_20[7:0]),.cy(-9'sd1),.dx(input_fmap_25[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O38_N0_S1),.chainout(chainout_0_O38));
logic signed [63:0] chainout_2_O38; 
logic signed [63:0] O38_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O38(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_27[7:0]),.ay(-9'sd1),.bx(input_fmap_33[7:0]),.by(-9'sd1),.cx(input_fmap_34[7:0]),.cy(-9'sd1),.dx(input_fmap_36[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O38_N2_S1),.chainout(chainout_2_O38));
logic signed [63:0] chainout_4_O38; 
logic signed [63:0] O38_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O38(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_37[7:0]),.ay(-9'sd1),.bx(input_fmap_40[7:0]),.by(-9'sd1),.cx(input_fmap_46[7:0]),.cy(-9'sd1),.dx(input_fmap_50[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O38_N4_S1),.chainout(chainout_4_O38));
logic signed [63:0] chainout_6_O38; 
logic signed [63:0] O38_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O38(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_52[7:0]),.ay( 9'sd3),.bx(input_fmap_54[7:0]),.by( 9'sd1),.cx(input_fmap_55[7:0]),.cy( 9'sd1),.dx(input_fmap_57[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O38_N6_S1),.chainout(chainout_6_O38));
logic signed [63:0] chainout_8_O38; 
logic signed [63:0] O38_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O38(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_58[7:0]),.ay(-9'sd1),.bx(input_fmap_61[7:0]),.by( 9'sd1),.cx(input_fmap_62[7:0]),.cy( 9'sd1),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O38_N8_S1),.chainout(chainout_8_O38));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O38_N0_S2;		always @(posedge clk) O38_N0_S2 <=     O38_N0_S1  +  O38_N2_S1 ;
 logic signed [21:0] O38_N2_S2;		always @(posedge clk) O38_N2_S2 <=     O38_N4_S1  +  O38_N6_S1 ;
 logic signed [21:0] O38_N4_S2;		always @(posedge clk) O38_N4_S2 <=     O38_N8_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O38_N0_S3;		always @(posedge clk) O38_N0_S3 <=     O38_N0_S2  +  O38_N2_S2 ;
 logic signed [22:0] O38_N2_S3;		always @(posedge clk) O38_N2_S3 <=     O38_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O38_N0_S4;		always @(posedge clk) O38_N0_S4 <=     O38_N0_S3  +  O38_N2_S3 ;
 assign conv_mac_38 = O38_N0_S4;

logic signed [31:0] conv_mac_39;
logic signed [63:0] chainout_0_O39; 
logic signed [63:0] O39_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O39(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd1),.bx(input_fmap_2[7:0]),.by( 9'sd1),.cx(input_fmap_3[7:0]),.cy(-9'sd1),.dx(input_fmap_5[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O39_N0_S1),.chainout(chainout_0_O39));
logic signed [63:0] chainout_2_O39; 
logic signed [63:0] O39_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O39(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_7[7:0]),.ay(-9'sd2),.bx(input_fmap_8[7:0]),.by( 9'sd1),.cx(input_fmap_10[7:0]),.cy(-9'sd1),.dx(input_fmap_11[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O39_N2_S1),.chainout(chainout_2_O39));
logic signed [63:0] chainout_4_O39; 
logic signed [63:0] O39_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O39(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_12[7:0]),.ay(-9'sd1),.bx(input_fmap_14[7:0]),.by( 9'sd1),.cx(input_fmap_15[7:0]),.cy(-9'sd1),.dx(input_fmap_17[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O39_N4_S1),.chainout(chainout_4_O39));
logic signed [63:0] chainout_6_O39; 
logic signed [63:0] O39_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O39(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_18[7:0]),.ay(-9'sd1),.bx(input_fmap_19[7:0]),.by(-9'sd1),.cx(input_fmap_20[7:0]),.cy( 9'sd1),.dx(input_fmap_23[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O39_N6_S1),.chainout(chainout_6_O39));
logic signed [63:0] chainout_8_O39; 
logic signed [63:0] O39_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O39(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_24[7:0]),.ay(-9'sd1),.bx(input_fmap_25[7:0]),.by( 9'sd2),.cx(input_fmap_26[7:0]),.cy( 9'sd1),.dx(input_fmap_27[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O39_N8_S1),.chainout(chainout_8_O39));
logic signed [63:0] chainout_10_O39; 
logic signed [63:0] O39_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O39(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_28[7:0]),.ay(-9'sd1),.bx(input_fmap_29[7:0]),.by( 9'sd2),.cx(input_fmap_30[7:0]),.cy( 9'sd2),.dx(input_fmap_31[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O39_N10_S1),.chainout(chainout_10_O39));
logic signed [63:0] chainout_12_O39; 
logic signed [63:0] O39_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O39(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_36[7:0]),.ay( 9'sd1),.bx(input_fmap_37[7:0]),.by( 9'sd1),.cx(input_fmap_38[7:0]),.cy( 9'sd1),.dx(input_fmap_39[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O39_N12_S1),.chainout(chainout_12_O39));
logic signed [63:0] chainout_14_O39; 
logic signed [63:0] O39_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O39(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_44[7:0]),.ay( 9'sd1),.bx(input_fmap_45[7:0]),.by( 9'sd1),.cx(input_fmap_48[7:0]),.cy( 9'sd1),.dx(input_fmap_49[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O39_N14_S1),.chainout(chainout_14_O39));
logic signed [63:0] chainout_16_O39; 
logic signed [63:0] O39_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O39(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_51[7:0]),.ay(-9'sd2),.bx(input_fmap_52[7:0]),.by( 9'sd1),.cx(input_fmap_55[7:0]),.cy(-9'sd1),.dx(input_fmap_58[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O39_N16_S1),.chainout(chainout_16_O39));
logic signed [63:0] chainout_18_O39; 
logic signed [63:0] O39_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O39(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_59[7:0]),.ay( 9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O39_N18_S1),.chainout(chainout_18_O39));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O39_N0_S2;		always @(posedge clk) O39_N0_S2 <=     O39_N0_S1  +  O39_N2_S1 ;
 logic signed [21:0] O39_N2_S2;		always @(posedge clk) O39_N2_S2 <=     O39_N4_S1  +  O39_N6_S1 ;
 logic signed [21:0] O39_N4_S2;		always @(posedge clk) O39_N4_S2 <=     O39_N8_S1  +  O39_N10_S1 ;
 logic signed [21:0] O39_N6_S2;		always @(posedge clk) O39_N6_S2 <=     O39_N12_S1  +  O39_N14_S1 ;
 logic signed [21:0] O39_N8_S2;		always @(posedge clk) O39_N8_S2 <=     O39_N16_S1  +  O39_N18_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O39_N0_S3;		always @(posedge clk) O39_N0_S3 <=     O39_N0_S2  +  O39_N2_S2 ;
 logic signed [22:0] O39_N2_S3;		always @(posedge clk) O39_N2_S3 <=     O39_N4_S2  +  O39_N6_S2 ;
 logic signed [22:0] O39_N4_S3;		always @(posedge clk) O39_N4_S3 <=     O39_N8_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O39_N0_S4;		always @(posedge clk) O39_N0_S4 <=     O39_N0_S3  +  O39_N2_S3 ;
 logic signed [23:0] O39_N2_S4;		always @(posedge clk) O39_N2_S4 <=     O39_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O39_N0_S5;		always @(posedge clk) O39_N0_S5 <=     O39_N0_S4  +  O39_N2_S4 ;
 assign conv_mac_39 = O39_N0_S5;

logic signed [31:0] conv_mac_40;
logic signed [63:0] chainout_0_O40; 
logic signed [63:0] O40_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O40(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay( 9'sd1),.bx(input_fmap_2[7:0]),.by( 9'sd1),.cx(input_fmap_3[7:0]),.cy(-9'sd1),.dx(input_fmap_4[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O40_N0_S1),.chainout(chainout_0_O40));
logic signed [63:0] chainout_2_O40; 
logic signed [63:0] O40_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O40(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_8[7:0]),.ay( 9'sd1),.bx(input_fmap_9[7:0]),.by(-9'sd1),.cx(input_fmap_13[7:0]),.cy( 9'sd1),.dx(input_fmap_14[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O40_N2_S1),.chainout(chainout_2_O40));
logic signed [63:0] chainout_4_O40; 
logic signed [63:0] O40_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O40(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_15[7:0]),.ay(-9'sd2),.bx(input_fmap_17[7:0]),.by( 9'sd1),.cx(input_fmap_20[7:0]),.cy( 9'sd1),.dx(input_fmap_26[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O40_N4_S1),.chainout(chainout_4_O40));
logic signed [63:0] chainout_6_O40; 
logic signed [63:0] O40_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O40(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_28[7:0]),.ay( 9'sd2),.bx(input_fmap_30[7:0]),.by(-9'sd2),.cx(input_fmap_31[7:0]),.cy( 9'sd1),.dx(input_fmap_32[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O40_N6_S1),.chainout(chainout_6_O40));
logic signed [63:0] chainout_8_O40; 
logic signed [63:0] O40_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O40(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_34[7:0]),.ay(-9'sd1),.bx(input_fmap_35[7:0]),.by(-9'sd1),.cx(input_fmap_36[7:0]),.cy(-9'sd1),.dx(input_fmap_39[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O40_N8_S1),.chainout(chainout_8_O40));
logic signed [63:0] chainout_10_O40; 
logic signed [63:0] O40_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O40(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_41[7:0]),.ay( 9'sd1),.bx(input_fmap_42[7:0]),.by(-9'sd1),.cx(input_fmap_43[7:0]),.cy( 9'sd1),.dx(input_fmap_46[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O40_N10_S1),.chainout(chainout_10_O40));
logic signed [63:0] chainout_12_O40; 
logic signed [63:0] O40_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O40(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_47[7:0]),.ay( 9'sd1),.bx(input_fmap_51[7:0]),.by(-9'sd1),.cx(input_fmap_52[7:0]),.cy(-9'sd1),.dx(input_fmap_53[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O40_N12_S1),.chainout(chainout_12_O40));
logic signed [63:0] chainout_14_O40; 
logic signed [63:0] O40_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O40(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_56[7:0]),.ay(-9'sd1),.bx(input_fmap_57[7:0]),.by(-9'sd2),.cx(input_fmap_60[7:0]),.cy(-9'sd1),.dx(input_fmap_61[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O40_N14_S1),.chainout(chainout_14_O40));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O40_N0_S2;		always @(posedge clk) O40_N0_S2 <=     O40_N0_S1  +  O40_N2_S1 ;
 logic signed [21:0] O40_N2_S2;		always @(posedge clk) O40_N2_S2 <=     O40_N4_S1  +  O40_N6_S1 ;
 logic signed [21:0] O40_N4_S2;		always @(posedge clk) O40_N4_S2 <=     O40_N8_S1  +  O40_N10_S1 ;
 logic signed [21:0] O40_N6_S2;		always @(posedge clk) O40_N6_S2 <=     O40_N12_S1  +  O40_N14_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O40_N0_S3;		always @(posedge clk) O40_N0_S3 <=     O40_N0_S2  +  O40_N2_S2 ;
 logic signed [22:0] O40_N2_S3;		always @(posedge clk) O40_N2_S3 <=     O40_N4_S2  +  O40_N6_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O40_N0_S4;		always @(posedge clk) O40_N0_S4 <=     O40_N0_S3  +  O40_N2_S3 ;
 assign conv_mac_40 = O40_N0_S4;

logic signed [31:0] conv_mac_41;
logic signed [63:0] chainout_0_O41; 
logic signed [63:0] O41_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O41(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_2[7:0]),.ay( 9'sd1),.bx(input_fmap_3[7:0]),.by( 9'sd1),.cx(input_fmap_4[7:0]),.cy(-9'sd2),.dx(input_fmap_5[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O41_N0_S1),.chainout(chainout_0_O41));
logic signed [63:0] chainout_2_O41; 
logic signed [63:0] O41_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O41(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_8[7:0]),.ay(-9'sd1),.bx(input_fmap_11[7:0]),.by(-9'sd1),.cx(input_fmap_12[7:0]),.cy(-9'sd1),.dx(input_fmap_13[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O41_N2_S1),.chainout(chainout_2_O41));
logic signed [63:0] chainout_4_O41; 
logic signed [63:0] O41_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O41(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_17[7:0]),.ay( 9'sd1),.bx(input_fmap_20[7:0]),.by( 9'sd1),.cx(input_fmap_23[7:0]),.cy( 9'sd1),.dx(input_fmap_27[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O41_N4_S1),.chainout(chainout_4_O41));
logic signed [63:0] chainout_6_O41; 
logic signed [63:0] O41_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O41(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_30[7:0]),.ay( 9'sd1),.bx(input_fmap_31[7:0]),.by( 9'sd2),.cx(input_fmap_33[7:0]),.cy( 9'sd1),.dx(input_fmap_36[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O41_N6_S1),.chainout(chainout_6_O41));
logic signed [63:0] chainout_8_O41; 
logic signed [63:0] O41_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O41(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_37[7:0]),.ay( 9'sd1),.bx(input_fmap_39[7:0]),.by( 9'sd2),.cx(input_fmap_40[7:0]),.cy( 9'sd1),.dx(input_fmap_42[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O41_N8_S1),.chainout(chainout_8_O41));
logic signed [63:0] chainout_10_O41; 
logic signed [63:0] O41_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O41(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_46[7:0]),.ay(-9'sd1),.bx(input_fmap_47[7:0]),.by( 9'sd2),.cx(input_fmap_48[7:0]),.cy(-9'sd1),.dx(input_fmap_51[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O41_N10_S1),.chainout(chainout_10_O41));
logic signed [63:0] chainout_12_O41; 
logic signed [63:0] O41_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O41(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_54[7:0]),.ay( 9'sd2),.bx(input_fmap_57[7:0]),.by( 9'sd1),.cx(input_fmap_58[7:0]),.cy(-9'sd1),.dx(input_fmap_61[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O41_N12_S1),.chainout(chainout_12_O41));
logic signed [63:0] chainout_14_O41; 
logic signed [63:0] O41_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O41(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_62[7:0]),.ay(-9'sd1),.bx(input_fmap_63[7:0]),.by( 9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O41_N14_S1),.chainout(chainout_14_O41));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O41_N0_S2;		always @(posedge clk) O41_N0_S2 <=     O41_N0_S1  +  O41_N2_S1 ;
 logic signed [21:0] O41_N2_S2;		always @(posedge clk) O41_N2_S2 <=     O41_N4_S1  +  O41_N6_S1 ;
 logic signed [21:0] O41_N4_S2;		always @(posedge clk) O41_N4_S2 <=     O41_N8_S1  +  O41_N10_S1 ;
 logic signed [21:0] O41_N6_S2;		always @(posedge clk) O41_N6_S2 <=     O41_N12_S1  +  O41_N14_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O41_N0_S3;		always @(posedge clk) O41_N0_S3 <=     O41_N0_S2  +  O41_N2_S2 ;
 logic signed [22:0] O41_N2_S3;		always @(posedge clk) O41_N2_S3 <=     O41_N4_S2  +  O41_N6_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O41_N0_S4;		always @(posedge clk) O41_N0_S4 <=     O41_N0_S3  +  O41_N2_S3 ;
 assign conv_mac_41 = O41_N0_S4;

logic signed [31:0] conv_mac_42;
logic signed [63:0] chainout_0_O42; 
logic signed [63:0] O42_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O42(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd1),.bx(input_fmap_4[7:0]),.by( 9'sd1),.cx(input_fmap_7[7:0]),.cy(-9'sd1),.dx(input_fmap_8[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O42_N0_S1),.chainout(chainout_0_O42));
logic signed [63:0] chainout_2_O42; 
logic signed [63:0] O42_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O42(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_10[7:0]),.ay(-9'sd1),.bx(input_fmap_11[7:0]),.by(-9'sd1),.cx(input_fmap_13[7:0]),.cy( 9'sd1),.dx(input_fmap_16[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O42_N2_S1),.chainout(chainout_2_O42));
logic signed [63:0] chainout_4_O42; 
logic signed [63:0] O42_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O42(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_17[7:0]),.ay(-9'sd1),.bx(input_fmap_18[7:0]),.by( 9'sd1),.cx(input_fmap_21[7:0]),.cy(-9'sd1),.dx(input_fmap_22[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O42_N4_S1),.chainout(chainout_4_O42));
logic signed [63:0] chainout_6_O42; 
logic signed [63:0] O42_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O42(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_23[7:0]),.ay(-9'sd1),.bx(input_fmap_24[7:0]),.by( 9'sd1),.cx(input_fmap_25[7:0]),.cy(-9'sd2),.dx(input_fmap_26[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O42_N6_S1),.chainout(chainout_6_O42));
logic signed [63:0] chainout_8_O42; 
logic signed [63:0] O42_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O42(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_27[7:0]),.ay(-9'sd1),.bx(input_fmap_29[7:0]),.by( 9'sd1),.cx(input_fmap_33[7:0]),.cy( 9'sd2),.dx(input_fmap_34[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O42_N8_S1),.chainout(chainout_8_O42));
logic signed [63:0] chainout_10_O42; 
logic signed [63:0] O42_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O42(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_35[7:0]),.ay(-9'sd1),.bx(input_fmap_36[7:0]),.by(-9'sd1),.cx(input_fmap_37[7:0]),.cy(-9'sd1),.dx(input_fmap_38[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O42_N10_S1),.chainout(chainout_10_O42));
logic signed [63:0] chainout_12_O42; 
logic signed [63:0] O42_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O42(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_39[7:0]),.ay( 9'sd1),.bx(input_fmap_42[7:0]),.by(-9'sd1),.cx(input_fmap_45[7:0]),.cy( 9'sd2),.dx(input_fmap_46[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O42_N12_S1),.chainout(chainout_12_O42));
logic signed [63:0] chainout_14_O42; 
logic signed [63:0] O42_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O42(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_47[7:0]),.ay(-9'sd2),.bx(input_fmap_50[7:0]),.by( 9'sd1),.cx(input_fmap_52[7:0]),.cy( 9'sd1),.dx(input_fmap_53[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O42_N14_S1),.chainout(chainout_14_O42));
logic signed [63:0] chainout_16_O42; 
logic signed [63:0] O42_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O42(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_55[7:0]),.ay(-9'sd1),.bx(input_fmap_57[7:0]),.by( 9'sd2),.cx(input_fmap_60[7:0]),.cy(-9'sd1),.dx(input_fmap_61[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O42_N16_S1),.chainout(chainout_16_O42));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O42_N0_S2;		always @(posedge clk) O42_N0_S2 <=     O42_N0_S1  +  O42_N2_S1 ;
 logic signed [21:0] O42_N2_S2;		always @(posedge clk) O42_N2_S2 <=     O42_N4_S1  +  O42_N6_S1 ;
 logic signed [21:0] O42_N4_S2;		always @(posedge clk) O42_N4_S2 <=     O42_N8_S1  +  O42_N10_S1 ;
 logic signed [21:0] O42_N6_S2;		always @(posedge clk) O42_N6_S2 <=     O42_N12_S1  +  O42_N14_S1 ;
 logic signed [21:0] O42_N8_S2;		always @(posedge clk) O42_N8_S2 <=     O42_N16_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O42_N0_S3;		always @(posedge clk) O42_N0_S3 <=     O42_N0_S2  +  O42_N2_S2 ;
 logic signed [22:0] O42_N2_S3;		always @(posedge clk) O42_N2_S3 <=     O42_N4_S2  +  O42_N6_S2 ;
 logic signed [22:0] O42_N4_S3;		always @(posedge clk) O42_N4_S3 <=     O42_N8_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O42_N0_S4;		always @(posedge clk) O42_N0_S4 <=     O42_N0_S3  +  O42_N2_S3 ;
 logic signed [23:0] O42_N2_S4;		always @(posedge clk) O42_N2_S4 <=     O42_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O42_N0_S5;		always @(posedge clk) O42_N0_S5 <=     O42_N0_S4  +  O42_N2_S4 ;
 assign conv_mac_42 = O42_N0_S5;

logic signed [31:0] conv_mac_43;
logic signed [63:0] chainout_0_O43; 
logic signed [63:0] O43_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O43(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay( 9'sd1),.bx(input_fmap_2[7:0]),.by(-9'sd1),.cx(input_fmap_3[7:0]),.cy(-9'sd1),.dx(input_fmap_4[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O43_N0_S1),.chainout(chainout_0_O43));
logic signed [63:0] chainout_2_O43; 
logic signed [63:0] O43_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O43(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_6[7:0]),.ay( 9'sd1),.bx(input_fmap_12[7:0]),.by( 9'sd1),.cx(input_fmap_13[7:0]),.cy(-9'sd1),.dx(input_fmap_15[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O43_N2_S1),.chainout(chainout_2_O43));
logic signed [63:0] chainout_4_O43; 
logic signed [63:0] O43_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O43(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_18[7:0]),.ay( 9'sd1),.bx(input_fmap_19[7:0]),.by( 9'sd1),.cx(input_fmap_21[7:0]),.cy( 9'sd1),.dx(input_fmap_22[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O43_N4_S1),.chainout(chainout_4_O43));
logic signed [63:0] chainout_6_O43; 
logic signed [63:0] O43_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O43(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_24[7:0]),.ay( 9'sd1),.bx(input_fmap_25[7:0]),.by( 9'sd1),.cx(input_fmap_26[7:0]),.cy( 9'sd1),.dx(input_fmap_29[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O43_N6_S1),.chainout(chainout_6_O43));
logic signed [63:0] chainout_8_O43; 
logic signed [63:0] O43_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O43(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_31[7:0]),.ay( 9'sd1),.bx(input_fmap_32[7:0]),.by(-9'sd1),.cx(input_fmap_33[7:0]),.cy(-9'sd1),.dx(input_fmap_34[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O43_N8_S1),.chainout(chainout_8_O43));
logic signed [63:0] chainout_10_O43; 
logic signed [63:0] O43_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O43(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_36[7:0]),.ay( 9'sd3),.bx(input_fmap_37[7:0]),.by( 9'sd2),.cx(input_fmap_38[7:0]),.cy( 9'sd1),.dx(input_fmap_40[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O43_N10_S1),.chainout(chainout_10_O43));
logic signed [63:0] chainout_12_O43; 
logic signed [63:0] O43_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O43(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_44[7:0]),.ay(-9'sd1),.bx(input_fmap_46[7:0]),.by(-9'sd2),.cx(input_fmap_49[7:0]),.cy( 9'sd2),.dx(input_fmap_51[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O43_N12_S1),.chainout(chainout_12_O43));
logic signed [63:0] chainout_14_O43; 
logic signed [63:0] O43_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O43(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_52[7:0]),.ay(-9'sd2),.bx(input_fmap_53[7:0]),.by( 9'sd1),.cx(input_fmap_60[7:0]),.cy(-9'sd1),.dx(input_fmap_61[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O43_N14_S1),.chainout(chainout_14_O43));
logic signed [63:0] chainout_16_O43; 
logic signed [63:0] O43_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O43(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_63[7:0]),.ay( 9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O43_N16_S1),.chainout(chainout_16_O43));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O43_N0_S2;		always @(posedge clk) O43_N0_S2 <=     O43_N0_S1  +  O43_N2_S1 ;
 logic signed [21:0] O43_N2_S2;		always @(posedge clk) O43_N2_S2 <=     O43_N4_S1  +  O43_N6_S1 ;
 logic signed [21:0] O43_N4_S2;		always @(posedge clk) O43_N4_S2 <=     O43_N8_S1  +  O43_N10_S1 ;
 logic signed [21:0] O43_N6_S2;		always @(posedge clk) O43_N6_S2 <=     O43_N12_S1  +  O43_N14_S1 ;
 logic signed [21:0] O43_N8_S2;		always @(posedge clk) O43_N8_S2 <=     O43_N16_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O43_N0_S3;		always @(posedge clk) O43_N0_S3 <=     O43_N0_S2  +  O43_N2_S2 ;
 logic signed [22:0] O43_N2_S3;		always @(posedge clk) O43_N2_S3 <=     O43_N4_S2  +  O43_N6_S2 ;
 logic signed [22:0] O43_N4_S3;		always @(posedge clk) O43_N4_S3 <=     O43_N8_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O43_N0_S4;		always @(posedge clk) O43_N0_S4 <=     O43_N0_S3  +  O43_N2_S3 ;
 logic signed [23:0] O43_N2_S4;		always @(posedge clk) O43_N2_S4 <=     O43_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O43_N0_S5;		always @(posedge clk) O43_N0_S5 <=     O43_N0_S4  +  O43_N2_S4 ;
 assign conv_mac_43 = O43_N0_S5;

logic signed [31:0] conv_mac_44;
logic signed [63:0] chainout_0_O44; 
logic signed [63:0] O44_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O44(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd1),.bx(input_fmap_1[7:0]),.by(-9'sd1),.cx(input_fmap_2[7:0]),.cy( 9'sd2),.dx(input_fmap_3[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O44_N0_S1),.chainout(chainout_0_O44));
logic signed [63:0] chainout_2_O44; 
logic signed [63:0] O44_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O44(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_4[7:0]),.ay(-9'sd1),.bx(input_fmap_6[7:0]),.by(-9'sd1),.cx(input_fmap_8[7:0]),.cy(-9'sd1),.dx(input_fmap_9[7:0]),.dy( 9'sd3),.chainin(63'd0),.result(O44_N2_S1),.chainout(chainout_2_O44));
logic signed [63:0] chainout_4_O44; 
logic signed [63:0] O44_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O44(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_10[7:0]),.ay( 9'sd3),.bx(input_fmap_12[7:0]),.by( 9'sd3),.cx(input_fmap_14[7:0]),.cy( 9'sd3),.dx(input_fmap_15[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O44_N4_S1),.chainout(chainout_4_O44));
logic signed [63:0] chainout_6_O44; 
logic signed [63:0] O44_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O44(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_17[7:0]),.ay( 9'sd1),.bx(input_fmap_18[7:0]),.by( 9'sd1),.cx(input_fmap_19[7:0]),.cy(-9'sd2),.dx(input_fmap_20[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O44_N6_S1),.chainout(chainout_6_O44));
logic signed [63:0] chainout_8_O44; 
logic signed [63:0] O44_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O44(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_22[7:0]),.ay( 9'sd1),.bx(input_fmap_23[7:0]),.by( 9'sd1),.cx(input_fmap_25[7:0]),.cy(-9'sd1),.dx(input_fmap_26[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O44_N8_S1),.chainout(chainout_8_O44));
logic signed [63:0] chainout_10_O44; 
logic signed [63:0] O44_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O44(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_27[7:0]),.ay( 9'sd1),.bx(input_fmap_28[7:0]),.by(-9'sd1),.cx(input_fmap_29[7:0]),.cy(-9'sd4),.dx(input_fmap_31[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O44_N10_S1),.chainout(chainout_10_O44));
logic signed [63:0] chainout_12_O44; 
logic signed [63:0] O44_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O44(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_32[7:0]),.ay(-9'sd1),.bx(input_fmap_33[7:0]),.by( 9'sd1),.cx(input_fmap_34[7:0]),.cy( 9'sd1),.dx(input_fmap_35[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O44_N12_S1),.chainout(chainout_12_O44));
logic signed [63:0] chainout_14_O44; 
logic signed [63:0] O44_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O44(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_37[7:0]),.ay( 9'sd2),.bx(input_fmap_38[7:0]),.by( 9'sd2),.cx(input_fmap_39[7:0]),.cy(-9'sd1),.dx(input_fmap_40[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O44_N14_S1),.chainout(chainout_14_O44));
logic signed [63:0] chainout_16_O44; 
logic signed [63:0] O44_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O44(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_41[7:0]),.ay(-9'sd4),.bx(input_fmap_42[7:0]),.by(-9'sd2),.cx(input_fmap_43[7:0]),.cy(-9'sd1),.dx(input_fmap_44[7:0]),.dy(-9'sd3),.chainin(63'd0),.result(O44_N16_S1),.chainout(chainout_16_O44));
logic signed [63:0] chainout_18_O44; 
logic signed [63:0] O44_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O44(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_45[7:0]),.ay( 9'sd2),.bx(input_fmap_46[7:0]),.by(-9'sd3),.cx(input_fmap_47[7:0]),.cy( 9'sd2),.dx(input_fmap_49[7:0]),.dy( 9'sd6),.chainin(63'd0),.result(O44_N18_S1),.chainout(chainout_18_O44));
logic signed [63:0] chainout_20_O44; 
logic signed [63:0] O44_N20_S1; 
 int_sop_4_wrapper int_sop_4_inst_20_O44(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_50[7:0]),.ay( 9'sd1),.bx(input_fmap_51[7:0]),.by( 9'sd3),.cx(input_fmap_52[7:0]),.cy(-9'sd1),.dx(input_fmap_54[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O44_N20_S1),.chainout(chainout_20_O44));
logic signed [63:0] chainout_22_O44; 
logic signed [63:0] O44_N22_S1; 
 int_sop_4_wrapper int_sop_4_inst_22_O44(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_55[7:0]),.ay( 9'sd1),.bx(input_fmap_56[7:0]),.by(-9'sd2),.cx(input_fmap_58[7:0]),.cy(-9'sd1),.dx(input_fmap_59[7:0]),.dy( 9'sd4),.chainin(63'd0),.result(O44_N22_S1),.chainout(chainout_22_O44));
logic signed [63:0] chainout_24_O44; 
logic signed [63:0] O44_N24_S1; 
 int_sop_4_wrapper int_sop_4_inst_24_O44(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_60[7:0]),.ay( 9'sd1),.bx(input_fmap_61[7:0]),.by(-9'sd2),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O44_N24_S1),.chainout(chainout_24_O44));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O44_N0_S2;		always @(posedge clk) O44_N0_S2 <=     O44_N0_S1  +  O44_N2_S1 ;
 logic signed [21:0] O44_N2_S2;		always @(posedge clk) O44_N2_S2 <=     O44_N4_S1  +  O44_N6_S1 ;
 logic signed [21:0] O44_N4_S2;		always @(posedge clk) O44_N4_S2 <=     O44_N8_S1  +  O44_N10_S1 ;
 logic signed [21:0] O44_N6_S2;		always @(posedge clk) O44_N6_S2 <=     O44_N12_S1  +  O44_N14_S1 ;
 logic signed [21:0] O44_N8_S2;		always @(posedge clk) O44_N8_S2 <=     O44_N16_S1  +  O44_N18_S1 ;
 logic signed [21:0] O44_N10_S2;		always @(posedge clk) O44_N10_S2 <=     O44_N20_S1  +  O44_N22_S1 ;
 logic signed [21:0] O44_N12_S2;		always @(posedge clk) O44_N12_S2 <=     O44_N24_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O44_N0_S3;		always @(posedge clk) O44_N0_S3 <=     O44_N0_S2  +  O44_N2_S2 ;
 logic signed [22:0] O44_N2_S3;		always @(posedge clk) O44_N2_S3 <=     O44_N4_S2  +  O44_N6_S2 ;
 logic signed [22:0] O44_N4_S3;		always @(posedge clk) O44_N4_S3 <=     O44_N8_S2  +  O44_N10_S2 ;
 logic signed [22:0] O44_N6_S3;		always @(posedge clk) O44_N6_S3 <=     O44_N12_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O44_N0_S4;		always @(posedge clk) O44_N0_S4 <=     O44_N0_S3  +  O44_N2_S3 ;
 logic signed [23:0] O44_N2_S4;		always @(posedge clk) O44_N2_S4 <=     O44_N4_S3  +  O44_N6_S3 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O44_N0_S5;		always @(posedge clk) O44_N0_S5 <=     O44_N0_S4  +  O44_N2_S4 ;
 assign conv_mac_44 = O44_N0_S5;

logic signed [31:0] conv_mac_45;
logic signed [63:0] chainout_0_O45; 
logic signed [63:0] O45_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O45(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd1),.bx(input_fmap_1[7:0]),.by(-9'sd1),.cx(input_fmap_2[7:0]),.cy(-9'sd1),.dx(input_fmap_3[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O45_N0_S1),.chainout(chainout_0_O45));
logic signed [63:0] chainout_2_O45; 
logic signed [63:0] O45_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O45(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_4[7:0]),.ay(-9'sd2),.bx(input_fmap_5[7:0]),.by(-9'sd1),.cx(input_fmap_7[7:0]),.cy(-9'sd1),.dx(input_fmap_8[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O45_N2_S1),.chainout(chainout_2_O45));
logic signed [63:0] chainout_4_O45; 
logic signed [63:0] O45_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O45(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_9[7:0]),.ay( 9'sd1),.bx(input_fmap_10[7:0]),.by(-9'sd1),.cx(input_fmap_11[7:0]),.cy(-9'sd1),.dx(input_fmap_12[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O45_N4_S1),.chainout(chainout_4_O45));
logic signed [63:0] chainout_6_O45; 
logic signed [63:0] O45_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O45(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_13[7:0]),.ay(-9'sd1),.bx(input_fmap_14[7:0]),.by(-9'sd2),.cx(input_fmap_15[7:0]),.cy( 9'sd1),.dx(input_fmap_16[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O45_N6_S1),.chainout(chainout_6_O45));
logic signed [63:0] chainout_8_O45; 
logic signed [63:0] O45_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O45(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_17[7:0]),.ay(-9'sd1),.bx(input_fmap_21[7:0]),.by(-9'sd1),.cx(input_fmap_23[7:0]),.cy( 9'sd1),.dx(input_fmap_24[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O45_N8_S1),.chainout(chainout_8_O45));
logic signed [63:0] chainout_10_O45; 
logic signed [63:0] O45_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O45(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_27[7:0]),.ay( 9'sd2),.bx(input_fmap_28[7:0]),.by(-9'sd2),.cx(input_fmap_29[7:0]),.cy(-9'sd1),.dx(input_fmap_30[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O45_N10_S1),.chainout(chainout_10_O45));
logic signed [63:0] chainout_12_O45; 
logic signed [63:0] O45_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O45(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_32[7:0]),.ay( 9'sd1),.bx(input_fmap_33[7:0]),.by(-9'sd1),.cx(input_fmap_34[7:0]),.cy( 9'sd1),.dx(input_fmap_35[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O45_N12_S1),.chainout(chainout_12_O45));
logic signed [63:0] chainout_14_O45; 
logic signed [63:0] O45_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O45(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_37[7:0]),.ay( 9'sd1),.bx(input_fmap_38[7:0]),.by( 9'sd1),.cx(input_fmap_39[7:0]),.cy( 9'sd1),.dx(input_fmap_40[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O45_N14_S1),.chainout(chainout_14_O45));
logic signed [63:0] chainout_16_O45; 
logic signed [63:0] O45_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O45(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_42[7:0]),.ay( 9'sd1),.bx(input_fmap_44[7:0]),.by(-9'sd1),.cx(input_fmap_47[7:0]),.cy( 9'sd1),.dx(input_fmap_48[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O45_N16_S1),.chainout(chainout_16_O45));
logic signed [63:0] chainout_18_O45; 
logic signed [63:0] O45_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O45(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_52[7:0]),.ay(-9'sd1),.bx(input_fmap_53[7:0]),.by(-9'sd1),.cx(input_fmap_54[7:0]),.cy( 9'sd2),.dx(input_fmap_56[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O45_N18_S1),.chainout(chainout_18_O45));
logic signed [63:0] chainout_20_O45; 
logic signed [63:0] O45_N20_S1; 
 int_sop_4_wrapper int_sop_4_inst_20_O45(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_57[7:0]),.ay( 9'sd1),.bx(input_fmap_58[7:0]),.by( 9'sd1),.cx(input_fmap_59[7:0]),.cy(-9'sd2),.dx(input_fmap_60[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O45_N20_S1),.chainout(chainout_20_O45));
logic signed [63:0] chainout_22_O45; 
logic signed [63:0] O45_N22_S1; 
 int_sop_4_wrapper int_sop_4_inst_22_O45(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_61[7:0]),.ay( 9'sd6),.bx(input_fmap_62[7:0]),.by(-9'sd1),.cx(input_fmap_63[7:0]),.cy( 9'sd2),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O45_N22_S1),.chainout(chainout_22_O45));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O45_N0_S2;		always @(posedge clk) O45_N0_S2 <=     O45_N0_S1  +  O45_N2_S1 ;
 logic signed [21:0] O45_N2_S2;		always @(posedge clk) O45_N2_S2 <=     O45_N4_S1  +  O45_N6_S1 ;
 logic signed [21:0] O45_N4_S2;		always @(posedge clk) O45_N4_S2 <=     O45_N8_S1  +  O45_N10_S1 ;
 logic signed [21:0] O45_N6_S2;		always @(posedge clk) O45_N6_S2 <=     O45_N12_S1  +  O45_N14_S1 ;
 logic signed [21:0] O45_N8_S2;		always @(posedge clk) O45_N8_S2 <=     O45_N16_S1  +  O45_N18_S1 ;
 logic signed [21:0] O45_N10_S2;		always @(posedge clk) O45_N10_S2 <=     O45_N20_S1  +  O45_N22_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O45_N0_S3;		always @(posedge clk) O45_N0_S3 <=     O45_N0_S2  +  O45_N2_S2 ;
 logic signed [22:0] O45_N2_S3;		always @(posedge clk) O45_N2_S3 <=     O45_N4_S2  +  O45_N6_S2 ;
 logic signed [22:0] O45_N4_S3;		always @(posedge clk) O45_N4_S3 <=     O45_N8_S2  +  O45_N10_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O45_N0_S4;		always @(posedge clk) O45_N0_S4 <=     O45_N0_S3  +  O45_N2_S3 ;
 logic signed [23:0] O45_N2_S4;		always @(posedge clk) O45_N2_S4 <=     O45_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O45_N0_S5;		always @(posedge clk) O45_N0_S5 <=     O45_N0_S4  +  O45_N2_S4 ;
 assign conv_mac_45 = O45_N0_S5;

logic signed [31:0] conv_mac_46;
logic signed [63:0] chainout_0_O46; 
logic signed [63:0] O46_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O46(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_2[7:0]),.ay( 9'sd2),.bx(input_fmap_3[7:0]),.by( 9'sd1),.cx(input_fmap_10[7:0]),.cy(-9'sd1),.dx(input_fmap_11[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O46_N0_S1),.chainout(chainout_0_O46));
logic signed [63:0] chainout_2_O46; 
logic signed [63:0] O46_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O46(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_13[7:0]),.ay( 9'sd1),.bx(input_fmap_14[7:0]),.by( 9'sd1),.cx(input_fmap_18[7:0]),.cy(-9'sd1),.dx(input_fmap_20[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O46_N2_S1),.chainout(chainout_2_O46));
logic signed [63:0] chainout_4_O46; 
logic signed [63:0] O46_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O46(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_22[7:0]),.ay( 9'sd1),.bx(input_fmap_26[7:0]),.by( 9'sd1),.cx(input_fmap_28[7:0]),.cy(-9'sd1),.dx(input_fmap_30[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O46_N4_S1),.chainout(chainout_4_O46));
logic signed [63:0] chainout_6_O46; 
logic signed [63:0] O46_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O46(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_31[7:0]),.ay(-9'sd1),.bx(input_fmap_37[7:0]),.by( 9'sd1),.cx(input_fmap_48[7:0]),.cy( 9'sd1),.dx(input_fmap_50[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O46_N6_S1),.chainout(chainout_6_O46));
logic signed [63:0] chainout_8_O46; 
logic signed [63:0] O46_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O46(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_52[7:0]),.ay( 9'sd1),.bx(input_fmap_53[7:0]),.by(-9'sd1),.cx(input_fmap_56[7:0]),.cy( 9'sd1),.dx(input_fmap_59[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O46_N8_S1),.chainout(chainout_8_O46));
logic signed [63:0] chainout_10_O46; 
logic signed [63:0] O46_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O46(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_63[7:0]),.ay(-9'sd2),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O46_N10_S1),.chainout(chainout_10_O46));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O46_N0_S2;		always @(posedge clk) O46_N0_S2 <=     O46_N0_S1  +  O46_N2_S1 ;
 logic signed [21:0] O46_N2_S2;		always @(posedge clk) O46_N2_S2 <=     O46_N4_S1  +  O46_N6_S1 ;
 logic signed [21:0] O46_N4_S2;		always @(posedge clk) O46_N4_S2 <=     O46_N8_S1  +  O46_N10_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O46_N0_S3;		always @(posedge clk) O46_N0_S3 <=     O46_N0_S2  +  O46_N2_S2 ;
 logic signed [22:0] O46_N2_S3;		always @(posedge clk) O46_N2_S3 <=     O46_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O46_N0_S4;		always @(posedge clk) O46_N0_S4 <=     O46_N0_S3  +  O46_N2_S3 ;
 assign conv_mac_46 = O46_N0_S4;

logic signed [31:0] conv_mac_47;
logic signed [63:0] chainout_0_O47; 
logic signed [63:0] O47_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O47(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd1),.bx(input_fmap_3[7:0]),.by( 9'sd1),.cx(input_fmap_4[7:0]),.cy( 9'sd1),.dx(input_fmap_10[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O47_N0_S1),.chainout(chainout_0_O47));
logic signed [63:0] chainout_2_O47; 
logic signed [63:0] O47_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O47(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_12[7:0]),.ay( 9'sd1),.bx(input_fmap_13[7:0]),.by( 9'sd1),.cx(input_fmap_15[7:0]),.cy(-9'sd1),.dx(input_fmap_17[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O47_N2_S1),.chainout(chainout_2_O47));
logic signed [63:0] chainout_4_O47; 
logic signed [63:0] O47_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O47(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_19[7:0]),.ay(-9'sd1),.bx(input_fmap_21[7:0]),.by( 9'sd1),.cx(input_fmap_25[7:0]),.cy( 9'sd1),.dx(input_fmap_26[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O47_N4_S1),.chainout(chainout_4_O47));
logic signed [63:0] chainout_6_O47; 
logic signed [63:0] O47_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O47(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_27[7:0]),.ay(-9'sd1),.bx(input_fmap_31[7:0]),.by(-9'sd1),.cx(input_fmap_32[7:0]),.cy( 9'sd1),.dx(input_fmap_33[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O47_N6_S1),.chainout(chainout_6_O47));
logic signed [63:0] chainout_8_O47; 
logic signed [63:0] O47_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O47(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_34[7:0]),.ay( 9'sd1),.bx(input_fmap_40[7:0]),.by( 9'sd2),.cx(input_fmap_41[7:0]),.cy(-9'sd1),.dx(input_fmap_43[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O47_N8_S1),.chainout(chainout_8_O47));
logic signed [63:0] chainout_10_O47; 
logic signed [63:0] O47_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O47(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_45[7:0]),.ay( 9'sd1),.bx(input_fmap_46[7:0]),.by(-9'sd1),.cx(input_fmap_48[7:0]),.cy(-9'sd1),.dx(input_fmap_49[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O47_N10_S1),.chainout(chainout_10_O47));
logic signed [63:0] chainout_12_O47; 
logic signed [63:0] O47_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O47(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_50[7:0]),.ay( 9'sd1),.bx(input_fmap_52[7:0]),.by(-9'sd1),.cx(input_fmap_53[7:0]),.cy( 9'sd1),.dx(input_fmap_55[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O47_N12_S1),.chainout(chainout_12_O47));
logic signed [63:0] chainout_14_O47; 
logic signed [63:0] O47_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O47(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_59[7:0]),.ay(-9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O47_N14_S1),.chainout(chainout_14_O47));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O47_N0_S2;		always @(posedge clk) O47_N0_S2 <=     O47_N0_S1  +  O47_N2_S1 ;
 logic signed [21:0] O47_N2_S2;		always @(posedge clk) O47_N2_S2 <=     O47_N4_S1  +  O47_N6_S1 ;
 logic signed [21:0] O47_N4_S2;		always @(posedge clk) O47_N4_S2 <=     O47_N8_S1  +  O47_N10_S1 ;
 logic signed [21:0] O47_N6_S2;		always @(posedge clk) O47_N6_S2 <=     O47_N12_S1  +  O47_N14_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O47_N0_S3;		always @(posedge clk) O47_N0_S3 <=     O47_N0_S2  +  O47_N2_S2 ;
 logic signed [22:0] O47_N2_S3;		always @(posedge clk) O47_N2_S3 <=     O47_N4_S2  +  O47_N6_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O47_N0_S4;		always @(posedge clk) O47_N0_S4 <=     O47_N0_S3  +  O47_N2_S3 ;
 assign conv_mac_47 = O47_N0_S4;

logic signed [31:0] conv_mac_48;
logic signed [63:0] chainout_0_O48; 
logic signed [63:0] O48_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O48(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd1),.bx(input_fmap_1[7:0]),.by(-9'sd1),.cx(input_fmap_2[7:0]),.cy( 9'sd2),.dx(input_fmap_3[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O48_N0_S1),.chainout(chainout_0_O48));
logic signed [63:0] chainout_2_O48; 
logic signed [63:0] O48_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O48(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_4[7:0]),.ay( 9'sd1),.bx(input_fmap_6[7:0]),.by(-9'sd1),.cx(input_fmap_8[7:0]),.cy(-9'sd1),.dx(input_fmap_10[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O48_N2_S1),.chainout(chainout_2_O48));
logic signed [63:0] chainout_4_O48; 
logic signed [63:0] O48_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O48(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_11[7:0]),.ay(-9'sd1),.bx(input_fmap_12[7:0]),.by( 9'sd1),.cx(input_fmap_13[7:0]),.cy( 9'sd1),.dx(input_fmap_14[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O48_N4_S1),.chainout(chainout_4_O48));
logic signed [63:0] chainout_6_O48; 
logic signed [63:0] O48_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O48(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_15[7:0]),.ay( 9'sd1),.bx(input_fmap_16[7:0]),.by(-9'sd3),.cx(input_fmap_17[7:0]),.cy(-9'sd1),.dx(input_fmap_18[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O48_N6_S1),.chainout(chainout_6_O48));
logic signed [63:0] chainout_8_O48; 
logic signed [63:0] O48_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O48(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_21[7:0]),.ay( 9'sd2),.bx(input_fmap_24[7:0]),.by(-9'sd2),.cx(input_fmap_25[7:0]),.cy(-9'sd2),.dx(input_fmap_26[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O48_N8_S1),.chainout(chainout_8_O48));
logic signed [63:0] chainout_10_O48; 
logic signed [63:0] O48_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O48(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_28[7:0]),.ay(-9'sd1),.bx(input_fmap_31[7:0]),.by( 9'sd1),.cx(input_fmap_32[7:0]),.cy( 9'sd1),.dx(input_fmap_33[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O48_N10_S1),.chainout(chainout_10_O48));
logic signed [63:0] chainout_12_O48; 
logic signed [63:0] O48_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O48(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_34[7:0]),.ay(-9'sd2),.bx(input_fmap_35[7:0]),.by( 9'sd2),.cx(input_fmap_36[7:0]),.cy(-9'sd1),.dx(input_fmap_37[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O48_N12_S1),.chainout(chainout_12_O48));
logic signed [63:0] chainout_14_O48; 
logic signed [63:0] O48_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O48(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_38[7:0]),.ay( 9'sd1),.bx(input_fmap_39[7:0]),.by(-9'sd1),.cx(input_fmap_41[7:0]),.cy( 9'sd1),.dx(input_fmap_42[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O48_N14_S1),.chainout(chainout_14_O48));
logic signed [63:0] chainout_16_O48; 
logic signed [63:0] O48_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O48(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_43[7:0]),.ay(-9'sd2),.bx(input_fmap_45[7:0]),.by(-9'sd3),.cx(input_fmap_46[7:0]),.cy(-9'sd1),.dx(input_fmap_47[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O48_N16_S1),.chainout(chainout_16_O48));
logic signed [63:0] chainout_18_O48; 
logic signed [63:0] O48_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O48(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_49[7:0]),.ay(-9'sd1),.bx(input_fmap_50[7:0]),.by(-9'sd1),.cx(input_fmap_53[7:0]),.cy(-9'sd1),.dx(input_fmap_54[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O48_N18_S1),.chainout(chainout_18_O48));
logic signed [63:0] chainout_20_O48; 
logic signed [63:0] O48_N20_S1; 
 int_sop_4_wrapper int_sop_4_inst_20_O48(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_56[7:0]),.ay( 9'sd1),.bx(input_fmap_59[7:0]),.by(-9'sd1),.cx(input_fmap_60[7:0]),.cy(-9'sd2),.dx(input_fmap_61[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O48_N20_S1),.chainout(chainout_20_O48));
logic signed [63:0] chainout_22_O48; 
logic signed [63:0] O48_N22_S1; 
 int_sop_4_wrapper int_sop_4_inst_22_O48(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_62[7:0]),.ay( 9'sd1),.bx(input_fmap_63[7:0]),.by( 9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O48_N22_S1),.chainout(chainout_22_O48));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O48_N0_S2;		always @(posedge clk) O48_N0_S2 <=     O48_N0_S1  +  O48_N2_S1 ;
 logic signed [21:0] O48_N2_S2;		always @(posedge clk) O48_N2_S2 <=     O48_N4_S1  +  O48_N6_S1 ;
 logic signed [21:0] O48_N4_S2;		always @(posedge clk) O48_N4_S2 <=     O48_N8_S1  +  O48_N10_S1 ;
 logic signed [21:0] O48_N6_S2;		always @(posedge clk) O48_N6_S2 <=     O48_N12_S1  +  O48_N14_S1 ;
 logic signed [21:0] O48_N8_S2;		always @(posedge clk) O48_N8_S2 <=     O48_N16_S1  +  O48_N18_S1 ;
 logic signed [21:0] O48_N10_S2;		always @(posedge clk) O48_N10_S2 <=     O48_N20_S1  +  O48_N22_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O48_N0_S3;		always @(posedge clk) O48_N0_S3 <=     O48_N0_S2  +  O48_N2_S2 ;
 logic signed [22:0] O48_N2_S3;		always @(posedge clk) O48_N2_S3 <=     O48_N4_S2  +  O48_N6_S2 ;
 logic signed [22:0] O48_N4_S3;		always @(posedge clk) O48_N4_S3 <=     O48_N8_S2  +  O48_N10_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O48_N0_S4;		always @(posedge clk) O48_N0_S4 <=     O48_N0_S3  +  O48_N2_S3 ;
 logic signed [23:0] O48_N2_S4;		always @(posedge clk) O48_N2_S4 <=     O48_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O48_N0_S5;		always @(posedge clk) O48_N0_S5 <=     O48_N0_S4  +  O48_N2_S4 ;
 assign conv_mac_48 = O48_N0_S5;

logic signed [31:0] conv_mac_49;
logic signed [63:0] chainout_0_O49; 
logic signed [63:0] O49_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O49(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd2),.bx(input_fmap_4[7:0]),.by( 9'sd3),.cx(input_fmap_5[7:0]),.cy(-9'sd1),.dx(input_fmap_6[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O49_N0_S1),.chainout(chainout_0_O49));
logic signed [63:0] chainout_2_O49; 
logic signed [63:0] O49_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O49(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_7[7:0]),.ay( 9'sd1),.bx(input_fmap_10[7:0]),.by(-9'sd1),.cx(input_fmap_11[7:0]),.cy( 9'sd1),.dx(input_fmap_12[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O49_N2_S1),.chainout(chainout_2_O49));
logic signed [63:0] chainout_4_O49; 
logic signed [63:0] O49_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O49(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_13[7:0]),.ay( 9'sd1),.bx(input_fmap_17[7:0]),.by( 9'sd1),.cx(input_fmap_19[7:0]),.cy( 9'sd1),.dx(input_fmap_21[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O49_N4_S1),.chainout(chainout_4_O49));
logic signed [63:0] chainout_6_O49; 
logic signed [63:0] O49_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O49(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_23[7:0]),.ay(-9'sd1),.bx(input_fmap_24[7:0]),.by( 9'sd2),.cx(input_fmap_25[7:0]),.cy( 9'sd1),.dx(input_fmap_26[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O49_N6_S1),.chainout(chainout_6_O49));
logic signed [63:0] chainout_8_O49; 
logic signed [63:0] O49_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O49(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_27[7:0]),.ay( 9'sd1),.bx(input_fmap_28[7:0]),.by(-9'sd1),.cx(input_fmap_29[7:0]),.cy(-9'sd1),.dx(input_fmap_31[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O49_N8_S1),.chainout(chainout_8_O49));
logic signed [63:0] chainout_10_O49; 
logic signed [63:0] O49_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O49(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_32[7:0]),.ay( 9'sd3),.bx(input_fmap_33[7:0]),.by( 9'sd1),.cx(input_fmap_34[7:0]),.cy(-9'sd1),.dx(input_fmap_35[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O49_N10_S1),.chainout(chainout_10_O49));
logic signed [63:0] chainout_12_O49; 
logic signed [63:0] O49_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O49(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_36[7:0]),.ay(-9'sd1),.bx(input_fmap_38[7:0]),.by(-9'sd1),.cx(input_fmap_40[7:0]),.cy( 9'sd1),.dx(input_fmap_42[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O49_N12_S1),.chainout(chainout_12_O49));
logic signed [63:0] chainout_14_O49; 
logic signed [63:0] O49_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O49(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_43[7:0]),.ay( 9'sd1),.bx(input_fmap_46[7:0]),.by(-9'sd1),.cx(input_fmap_47[7:0]),.cy(-9'sd1),.dx(input_fmap_49[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O49_N14_S1),.chainout(chainout_14_O49));
logic signed [63:0] chainout_16_O49; 
logic signed [63:0] O49_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O49(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_53[7:0]),.ay( 9'sd1),.bx(input_fmap_54[7:0]),.by(-9'sd1),.cx(input_fmap_58[7:0]),.cy(-9'sd1),.dx(input_fmap_59[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O49_N16_S1),.chainout(chainout_16_O49));
logic signed [63:0] chainout_18_O49; 
logic signed [63:0] O49_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O49(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_61[7:0]),.ay(-9'sd2),.bx(input_fmap_62[7:0]),.by( 9'sd2),.cx(input_fmap_63[7:0]),.cy( 9'sd1),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O49_N18_S1),.chainout(chainout_18_O49));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O49_N0_S2;		always @(posedge clk) O49_N0_S2 <=     O49_N0_S1  +  O49_N2_S1 ;
 logic signed [21:0] O49_N2_S2;		always @(posedge clk) O49_N2_S2 <=     O49_N4_S1  +  O49_N6_S1 ;
 logic signed [21:0] O49_N4_S2;		always @(posedge clk) O49_N4_S2 <=     O49_N8_S1  +  O49_N10_S1 ;
 logic signed [21:0] O49_N6_S2;		always @(posedge clk) O49_N6_S2 <=     O49_N12_S1  +  O49_N14_S1 ;
 logic signed [21:0] O49_N8_S2;		always @(posedge clk) O49_N8_S2 <=     O49_N16_S1  +  O49_N18_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O49_N0_S3;		always @(posedge clk) O49_N0_S3 <=     O49_N0_S2  +  O49_N2_S2 ;
 logic signed [22:0] O49_N2_S3;		always @(posedge clk) O49_N2_S3 <=     O49_N4_S2  +  O49_N6_S2 ;
 logic signed [22:0] O49_N4_S3;		always @(posedge clk) O49_N4_S3 <=     O49_N8_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O49_N0_S4;		always @(posedge clk) O49_N0_S4 <=     O49_N0_S3  +  O49_N2_S3 ;
 logic signed [23:0] O49_N2_S4;		always @(posedge clk) O49_N2_S4 <=     O49_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O49_N0_S5;		always @(posedge clk) O49_N0_S5 <=     O49_N0_S4  +  O49_N2_S4 ;
 assign conv_mac_49 = O49_N0_S5;

logic signed [31:0] conv_mac_50;
logic signed [63:0] chainout_0_O50; 
logic signed [63:0] O50_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O50(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd1),.bx(input_fmap_1[7:0]),.by(-9'sd1),.cx(input_fmap_4[7:0]),.cy( 9'sd1),.dx(input_fmap_6[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O50_N0_S1),.chainout(chainout_0_O50));
logic signed [63:0] chainout_2_O50; 
logic signed [63:0] O50_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O50(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_9[7:0]),.ay(-9'sd2),.bx(input_fmap_10[7:0]),.by(-9'sd1),.cx(input_fmap_12[7:0]),.cy(-9'sd1),.dx(input_fmap_13[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O50_N2_S1),.chainout(chainout_2_O50));
logic signed [63:0] chainout_4_O50; 
logic signed [63:0] O50_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O50(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_14[7:0]),.ay( 9'sd1),.bx(input_fmap_16[7:0]),.by(-9'sd1),.cx(input_fmap_17[7:0]),.cy(-9'sd1),.dx(input_fmap_21[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O50_N4_S1),.chainout(chainout_4_O50));
logic signed [63:0] chainout_6_O50; 
logic signed [63:0] O50_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O50(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_23[7:0]),.ay( 9'sd4),.bx(input_fmap_29[7:0]),.by( 9'sd2),.cx(input_fmap_30[7:0]),.cy( 9'sd3),.dx(input_fmap_31[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O50_N6_S1),.chainout(chainout_6_O50));
logic signed [63:0] chainout_8_O50; 
logic signed [63:0] O50_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O50(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_32[7:0]),.ay(-9'sd1),.bx(input_fmap_34[7:0]),.by( 9'sd1),.cx(input_fmap_35[7:0]),.cy(-9'sd1),.dx(input_fmap_38[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O50_N8_S1),.chainout(chainout_8_O50));
logic signed [63:0] chainout_10_O50; 
logic signed [63:0] O50_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O50(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_39[7:0]),.ay( 9'sd1),.bx(input_fmap_42[7:0]),.by(-9'sd1),.cx(input_fmap_43[7:0]),.cy(-9'sd1),.dx(input_fmap_45[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O50_N10_S1),.chainout(chainout_10_O50));
logic signed [63:0] chainout_12_O50; 
logic signed [63:0] O50_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O50(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_48[7:0]),.ay( 9'sd2),.bx(input_fmap_49[7:0]),.by(-9'sd1),.cx(input_fmap_50[7:0]),.cy( 9'sd1),.dx(input_fmap_51[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O50_N12_S1),.chainout(chainout_12_O50));
logic signed [63:0] chainout_14_O50; 
logic signed [63:0] O50_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O50(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_55[7:0]),.ay(-9'sd1),.bx(input_fmap_56[7:0]),.by(-9'sd2),.cx(input_fmap_58[7:0]),.cy( 9'sd1),.dx(input_fmap_60[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O50_N14_S1),.chainout(chainout_14_O50));
logic signed [63:0] chainout_16_O50; 
logic signed [63:0] O50_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O50(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_61[7:0]),.ay(-9'sd3),.bx(input_fmap_62[7:0]),.by( 9'sd2),.cx(input_fmap_63[7:0]),.cy( 9'sd1),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O50_N16_S1),.chainout(chainout_16_O50));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O50_N0_S2;		always @(posedge clk) O50_N0_S2 <=     O50_N0_S1  +  O50_N2_S1 ;
 logic signed [21:0] O50_N2_S2;		always @(posedge clk) O50_N2_S2 <=     O50_N4_S1  +  O50_N6_S1 ;
 logic signed [21:0] O50_N4_S2;		always @(posedge clk) O50_N4_S2 <=     O50_N8_S1  +  O50_N10_S1 ;
 logic signed [21:0] O50_N6_S2;		always @(posedge clk) O50_N6_S2 <=     O50_N12_S1  +  O50_N14_S1 ;
 logic signed [21:0] O50_N8_S2;		always @(posedge clk) O50_N8_S2 <=     O50_N16_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O50_N0_S3;		always @(posedge clk) O50_N0_S3 <=     O50_N0_S2  +  O50_N2_S2 ;
 logic signed [22:0] O50_N2_S3;		always @(posedge clk) O50_N2_S3 <=     O50_N4_S2  +  O50_N6_S2 ;
 logic signed [22:0] O50_N4_S3;		always @(posedge clk) O50_N4_S3 <=     O50_N8_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O50_N0_S4;		always @(posedge clk) O50_N0_S4 <=     O50_N0_S3  +  O50_N2_S3 ;
 logic signed [23:0] O50_N2_S4;		always @(posedge clk) O50_N2_S4 <=     O50_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O50_N0_S5;		always @(posedge clk) O50_N0_S5 <=     O50_N0_S4  +  O50_N2_S4 ;
 assign conv_mac_50 = O50_N0_S5;

logic signed [31:0] conv_mac_51;
logic signed [63:0] chainout_0_O51; 
logic signed [63:0] O51_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O51(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_3[7:0]),.ay(-9'sd1),.bx(input_fmap_4[7:0]),.by( 9'sd4),.cx(input_fmap_7[7:0]),.cy( 9'sd1),.dx(input_fmap_8[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O51_N0_S1),.chainout(chainout_0_O51));
logic signed [63:0] chainout_2_O51; 
logic signed [63:0] O51_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O51(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_10[7:0]),.ay(-9'sd2),.bx(input_fmap_12[7:0]),.by( 9'sd2),.cx(input_fmap_13[7:0]),.cy(-9'sd1),.dx(input_fmap_14[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O51_N2_S1),.chainout(chainout_2_O51));
logic signed [63:0] chainout_4_O51; 
logic signed [63:0] O51_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O51(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_15[7:0]),.ay(-9'sd1),.bx(input_fmap_16[7:0]),.by( 9'sd1),.cx(input_fmap_17[7:0]),.cy(-9'sd1),.dx(input_fmap_19[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O51_N4_S1),.chainout(chainout_4_O51));
logic signed [63:0] chainout_6_O51; 
logic signed [63:0] O51_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O51(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_23[7:0]),.ay( 9'sd1),.bx(input_fmap_27[7:0]),.by(-9'sd1),.cx(input_fmap_31[7:0]),.cy(-9'sd1),.dx(input_fmap_33[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O51_N6_S1),.chainout(chainout_6_O51));
logic signed [63:0] chainout_8_O51; 
logic signed [63:0] O51_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O51(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_34[7:0]),.ay( 9'sd2),.bx(input_fmap_36[7:0]),.by( 9'sd1),.cx(input_fmap_39[7:0]),.cy( 9'sd3),.dx(input_fmap_43[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O51_N8_S1),.chainout(chainout_8_O51));
logic signed [63:0] chainout_10_O51; 
logic signed [63:0] O51_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O51(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_51[7:0]),.ay(-9'sd2),.bx(input_fmap_52[7:0]),.by(-9'sd1),.cx(input_fmap_54[7:0]),.cy( 9'sd2),.dx(input_fmap_60[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O51_N10_S1),.chainout(chainout_10_O51));
logic signed [63:0] chainout_12_O51; 
logic signed [63:0] O51_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O51(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_61[7:0]),.ay(-9'sd1),.bx(input_fmap_62[7:0]),.by( 9'sd3),.cx(input_fmap_63[7:0]),.cy( 9'sd1),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O51_N12_S1),.chainout(chainout_12_O51));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O51_N0_S2;		always @(posedge clk) O51_N0_S2 <=     O51_N0_S1  +  O51_N2_S1 ;
 logic signed [21:0] O51_N2_S2;		always @(posedge clk) O51_N2_S2 <=     O51_N4_S1  +  O51_N6_S1 ;
 logic signed [21:0] O51_N4_S2;		always @(posedge clk) O51_N4_S2 <=     O51_N8_S1  +  O51_N10_S1 ;
 logic signed [21:0] O51_N6_S2;		always @(posedge clk) O51_N6_S2 <=     O51_N12_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O51_N0_S3;		always @(posedge clk) O51_N0_S3 <=     O51_N0_S2  +  O51_N2_S2 ;
 logic signed [22:0] O51_N2_S3;		always @(posedge clk) O51_N2_S3 <=     O51_N4_S2  +  O51_N6_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O51_N0_S4;		always @(posedge clk) O51_N0_S4 <=     O51_N0_S3  +  O51_N2_S3 ;
 assign conv_mac_51 = O51_N0_S4;

logic signed [31:0] conv_mac_52;
logic signed [63:0] chainout_0_O52; 
logic signed [63:0] O52_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O52(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd1),.bx(input_fmap_1[7:0]),.by(-9'sd1),.cx(input_fmap_2[7:0]),.cy( 9'sd1),.dx(input_fmap_3[7:0]),.dy( 9'sd3),.chainin(63'd0),.result(O52_N0_S1),.chainout(chainout_0_O52));
logic signed [63:0] chainout_2_O52; 
logic signed [63:0] O52_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O52(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_4[7:0]),.ay(-9'sd3),.bx(input_fmap_5[7:0]),.by(-9'sd1),.cx(input_fmap_6[7:0]),.cy(-9'sd1),.dx(input_fmap_7[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O52_N2_S1),.chainout(chainout_2_O52));
logic signed [63:0] chainout_4_O52; 
logic signed [63:0] O52_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O52(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_8[7:0]),.ay(-9'sd1),.bx(input_fmap_9[7:0]),.by(-9'sd1),.cx(input_fmap_10[7:0]),.cy(-9'sd2),.dx(input_fmap_11[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O52_N4_S1),.chainout(chainout_4_O52));
logic signed [63:0] chainout_6_O52; 
logic signed [63:0] O52_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O52(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_13[7:0]),.ay( 9'sd1),.bx(input_fmap_14[7:0]),.by( 9'sd1),.cx(input_fmap_15[7:0]),.cy(-9'sd2),.dx(input_fmap_16[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O52_N6_S1),.chainout(chainout_6_O52));
logic signed [63:0] chainout_8_O52; 
logic signed [63:0] O52_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O52(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_20[7:0]),.ay( 9'sd3),.bx(input_fmap_21[7:0]),.by(-9'sd1),.cx(input_fmap_23[7:0]),.cy( 9'sd1),.dx(input_fmap_24[7:0]),.dy( 9'sd3),.chainin(63'd0),.result(O52_N8_S1),.chainout(chainout_8_O52));
logic signed [63:0] chainout_10_O52; 
logic signed [63:0] O52_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O52(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_25[7:0]),.ay( 9'sd2),.bx(input_fmap_26[7:0]),.by( 9'sd2),.cx(input_fmap_27[7:0]),.cy( 9'sd2),.dx(input_fmap_34[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O52_N10_S1),.chainout(chainout_10_O52));
logic signed [63:0] chainout_12_O52; 
logic signed [63:0] O52_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O52(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_35[7:0]),.ay(-9'sd1),.bx(input_fmap_37[7:0]),.by(-9'sd4),.cx(input_fmap_38[7:0]),.cy( 9'sd1),.dx(input_fmap_40[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O52_N12_S1),.chainout(chainout_12_O52));
logic signed [63:0] chainout_14_O52; 
logic signed [63:0] O52_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O52(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_41[7:0]),.ay(-9'sd1),.bx(input_fmap_42[7:0]),.by(-9'sd1),.cx(input_fmap_43[7:0]),.cy(-9'sd1),.dx(input_fmap_45[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O52_N14_S1),.chainout(chainout_14_O52));
logic signed [63:0] chainout_16_O52; 
logic signed [63:0] O52_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O52(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_46[7:0]),.ay( 9'sd1),.bx(input_fmap_50[7:0]),.by( 9'sd1),.cx(input_fmap_51[7:0]),.cy(-9'sd4),.dx(input_fmap_52[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O52_N16_S1),.chainout(chainout_16_O52));
logic signed [63:0] chainout_18_O52; 
logic signed [63:0] O52_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O52(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_53[7:0]),.ay(-9'sd1),.bx(input_fmap_54[7:0]),.by(-9'sd1),.cx(input_fmap_55[7:0]),.cy( 9'sd3),.dx(input_fmap_56[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O52_N18_S1),.chainout(chainout_18_O52));
logic signed [63:0] chainout_20_O52; 
logic signed [63:0] O52_N20_S1; 
 int_sop_4_wrapper int_sop_4_inst_20_O52(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_57[7:0]),.ay( 9'sd4),.bx(input_fmap_58[7:0]),.by( 9'sd2),.cx(input_fmap_59[7:0]),.cy( 9'sd2),.dx(input_fmap_61[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O52_N20_S1),.chainout(chainout_20_O52));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O52_N0_S2;		always @(posedge clk) O52_N0_S2 <=     O52_N0_S1  +  O52_N2_S1 ;
 logic signed [21:0] O52_N2_S2;		always @(posedge clk) O52_N2_S2 <=     O52_N4_S1  +  O52_N6_S1 ;
 logic signed [21:0] O52_N4_S2;		always @(posedge clk) O52_N4_S2 <=     O52_N8_S1  +  O52_N10_S1 ;
 logic signed [21:0] O52_N6_S2;		always @(posedge clk) O52_N6_S2 <=     O52_N12_S1  +  O52_N14_S1 ;
 logic signed [21:0] O52_N8_S2;		always @(posedge clk) O52_N8_S2 <=     O52_N16_S1  +  O52_N18_S1 ;
 logic signed [21:0] O52_N10_S2;		always @(posedge clk) O52_N10_S2 <=     O52_N20_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O52_N0_S3;		always @(posedge clk) O52_N0_S3 <=     O52_N0_S2  +  O52_N2_S2 ;
 logic signed [22:0] O52_N2_S3;		always @(posedge clk) O52_N2_S3 <=     O52_N4_S2  +  O52_N6_S2 ;
 logic signed [22:0] O52_N4_S3;		always @(posedge clk) O52_N4_S3 <=     O52_N8_S2  +  O52_N10_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O52_N0_S4;		always @(posedge clk) O52_N0_S4 <=     O52_N0_S3  +  O52_N2_S3 ;
 logic signed [23:0] O52_N2_S4;		always @(posedge clk) O52_N2_S4 <=     O52_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O52_N0_S5;		always @(posedge clk) O52_N0_S5 <=     O52_N0_S4  +  O52_N2_S4 ;
 assign conv_mac_52 = O52_N0_S5;

logic signed [31:0] conv_mac_53;
logic signed [63:0] chainout_0_O53; 
logic signed [63:0] O53_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O53(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd1),.bx(input_fmap_1[7:0]),.by(-9'sd2),.cx(input_fmap_2[7:0]),.cy( 9'sd1),.dx(input_fmap_3[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O53_N0_S1),.chainout(chainout_0_O53));
logic signed [63:0] chainout_2_O53; 
logic signed [63:0] O53_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O53(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_4[7:0]),.ay(-9'sd2),.bx(input_fmap_6[7:0]),.by( 9'sd1),.cx(input_fmap_8[7:0]),.cy( 9'sd2),.dx(input_fmap_9[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O53_N2_S1),.chainout(chainout_2_O53));
logic signed [63:0] chainout_4_O53; 
logic signed [63:0] O53_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O53(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_10[7:0]),.ay(-9'sd1),.bx(input_fmap_12[7:0]),.by(-9'sd2),.cx(input_fmap_13[7:0]),.cy( 9'sd2),.dx(input_fmap_16[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O53_N4_S1),.chainout(chainout_4_O53));
logic signed [63:0] chainout_6_O53; 
logic signed [63:0] O53_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O53(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_17[7:0]),.ay( 9'sd3),.bx(input_fmap_19[7:0]),.by( 9'sd2),.cx(input_fmap_23[7:0]),.cy(-9'sd1),.dx(input_fmap_24[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O53_N6_S1),.chainout(chainout_6_O53));
logic signed [63:0] chainout_8_O53; 
logic signed [63:0] O53_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O53(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_25[7:0]),.ay( 9'sd1),.bx(input_fmap_26[7:0]),.by( 9'sd1),.cx(input_fmap_27[7:0]),.cy(-9'sd1),.dx(input_fmap_28[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O53_N8_S1),.chainout(chainout_8_O53));
logic signed [63:0] chainout_10_O53; 
logic signed [63:0] O53_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O53(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_29[7:0]),.ay( 9'sd1),.bx(input_fmap_31[7:0]),.by(-9'sd1),.cx(input_fmap_32[7:0]),.cy( 9'sd2),.dx(input_fmap_34[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O53_N10_S1),.chainout(chainout_10_O53));
logic signed [63:0] chainout_12_O53; 
logic signed [63:0] O53_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O53(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_35[7:0]),.ay( 9'sd1),.bx(input_fmap_36[7:0]),.by(-9'sd1),.cx(input_fmap_37[7:0]),.cy( 9'sd1),.dx(input_fmap_39[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O53_N12_S1),.chainout(chainout_12_O53));
logic signed [63:0] chainout_14_O53; 
logic signed [63:0] O53_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O53(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_40[7:0]),.ay( 9'sd1),.bx(input_fmap_41[7:0]),.by(-9'sd1),.cx(input_fmap_43[7:0]),.cy(-9'sd2),.dx(input_fmap_44[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O53_N14_S1),.chainout(chainout_14_O53));
logic signed [63:0] chainout_16_O53; 
logic signed [63:0] O53_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O53(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_46[7:0]),.ay( 9'sd1),.bx(input_fmap_49[7:0]),.by( 9'sd2),.cx(input_fmap_50[7:0]),.cy(-9'sd3),.dx(input_fmap_51[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O53_N16_S1),.chainout(chainout_16_O53));
logic signed [63:0] chainout_18_O53; 
logic signed [63:0] O53_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O53(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_54[7:0]),.ay(-9'sd1),.bx(input_fmap_55[7:0]),.by( 9'sd1),.cx(input_fmap_56[7:0]),.cy( 9'sd1),.dx(input_fmap_60[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O53_N18_S1),.chainout(chainout_18_O53));
logic signed [63:0] chainout_20_O53; 
logic signed [63:0] O53_N20_S1; 
 int_sop_4_wrapper int_sop_4_inst_20_O53(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_61[7:0]),.ay(-9'sd2),.bx(input_fmap_63[7:0]),.by( 9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O53_N20_S1),.chainout(chainout_20_O53));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O53_N0_S2;		always @(posedge clk) O53_N0_S2 <=     O53_N0_S1  +  O53_N2_S1 ;
 logic signed [21:0] O53_N2_S2;		always @(posedge clk) O53_N2_S2 <=     O53_N4_S1  +  O53_N6_S1 ;
 logic signed [21:0] O53_N4_S2;		always @(posedge clk) O53_N4_S2 <=     O53_N8_S1  +  O53_N10_S1 ;
 logic signed [21:0] O53_N6_S2;		always @(posedge clk) O53_N6_S2 <=     O53_N12_S1  +  O53_N14_S1 ;
 logic signed [21:0] O53_N8_S2;		always @(posedge clk) O53_N8_S2 <=     O53_N16_S1  +  O53_N18_S1 ;
 logic signed [21:0] O53_N10_S2;		always @(posedge clk) O53_N10_S2 <=     O53_N20_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O53_N0_S3;		always @(posedge clk) O53_N0_S3 <=     O53_N0_S2  +  O53_N2_S2 ;
 logic signed [22:0] O53_N2_S3;		always @(posedge clk) O53_N2_S3 <=     O53_N4_S2  +  O53_N6_S2 ;
 logic signed [22:0] O53_N4_S3;		always @(posedge clk) O53_N4_S3 <=     O53_N8_S2  +  O53_N10_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O53_N0_S4;		always @(posedge clk) O53_N0_S4 <=     O53_N0_S3  +  O53_N2_S3 ;
 logic signed [23:0] O53_N2_S4;		always @(posedge clk) O53_N2_S4 <=     O53_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O53_N0_S5;		always @(posedge clk) O53_N0_S5 <=     O53_N0_S4  +  O53_N2_S4 ;
 assign conv_mac_53 = O53_N0_S5;

logic signed [31:0] conv_mac_54;
logic signed [63:0] chainout_0_O54; 
logic signed [63:0] O54_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O54(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd1),.bx(input_fmap_2[7:0]),.by( 9'sd2),.cx(input_fmap_3[7:0]),.cy( 9'sd1),.dx(input_fmap_4[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O54_N0_S1),.chainout(chainout_0_O54));
logic signed [63:0] chainout_2_O54; 
logic signed [63:0] O54_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O54(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_10[7:0]),.ay(-9'sd1),.bx(input_fmap_11[7:0]),.by(-9'sd1),.cx(input_fmap_13[7:0]),.cy( 9'sd1),.dx(input_fmap_14[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O54_N2_S1),.chainout(chainout_2_O54));
logic signed [63:0] chainout_4_O54; 
logic signed [63:0] O54_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O54(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_15[7:0]),.ay( 9'sd1),.bx(input_fmap_16[7:0]),.by(-9'sd1),.cx(input_fmap_17[7:0]),.cy(-9'sd1),.dx(input_fmap_18[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O54_N4_S1),.chainout(chainout_4_O54));
logic signed [63:0] chainout_6_O54; 
logic signed [63:0] O54_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O54(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_19[7:0]),.ay( 9'sd2),.bx(input_fmap_20[7:0]),.by( 9'sd1),.cx(input_fmap_21[7:0]),.cy( 9'sd1),.dx(input_fmap_22[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O54_N6_S1),.chainout(chainout_6_O54));
logic signed [63:0] chainout_8_O54; 
logic signed [63:0] O54_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O54(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_28[7:0]),.ay( 9'sd1),.bx(input_fmap_29[7:0]),.by( 9'sd1),.cx(input_fmap_33[7:0]),.cy( 9'sd1),.dx(input_fmap_34[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O54_N8_S1),.chainout(chainout_8_O54));
logic signed [63:0] chainout_10_O54; 
logic signed [63:0] O54_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O54(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_37[7:0]),.ay( 9'sd1),.bx(input_fmap_38[7:0]),.by( 9'sd1),.cx(input_fmap_41[7:0]),.cy( 9'sd1),.dx(input_fmap_42[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O54_N10_S1),.chainout(chainout_10_O54));
logic signed [63:0] chainout_12_O54; 
logic signed [63:0] O54_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O54(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_43[7:0]),.ay( 9'sd2),.bx(input_fmap_44[7:0]),.by(-9'sd1),.cx(input_fmap_46[7:0]),.cy( 9'sd1),.dx(input_fmap_47[7:0]),.dy(-9'sd3),.chainin(63'd0),.result(O54_N12_S1),.chainout(chainout_12_O54));
logic signed [63:0] chainout_14_O54; 
logic signed [63:0] O54_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O54(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_51[7:0]),.ay( 9'sd1),.bx(input_fmap_52[7:0]),.by( 9'sd1),.cx(input_fmap_53[7:0]),.cy( 9'sd1),.dx(input_fmap_55[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O54_N14_S1),.chainout(chainout_14_O54));
logic signed [63:0] chainout_16_O54; 
logic signed [63:0] O54_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O54(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_57[7:0]),.ay( 9'sd1),.bx(input_fmap_58[7:0]),.by( 9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O54_N16_S1),.chainout(chainout_16_O54));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O54_N0_S2;		always @(posedge clk) O54_N0_S2 <=     O54_N0_S1  +  O54_N2_S1 ;
 logic signed [21:0] O54_N2_S2;		always @(posedge clk) O54_N2_S2 <=     O54_N4_S1  +  O54_N6_S1 ;
 logic signed [21:0] O54_N4_S2;		always @(posedge clk) O54_N4_S2 <=     O54_N8_S1  +  O54_N10_S1 ;
 logic signed [21:0] O54_N6_S2;		always @(posedge clk) O54_N6_S2 <=     O54_N12_S1  +  O54_N14_S1 ;
 logic signed [21:0] O54_N8_S2;		always @(posedge clk) O54_N8_S2 <=     O54_N16_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O54_N0_S3;		always @(posedge clk) O54_N0_S3 <=     O54_N0_S2  +  O54_N2_S2 ;
 logic signed [22:0] O54_N2_S3;		always @(posedge clk) O54_N2_S3 <=     O54_N4_S2  +  O54_N6_S2 ;
 logic signed [22:0] O54_N4_S3;		always @(posedge clk) O54_N4_S3 <=     O54_N8_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O54_N0_S4;		always @(posedge clk) O54_N0_S4 <=     O54_N0_S3  +  O54_N2_S3 ;
 logic signed [23:0] O54_N2_S4;		always @(posedge clk) O54_N2_S4 <=     O54_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O54_N0_S5;		always @(posedge clk) O54_N0_S5 <=     O54_N0_S4  +  O54_N2_S4 ;
 assign conv_mac_54 = O54_N0_S5;

logic signed [31:0] conv_mac_55;
logic signed [63:0] chainout_0_O55; 
logic signed [63:0] O55_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O55(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd1),.bx(input_fmap_2[7:0]),.by(-9'sd2),.cx(input_fmap_3[7:0]),.cy(-9'sd1),.dx(input_fmap_5[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O55_N0_S1),.chainout(chainout_0_O55));
logic signed [63:0] chainout_2_O55; 
logic signed [63:0] O55_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O55(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_6[7:0]),.ay( 9'sd1),.bx(input_fmap_7[7:0]),.by(-9'sd1),.cx(input_fmap_8[7:0]),.cy( 9'sd2),.dx(input_fmap_14[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O55_N2_S1),.chainout(chainout_2_O55));
logic signed [63:0] chainout_4_O55; 
logic signed [63:0] O55_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O55(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_15[7:0]),.ay(-9'sd1),.bx(input_fmap_16[7:0]),.by( 9'sd1),.cx(input_fmap_17[7:0]),.cy( 9'sd1),.dx(input_fmap_18[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O55_N4_S1),.chainout(chainout_4_O55));
logic signed [63:0] chainout_6_O55; 
logic signed [63:0] O55_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O55(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_20[7:0]),.ay(-9'sd1),.bx(input_fmap_21[7:0]),.by( 9'sd1),.cx(input_fmap_24[7:0]),.cy(-9'sd1),.dx(input_fmap_25[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O55_N6_S1),.chainout(chainout_6_O55));
logic signed [63:0] chainout_8_O55; 
logic signed [63:0] O55_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O55(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_26[7:0]),.ay(-9'sd1),.bx(input_fmap_30[7:0]),.by(-9'sd1),.cx(input_fmap_37[7:0]),.cy( 9'sd1),.dx(input_fmap_39[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O55_N8_S1),.chainout(chainout_8_O55));
logic signed [63:0] chainout_10_O55; 
logic signed [63:0] O55_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O55(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_40[7:0]),.ay( 9'sd1),.bx(input_fmap_43[7:0]),.by(-9'sd1),.cx(input_fmap_45[7:0]),.cy( 9'sd1),.dx(input_fmap_48[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O55_N10_S1),.chainout(chainout_10_O55));
logic signed [63:0] chainout_12_O55; 
logic signed [63:0] O55_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O55(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_50[7:0]),.ay(-9'sd1),.bx(input_fmap_52[7:0]),.by( 9'sd2),.cx(input_fmap_57[7:0]),.cy( 9'sd1),.dx(input_fmap_63[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O55_N12_S1),.chainout(chainout_12_O55));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O55_N0_S2;		always @(posedge clk) O55_N0_S2 <=     O55_N0_S1  +  O55_N2_S1 ;
 logic signed [21:0] O55_N2_S2;		always @(posedge clk) O55_N2_S2 <=     O55_N4_S1  +  O55_N6_S1 ;
 logic signed [21:0] O55_N4_S2;		always @(posedge clk) O55_N4_S2 <=     O55_N8_S1  +  O55_N10_S1 ;
 logic signed [21:0] O55_N6_S2;		always @(posedge clk) O55_N6_S2 <=     O55_N12_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O55_N0_S3;		always @(posedge clk) O55_N0_S3 <=     O55_N0_S2  +  O55_N2_S2 ;
 logic signed [22:0] O55_N2_S3;		always @(posedge clk) O55_N2_S3 <=     O55_N4_S2  +  O55_N6_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O55_N0_S4;		always @(posedge clk) O55_N0_S4 <=     O55_N0_S3  +  O55_N2_S3 ;
 assign conv_mac_55 = O55_N0_S4;

logic signed [31:0] conv_mac_56;
logic signed [63:0] chainout_0_O56; 
logic signed [63:0] O56_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O56(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd1),.bx(input_fmap_7[7:0]),.by(-9'sd1),.cx(input_fmap_8[7:0]),.cy(-9'sd1),.dx(input_fmap_10[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O56_N0_S1),.chainout(chainout_0_O56));
logic signed [63:0] chainout_2_O56; 
logic signed [63:0] O56_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O56(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_13[7:0]),.ay( 9'sd2),.bx(input_fmap_14[7:0]),.by( 9'sd1),.cx(input_fmap_17[7:0]),.cy(-9'sd1),.dx(input_fmap_18[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O56_N2_S1),.chainout(chainout_2_O56));
logic signed [63:0] chainout_4_O56; 
logic signed [63:0] O56_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O56(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_19[7:0]),.ay(-9'sd1),.bx(input_fmap_21[7:0]),.by( 9'sd2),.cx(input_fmap_22[7:0]),.cy(-9'sd2),.dx(input_fmap_23[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O56_N4_S1),.chainout(chainout_4_O56));
logic signed [63:0] chainout_6_O56; 
logic signed [63:0] O56_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O56(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_24[7:0]),.ay( 9'sd1),.bx(input_fmap_25[7:0]),.by(-9'sd1),.cx(input_fmap_27[7:0]),.cy(-9'sd1),.dx(input_fmap_28[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O56_N6_S1),.chainout(chainout_6_O56));
logic signed [63:0] chainout_8_O56; 
logic signed [63:0] O56_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O56(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_30[7:0]),.ay( 9'sd1),.bx(input_fmap_31[7:0]),.by( 9'sd2),.cx(input_fmap_32[7:0]),.cy(-9'sd1),.dx(input_fmap_35[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O56_N8_S1),.chainout(chainout_8_O56));
logic signed [63:0] chainout_10_O56; 
logic signed [63:0] O56_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O56(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_36[7:0]),.ay( 9'sd1),.bx(input_fmap_37[7:0]),.by(-9'sd1),.cx(input_fmap_38[7:0]),.cy( 9'sd1),.dx(input_fmap_41[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O56_N10_S1),.chainout(chainout_10_O56));
logic signed [63:0] chainout_12_O56; 
logic signed [63:0] O56_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O56(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_43[7:0]),.ay(-9'sd1),.bx(input_fmap_46[7:0]),.by( 9'sd1),.cx(input_fmap_47[7:0]),.cy( 9'sd1),.dx(input_fmap_49[7:0]),.dy( 9'sd3),.chainin(63'd0),.result(O56_N12_S1),.chainout(chainout_12_O56));
logic signed [63:0] chainout_14_O56; 
logic signed [63:0] O56_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O56(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_51[7:0]),.ay(-9'sd1),.bx(input_fmap_52[7:0]),.by( 9'sd1),.cx(input_fmap_57[7:0]),.cy( 9'sd2),.dx(input_fmap_59[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O56_N14_S1),.chainout(chainout_14_O56));
logic signed [63:0] chainout_16_O56; 
logic signed [63:0] O56_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O56(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_62[7:0]),.ay( 9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O56_N16_S1),.chainout(chainout_16_O56));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O56_N0_S2;		always @(posedge clk) O56_N0_S2 <=     O56_N0_S1  +  O56_N2_S1 ;
 logic signed [21:0] O56_N2_S2;		always @(posedge clk) O56_N2_S2 <=     O56_N4_S1  +  O56_N6_S1 ;
 logic signed [21:0] O56_N4_S2;		always @(posedge clk) O56_N4_S2 <=     O56_N8_S1  +  O56_N10_S1 ;
 logic signed [21:0] O56_N6_S2;		always @(posedge clk) O56_N6_S2 <=     O56_N12_S1  +  O56_N14_S1 ;
 logic signed [21:0] O56_N8_S2;		always @(posedge clk) O56_N8_S2 <=     O56_N16_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O56_N0_S3;		always @(posedge clk) O56_N0_S3 <=     O56_N0_S2  +  O56_N2_S2 ;
 logic signed [22:0] O56_N2_S3;		always @(posedge clk) O56_N2_S3 <=     O56_N4_S2  +  O56_N6_S2 ;
 logic signed [22:0] O56_N4_S3;		always @(posedge clk) O56_N4_S3 <=     O56_N8_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O56_N0_S4;		always @(posedge clk) O56_N0_S4 <=     O56_N0_S3  +  O56_N2_S3 ;
 logic signed [23:0] O56_N2_S4;		always @(posedge clk) O56_N2_S4 <=     O56_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O56_N0_S5;		always @(posedge clk) O56_N0_S5 <=     O56_N0_S4  +  O56_N2_S4 ;
 assign conv_mac_56 = O56_N0_S5;

logic signed [31:0] conv_mac_57;
logic signed [63:0] chainout_0_O57; 
logic signed [63:0] O57_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O57(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_6[7:0]),.ay( 9'sd1),.bx(input_fmap_8[7:0]),.by(-9'sd1),.cx(input_fmap_20[7:0]),.cy( 9'sd2),.dx(input_fmap_28[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O57_N0_S1),.chainout(chainout_0_O57));
logic signed [63:0] chainout_2_O57; 
logic signed [63:0] O57_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O57(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_30[7:0]),.ay( 9'sd1),.bx(input_fmap_46[7:0]),.by(-9'sd1),.cx(input_fmap_48[7:0]),.cy( 9'sd1),.dx(input_fmap_56[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O57_N2_S1),.chainout(chainout_2_O57));
logic signed [63:0] chainout_4_O57; 
logic signed [63:0] O57_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O57(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_61[7:0]),.ay(-9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O57_N4_S1),.chainout(chainout_4_O57));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O57_N0_S2;		always @(posedge clk) O57_N0_S2 <=     O57_N0_S1  +  O57_N2_S1 ;
 logic signed [21:0] O57_N2_S2;		always @(posedge clk) O57_N2_S2 <=     O57_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O57_N0_S3;		always @(posedge clk) O57_N0_S3 <=     O57_N0_S2  +  O57_N2_S2 ;
 assign conv_mac_57 = O57_N0_S3;

logic signed [31:0] conv_mac_58;
logic signed [63:0] chainout_0_O58; 
logic signed [63:0] O58_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O58(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd1),.bx(input_fmap_1[7:0]),.by( 9'sd2),.cx(input_fmap_6[7:0]),.cy( 9'sd1),.dx(input_fmap_7[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O58_N0_S1),.chainout(chainout_0_O58));
logic signed [63:0] chainout_2_O58; 
logic signed [63:0] O58_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O58(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_9[7:0]),.ay( 9'sd1),.bx(input_fmap_10[7:0]),.by(-9'sd1),.cx(input_fmap_11[7:0]),.cy( 9'sd2),.dx(input_fmap_13[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O58_N2_S1),.chainout(chainout_2_O58));
logic signed [63:0] chainout_4_O58; 
logic signed [63:0] O58_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O58(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_14[7:0]),.ay( 9'sd1),.bx(input_fmap_16[7:0]),.by( 9'sd2),.cx(input_fmap_17[7:0]),.cy(-9'sd1),.dx(input_fmap_18[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O58_N4_S1),.chainout(chainout_4_O58));
logic signed [63:0] chainout_6_O58; 
logic signed [63:0] O58_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O58(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_19[7:0]),.ay(-9'sd1),.bx(input_fmap_21[7:0]),.by(-9'sd1),.cx(input_fmap_27[7:0]),.cy(-9'sd1),.dx(input_fmap_29[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O58_N6_S1),.chainout(chainout_6_O58));
logic signed [63:0] chainout_8_O58; 
logic signed [63:0] O58_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O58(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_32[7:0]),.ay( 9'sd1),.bx(input_fmap_34[7:0]),.by(-9'sd1),.cx(input_fmap_35[7:0]),.cy(-9'sd1),.dx(input_fmap_38[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O58_N8_S1),.chainout(chainout_8_O58));
logic signed [63:0] chainout_10_O58; 
logic signed [63:0] O58_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O58(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_41[7:0]),.ay( 9'sd1),.bx(input_fmap_42[7:0]),.by(-9'sd1),.cx(input_fmap_43[7:0]),.cy(-9'sd1),.dx(input_fmap_44[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O58_N10_S1),.chainout(chainout_10_O58));
logic signed [63:0] chainout_12_O58; 
logic signed [63:0] O58_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O58(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_46[7:0]),.ay(-9'sd1),.bx(input_fmap_47[7:0]),.by(-9'sd1),.cx(input_fmap_48[7:0]),.cy(-9'sd1),.dx(input_fmap_50[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O58_N12_S1),.chainout(chainout_12_O58));
logic signed [63:0] chainout_14_O58; 
logic signed [63:0] O58_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O58(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_51[7:0]),.ay( 9'sd1),.bx(input_fmap_52[7:0]),.by( 9'sd1),.cx(input_fmap_54[7:0]),.cy( 9'sd1),.dx(input_fmap_56[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O58_N14_S1),.chainout(chainout_14_O58));
logic signed [63:0] chainout_16_O58; 
logic signed [63:0] O58_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O58(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_57[7:0]),.ay(-9'sd1),.bx(input_fmap_59[7:0]),.by( 9'sd1),.cx(input_fmap_60[7:0]),.cy( 9'sd1),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O58_N16_S1),.chainout(chainout_16_O58));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O58_N0_S2;		always @(posedge clk) O58_N0_S2 <=     O58_N0_S1  +  O58_N2_S1 ;
 logic signed [21:0] O58_N2_S2;		always @(posedge clk) O58_N2_S2 <=     O58_N4_S1  +  O58_N6_S1 ;
 logic signed [21:0] O58_N4_S2;		always @(posedge clk) O58_N4_S2 <=     O58_N8_S1  +  O58_N10_S1 ;
 logic signed [21:0] O58_N6_S2;		always @(posedge clk) O58_N6_S2 <=     O58_N12_S1  +  O58_N14_S1 ;
 logic signed [21:0] O58_N8_S2;		always @(posedge clk) O58_N8_S2 <=     O58_N16_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O58_N0_S3;		always @(posedge clk) O58_N0_S3 <=     O58_N0_S2  +  O58_N2_S2 ;
 logic signed [22:0] O58_N2_S3;		always @(posedge clk) O58_N2_S3 <=     O58_N4_S2  +  O58_N6_S2 ;
 logic signed [22:0] O58_N4_S3;		always @(posedge clk) O58_N4_S3 <=     O58_N8_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O58_N0_S4;		always @(posedge clk) O58_N0_S4 <=     O58_N0_S3  +  O58_N2_S3 ;
 logic signed [23:0] O58_N2_S4;		always @(posedge clk) O58_N2_S4 <=     O58_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O58_N0_S5;		always @(posedge clk) O58_N0_S5 <=     O58_N0_S4  +  O58_N2_S4 ;
 assign conv_mac_58 = O58_N0_S5;

logic signed [31:0] conv_mac_59;
logic signed [63:0] chainout_0_O59; 
logic signed [63:0] O59_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O59(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd1),.bx(input_fmap_4[7:0]),.by( 9'sd1),.cx(input_fmap_7[7:0]),.cy(-9'sd1),.dx(input_fmap_18[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O59_N0_S1),.chainout(chainout_0_O59));
logic signed [63:0] chainout_2_O59; 
logic signed [63:0] O59_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O59(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_23[7:0]),.ay( 9'sd1),.bx(input_fmap_27[7:0]),.by(-9'sd1),.cx(input_fmap_28[7:0]),.cy(-9'sd1),.dx(input_fmap_31[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O59_N2_S1),.chainout(chainout_2_O59));
logic signed [63:0] chainout_4_O59; 
logic signed [63:0] O59_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O59(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_35[7:0]),.ay(-9'sd1),.bx(input_fmap_43[7:0]),.by(-9'sd1),.cx(input_fmap_46[7:0]),.cy( 9'sd1),.dx(input_fmap_48[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O59_N4_S1),.chainout(chainout_4_O59));
logic signed [63:0] chainout_6_O59; 
logic signed [63:0] O59_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O59(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_51[7:0]),.ay( 9'sd1),.bx(input_fmap_56[7:0]),.by( 9'sd1),.cx(input_fmap_61[7:0]),.cy(-9'sd2),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O59_N6_S1),.chainout(chainout_6_O59));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O59_N0_S2;		always @(posedge clk) O59_N0_S2 <=     O59_N0_S1  +  O59_N2_S1 ;
 logic signed [21:0] O59_N2_S2;		always @(posedge clk) O59_N2_S2 <=     O59_N4_S1  +  O59_N6_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O59_N0_S3;		always @(posedge clk) O59_N0_S3 <=     O59_N0_S2  +  O59_N2_S2 ;
 assign conv_mac_59 = O59_N0_S3;

logic signed [31:0] conv_mac_60;
logic signed [63:0] chainout_0_O60; 
logic signed [63:0] O60_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O60(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd1),.bx(input_fmap_1[7:0]),.by( 9'sd1),.cx(input_fmap_2[7:0]),.cy(-9'sd2),.dx(input_fmap_4[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O60_N0_S1),.chainout(chainout_0_O60));
logic signed [63:0] chainout_2_O60; 
logic signed [63:0] O60_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O60(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_5[7:0]),.ay( 9'sd1),.bx(input_fmap_9[7:0]),.by(-9'sd1),.cx(input_fmap_10[7:0]),.cy( 9'sd1),.dx(input_fmap_12[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O60_N2_S1),.chainout(chainout_2_O60));
logic signed [63:0] chainout_4_O60; 
logic signed [63:0] O60_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O60(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_14[7:0]),.ay(-9'sd2),.bx(input_fmap_15[7:0]),.by(-9'sd1),.cx(input_fmap_17[7:0]),.cy(-9'sd2),.dx(input_fmap_18[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O60_N4_S1),.chainout(chainout_4_O60));
logic signed [63:0] chainout_6_O60; 
logic signed [63:0] O60_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O60(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_19[7:0]),.ay(-9'sd2),.bx(input_fmap_20[7:0]),.by(-9'sd1),.cx(input_fmap_21[7:0]),.cy( 9'sd1),.dx(input_fmap_23[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O60_N6_S1),.chainout(chainout_6_O60));
logic signed [63:0] chainout_8_O60; 
logic signed [63:0] O60_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O60(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_24[7:0]),.ay(-9'sd1),.bx(input_fmap_25[7:0]),.by(-9'sd1),.cx(input_fmap_27[7:0]),.cy(-9'sd1),.dx(input_fmap_28[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O60_N8_S1),.chainout(chainout_8_O60));
logic signed [63:0] chainout_10_O60; 
logic signed [63:0] O60_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O60(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_31[7:0]),.ay( 9'sd1),.bx(input_fmap_32[7:0]),.by( 9'sd2),.cx(input_fmap_34[7:0]),.cy( 9'sd1),.dx(input_fmap_35[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O60_N10_S1),.chainout(chainout_10_O60));
logic signed [63:0] chainout_12_O60; 
logic signed [63:0] O60_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O60(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_36[7:0]),.ay( 9'sd2),.bx(input_fmap_42[7:0]),.by(-9'sd1),.cx(input_fmap_43[7:0]),.cy(-9'sd1),.dx(input_fmap_44[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O60_N12_S1),.chainout(chainout_12_O60));
logic signed [63:0] chainout_14_O60; 
logic signed [63:0] O60_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O60(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_45[7:0]),.ay(-9'sd1),.bx(input_fmap_46[7:0]),.by( 9'sd2),.cx(input_fmap_49[7:0]),.cy( 9'sd1),.dx(input_fmap_50[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O60_N14_S1),.chainout(chainout_14_O60));
logic signed [63:0] chainout_16_O60; 
logic signed [63:0] O60_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O60(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_52[7:0]),.ay(-9'sd1),.bx(input_fmap_53[7:0]),.by( 9'sd1),.cx(input_fmap_56[7:0]),.cy( 9'sd1),.dx(input_fmap_58[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O60_N16_S1),.chainout(chainout_16_O60));
logic signed [63:0] chainout_18_O60; 
logic signed [63:0] O60_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O60(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_60[7:0]),.ay(-9'sd3),.bx(input_fmap_63[7:0]),.by(-9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O60_N18_S1),.chainout(chainout_18_O60));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O60_N0_S2;		always @(posedge clk) O60_N0_S2 <=     O60_N0_S1  +  O60_N2_S1 ;
 logic signed [21:0] O60_N2_S2;		always @(posedge clk) O60_N2_S2 <=     O60_N4_S1  +  O60_N6_S1 ;
 logic signed [21:0] O60_N4_S2;		always @(posedge clk) O60_N4_S2 <=     O60_N8_S1  +  O60_N10_S1 ;
 logic signed [21:0] O60_N6_S2;		always @(posedge clk) O60_N6_S2 <=     O60_N12_S1  +  O60_N14_S1 ;
 logic signed [21:0] O60_N8_S2;		always @(posedge clk) O60_N8_S2 <=     O60_N16_S1  +  O60_N18_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O60_N0_S3;		always @(posedge clk) O60_N0_S3 <=     O60_N0_S2  +  O60_N2_S2 ;
 logic signed [22:0] O60_N2_S3;		always @(posedge clk) O60_N2_S3 <=     O60_N4_S2  +  O60_N6_S2 ;
 logic signed [22:0] O60_N4_S3;		always @(posedge clk) O60_N4_S3 <=     O60_N8_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O60_N0_S4;		always @(posedge clk) O60_N0_S4 <=     O60_N0_S3  +  O60_N2_S3 ;
 logic signed [23:0] O60_N2_S4;		always @(posedge clk) O60_N2_S4 <=     O60_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O60_N0_S5;		always @(posedge clk) O60_N0_S5 <=     O60_N0_S4  +  O60_N2_S4 ;
 assign conv_mac_60 = O60_N0_S5;

logic signed [31:0] conv_mac_61;
logic signed [63:0] chainout_0_O61; 
logic signed [63:0] O61_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O61(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_3[7:0]),.ay(-9'sd1),.bx(input_fmap_5[7:0]),.by(-9'sd1),.cx(input_fmap_9[7:0]),.cy(-9'sd1),.dx(input_fmap_10[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O61_N0_S1),.chainout(chainout_0_O61));
logic signed [63:0] chainout_2_O61; 
logic signed [63:0] O61_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O61(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_11[7:0]),.ay( 9'sd1),.bx(input_fmap_15[7:0]),.by( 9'sd1),.cx(input_fmap_16[7:0]),.cy(-9'sd1),.dx(input_fmap_17[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O61_N2_S1),.chainout(chainout_2_O61));
logic signed [63:0] chainout_4_O61; 
logic signed [63:0] O61_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O61(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_19[7:0]),.ay(-9'sd2),.bx(input_fmap_21[7:0]),.by(-9'sd1),.cx(input_fmap_29[7:0]),.cy( 9'sd1),.dx(input_fmap_34[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O61_N4_S1),.chainout(chainout_4_O61));
logic signed [63:0] chainout_6_O61; 
logic signed [63:0] O61_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O61(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_38[7:0]),.ay(-9'sd1),.bx(input_fmap_39[7:0]),.by(-9'sd1),.cx(input_fmap_45[7:0]),.cy( 9'sd1),.dx(input_fmap_46[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O61_N6_S1),.chainout(chainout_6_O61));
logic signed [63:0] chainout_8_O61; 
logic signed [63:0] O61_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O61(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_47[7:0]),.ay( 9'sd2),.bx(input_fmap_48[7:0]),.by( 9'sd1),.cx(input_fmap_49[7:0]),.cy(-9'sd2),.dx(input_fmap_50[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O61_N8_S1),.chainout(chainout_8_O61));
logic signed [63:0] chainout_10_O61; 
logic signed [63:0] O61_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O61(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_51[7:0]),.ay(-9'sd2),.bx(input_fmap_52[7:0]),.by( 9'sd1),.cx(input_fmap_61[7:0]),.cy(-9'sd2),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O61_N10_S1),.chainout(chainout_10_O61));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O61_N0_S2;		always @(posedge clk) O61_N0_S2 <=     O61_N0_S1  +  O61_N2_S1 ;
 logic signed [21:0] O61_N2_S2;		always @(posedge clk) O61_N2_S2 <=     O61_N4_S1  +  O61_N6_S1 ;
 logic signed [21:0] O61_N4_S2;		always @(posedge clk) O61_N4_S2 <=     O61_N8_S1  +  O61_N10_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O61_N0_S3;		always @(posedge clk) O61_N0_S3 <=     O61_N0_S2  +  O61_N2_S2 ;
 logic signed [22:0] O61_N2_S3;		always @(posedge clk) O61_N2_S3 <=     O61_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O61_N0_S4;		always @(posedge clk) O61_N0_S4 <=     O61_N0_S3  +  O61_N2_S3 ;
 assign conv_mac_61 = O61_N0_S4;

logic signed [31:0] conv_mac_62;
logic signed [63:0] chainout_0_O62; 
logic signed [63:0] O62_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O62(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd1),.bx(input_fmap_1[7:0]),.by( 9'sd2),.cx(input_fmap_2[7:0]),.cy( 9'sd1),.dx(input_fmap_4[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O62_N0_S1),.chainout(chainout_0_O62));
logic signed [63:0] chainout_2_O62; 
logic signed [63:0] O62_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O62(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_5[7:0]),.ay(-9'sd1),.bx(input_fmap_6[7:0]),.by(-9'sd1),.cx(input_fmap_7[7:0]),.cy(-9'sd2),.dx(input_fmap_8[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O62_N2_S1),.chainout(chainout_2_O62));
logic signed [63:0] chainout_4_O62; 
logic signed [63:0] O62_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O62(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_10[7:0]),.ay(-9'sd3),.bx(input_fmap_11[7:0]),.by(-9'sd2),.cx(input_fmap_12[7:0]),.cy( 9'sd4),.dx(input_fmap_13[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O62_N4_S1),.chainout(chainout_4_O62));
logic signed [63:0] chainout_6_O62; 
logic signed [63:0] O62_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O62(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_16[7:0]),.ay( 9'sd1),.bx(input_fmap_17[7:0]),.by(-9'sd1),.cx(input_fmap_18[7:0]),.cy(-9'sd2),.dx(input_fmap_19[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O62_N6_S1),.chainout(chainout_6_O62));
logic signed [63:0] chainout_8_O62; 
logic signed [63:0] O62_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O62(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_21[7:0]),.ay( 9'sd2),.bx(input_fmap_22[7:0]),.by(-9'sd1),.cx(input_fmap_25[7:0]),.cy( 9'sd2),.dx(input_fmap_27[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O62_N8_S1),.chainout(chainout_8_O62));
logic signed [63:0] chainout_10_O62; 
logic signed [63:0] O62_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O62(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_28[7:0]),.ay(-9'sd1),.bx(input_fmap_29[7:0]),.by( 9'sd2),.cx(input_fmap_30[7:0]),.cy( 9'sd2),.dx(input_fmap_31[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O62_N10_S1),.chainout(chainout_10_O62));
logic signed [63:0] chainout_12_O62; 
logic signed [63:0] O62_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O62(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_32[7:0]),.ay(-9'sd1),.bx(input_fmap_33[7:0]),.by(-9'sd3),.cx(input_fmap_35[7:0]),.cy(-9'sd3),.dx(input_fmap_36[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O62_N12_S1),.chainout(chainout_12_O62));
logic signed [63:0] chainout_14_O62; 
logic signed [63:0] O62_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O62(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_37[7:0]),.ay( 9'sd2),.bx(input_fmap_38[7:0]),.by( 9'sd2),.cx(input_fmap_39[7:0]),.cy( 9'sd3),.dx(input_fmap_40[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O62_N14_S1),.chainout(chainout_14_O62));
logic signed [63:0] chainout_16_O62; 
logic signed [63:0] O62_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O62(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_41[7:0]),.ay(-9'sd1),.bx(input_fmap_42[7:0]),.by(-9'sd1),.cx(input_fmap_43[7:0]),.cy( 9'sd1),.dx(input_fmap_44[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O62_N16_S1),.chainout(chainout_16_O62));
logic signed [63:0] chainout_18_O62; 
logic signed [63:0] O62_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O62(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_45[7:0]),.ay( 9'sd1),.bx(input_fmap_46[7:0]),.by( 9'sd1),.cx(input_fmap_47[7:0]),.cy(-9'sd1),.dx(input_fmap_48[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O62_N18_S1),.chainout(chainout_18_O62));
logic signed [63:0] chainout_20_O62; 
logic signed [63:0] O62_N20_S1; 
 int_sop_4_wrapper int_sop_4_inst_20_O62(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_49[7:0]),.ay(-9'sd1),.bx(input_fmap_51[7:0]),.by(-9'sd3),.cx(input_fmap_52[7:0]),.cy(-9'sd1),.dx(input_fmap_53[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O62_N20_S1),.chainout(chainout_20_O62));
logic signed [63:0] chainout_22_O62; 
logic signed [63:0] O62_N22_S1; 
 int_sop_4_wrapper int_sop_4_inst_22_O62(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_54[7:0]),.ay(-9'sd2),.bx(input_fmap_55[7:0]),.by(-9'sd3),.cx(input_fmap_56[7:0]),.cy(-9'sd1),.dx(input_fmap_57[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O62_N22_S1),.chainout(chainout_22_O62));
logic signed [63:0] chainout_24_O62; 
logic signed [63:0] O62_N24_S1; 
 int_sop_4_wrapper int_sop_4_inst_24_O62(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_58[7:0]),.ay( 9'sd2),.bx(input_fmap_60[7:0]),.by( 9'sd1),.cx(input_fmap_62[7:0]),.cy(-9'sd1),.dx(input_fmap_63[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O62_N24_S1),.chainout(chainout_24_O62));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O62_N0_S2;		always @(posedge clk) O62_N0_S2 <=     O62_N0_S1  +  O62_N2_S1 ;
 logic signed [21:0] O62_N2_S2;		always @(posedge clk) O62_N2_S2 <=     O62_N4_S1  +  O62_N6_S1 ;
 logic signed [21:0] O62_N4_S2;		always @(posedge clk) O62_N4_S2 <=     O62_N8_S1  +  O62_N10_S1 ;
 logic signed [21:0] O62_N6_S2;		always @(posedge clk) O62_N6_S2 <=     O62_N12_S1  +  O62_N14_S1 ;
 logic signed [21:0] O62_N8_S2;		always @(posedge clk) O62_N8_S2 <=     O62_N16_S1  +  O62_N18_S1 ;
 logic signed [21:0] O62_N10_S2;		always @(posedge clk) O62_N10_S2 <=     O62_N20_S1  +  O62_N22_S1 ;
 logic signed [21:0] O62_N12_S2;		always @(posedge clk) O62_N12_S2 <=     O62_N24_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O62_N0_S3;		always @(posedge clk) O62_N0_S3 <=     O62_N0_S2  +  O62_N2_S2 ;
 logic signed [22:0] O62_N2_S3;		always @(posedge clk) O62_N2_S3 <=     O62_N4_S2  +  O62_N6_S2 ;
 logic signed [22:0] O62_N4_S3;		always @(posedge clk) O62_N4_S3 <=     O62_N8_S2  +  O62_N10_S2 ;
 logic signed [22:0] O62_N6_S3;		always @(posedge clk) O62_N6_S3 <=     O62_N12_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O62_N0_S4;		always @(posedge clk) O62_N0_S4 <=     O62_N0_S3  +  O62_N2_S3 ;
 logic signed [23:0] O62_N2_S4;		always @(posedge clk) O62_N2_S4 <=     O62_N4_S3  +  O62_N6_S3 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O62_N0_S5;		always @(posedge clk) O62_N0_S5 <=     O62_N0_S4  +  O62_N2_S4 ;
 assign conv_mac_62 = O62_N0_S5;

logic signed [31:0] conv_mac_63;
logic signed [63:0] chainout_0_O63; 
logic signed [63:0] O63_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O63(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay(-9'sd2),.bx(input_fmap_5[7:0]),.by(-9'sd2),.cx(input_fmap_7[7:0]),.cy( 9'sd2),.dx(input_fmap_8[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O63_N0_S1),.chainout(chainout_0_O63));
logic signed [63:0] chainout_2_O63; 
logic signed [63:0] O63_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O63(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_14[7:0]),.ay( 9'sd1),.bx(input_fmap_15[7:0]),.by( 9'sd3),.cx(input_fmap_16[7:0]),.cy(-9'sd1),.dx(input_fmap_18[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O63_N2_S1),.chainout(chainout_2_O63));
logic signed [63:0] chainout_4_O63; 
logic signed [63:0] O63_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O63(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_20[7:0]),.ay( 9'sd6),.bx(input_fmap_21[7:0]),.by(-9'sd1),.cx(input_fmap_22[7:0]),.cy( 9'sd1),.dx(input_fmap_23[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O63_N4_S1),.chainout(chainout_4_O63));
logic signed [63:0] chainout_6_O63; 
logic signed [63:0] O63_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O63(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_24[7:0]),.ay( 9'sd1),.bx(input_fmap_26[7:0]),.by(-9'sd1),.cx(input_fmap_27[7:0]),.cy( 9'sd1),.dx(input_fmap_30[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O63_N6_S1),.chainout(chainout_6_O63));
logic signed [63:0] chainout_8_O63; 
logic signed [63:0] O63_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O63(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_32[7:0]),.ay( 9'sd1),.bx(input_fmap_35[7:0]),.by(-9'sd1),.cx(input_fmap_37[7:0]),.cy( 9'sd5),.dx(input_fmap_40[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O63_N8_S1),.chainout(chainout_8_O63));
logic signed [63:0] chainout_10_O63; 
logic signed [63:0] O63_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O63(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_41[7:0]),.ay(-9'sd1),.bx(input_fmap_42[7:0]),.by( 9'sd1),.cx(input_fmap_43[7:0]),.cy( 9'sd3),.dx(input_fmap_45[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O63_N10_S1),.chainout(chainout_10_O63));
logic signed [63:0] chainout_12_O63; 
logic signed [63:0] O63_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O63(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_46[7:0]),.ay(-9'sd2),.bx(input_fmap_47[7:0]),.by( 9'sd1),.cx(input_fmap_48[7:0]),.cy(-9'sd1),.dx(input_fmap_49[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O63_N12_S1),.chainout(chainout_12_O63));
logic signed [63:0] chainout_14_O63; 
logic signed [63:0] O63_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O63(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_51[7:0]),.ay( 9'sd2),.bx(input_fmap_52[7:0]),.by(-9'sd3),.cx(input_fmap_53[7:0]),.cy(-9'sd1),.dx(input_fmap_54[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O63_N14_S1),.chainout(chainout_14_O63));
logic signed [63:0] chainout_16_O63; 
logic signed [63:0] O63_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O63(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_55[7:0]),.ay(-9'sd4),.bx(input_fmap_56[7:0]),.by(-9'sd1),.cx(input_fmap_57[7:0]),.cy( 9'sd1),.dx(input_fmap_58[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O63_N16_S1),.chainout(chainout_16_O63));
logic signed [63:0] chainout_18_O63; 
logic signed [63:0] O63_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O63(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_59[7:0]),.ay(-9'sd1),.bx(input_fmap_62[7:0]),.by( 9'sd2),.cx(input_fmap_63[7:0]),.cy( 9'sd3),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O63_N18_S1),.chainout(chainout_18_O63));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O63_N0_S2;		always @(posedge clk) O63_N0_S2 <=     O63_N0_S1  +  O63_N2_S1 ;
 logic signed [21:0] O63_N2_S2;		always @(posedge clk) O63_N2_S2 <=     O63_N4_S1  +  O63_N6_S1 ;
 logic signed [21:0] O63_N4_S2;		always @(posedge clk) O63_N4_S2 <=     O63_N8_S1  +  O63_N10_S1 ;
 logic signed [21:0] O63_N6_S2;		always @(posedge clk) O63_N6_S2 <=     O63_N12_S1  +  O63_N14_S1 ;
 logic signed [21:0] O63_N8_S2;		always @(posedge clk) O63_N8_S2 <=     O63_N16_S1  +  O63_N18_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O63_N0_S3;		always @(posedge clk) O63_N0_S3 <=     O63_N0_S2  +  O63_N2_S2 ;
 logic signed [22:0] O63_N2_S3;		always @(posedge clk) O63_N2_S3 <=     O63_N4_S2  +  O63_N6_S2 ;
 logic signed [22:0] O63_N4_S3;		always @(posedge clk) O63_N4_S3 <=     O63_N8_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O63_N0_S4;		always @(posedge clk) O63_N0_S4 <=     O63_N0_S3  +  O63_N2_S3 ;
 logic signed [23:0] O63_N2_S4;		always @(posedge clk) O63_N2_S4 <=     O63_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O63_N0_S5;		always @(posedge clk) O63_N0_S5 <=     O63_N0_S4  +  O63_N2_S4 ;
 assign conv_mac_63 = O63_N0_S5;

logic valid_D1;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D1<= 0 ;
	else valid_D1<=valid;
end
logic valid_D2;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D2<= 0 ;
	else valid_D2<=valid_D1;
end
logic valid_D3;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D3<= 0 ;
	else valid_D3<=valid_D2;
end
logic valid_D4;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D4<= 0 ;
	else valid_D4<=valid_D3;
end
logic valid_D5;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D5<= 0 ;
	else valid_D5<=valid_D4;
end
logic valid_D6;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D6<= 0 ;
	else valid_D6<=valid_D5;
end
always_ff @(posedge clk) begin
	if (rstn == 0) ready <= 0 ;
	else ready <=valid_D6;
end
logic [31:0] bias_add_0;
assign bias_add_0 = conv_mac_0 + 4'd7;
logic [31:0] bias_add_1;
assign bias_add_1 = conv_mac_1 + 5'd11;
logic [31:0] bias_add_2;
assign bias_add_2 = conv_mac_2 + 5'd12;
logic [31:0] bias_add_3;
assign bias_add_3 = conv_mac_3 + 5'd15;
logic [31:0] bias_add_4;
assign bias_add_4 = conv_mac_4 + 3'd3;
logic [31:0] bias_add_5;
assign bias_add_5 = conv_mac_5 + 5'd8;
logic [31:0] bias_add_6;
assign bias_add_6 = conv_mac_6 + 5'd12;
logic [31:0] bias_add_7;
assign bias_add_7 = conv_mac_7 + 7'd32;
logic [31:0] bias_add_8;
assign bias_add_8 = conv_mac_8 + 5'd14;
logic [31:0] bias_add_9;
assign bias_add_9 = conv_mac_9 + 6'd22;
logic [31:0] bias_add_10;
assign bias_add_10 = conv_mac_10 + 5'd10;
logic [31:0] bias_add_11;
assign bias_add_11 = conv_mac_11 + 6'd16;
logic [31:0] bias_add_12;
assign bias_add_12 = conv_mac_12 - 5'd9;
logic [31:0] bias_add_13;
assign bias_add_13 = conv_mac_13 + 6'd17;
logic [31:0] bias_add_14;
assign bias_add_14 = conv_mac_14 + 6'd25;
logic [31:0] bias_add_15;
assign bias_add_15 = conv_mac_15 + 5'd15;
logic [31:0] bias_add_16;
assign bias_add_16 = conv_mac_16 + 5'd14;
logic [31:0] bias_add_17;
assign bias_add_17 = conv_mac_17 + 6'd24;
logic [31:0] bias_add_18;
assign bias_add_18 = conv_mac_18 + 6'd18;
logic [31:0] bias_add_19;
assign bias_add_19 = conv_mac_19 + 6'd19;
logic [31:0] bias_add_20;
assign bias_add_20 = conv_mac_20 + 5'd13;
logic [31:0] bias_add_21;
assign bias_add_21 = conv_mac_21 + 5'd13;
logic [31:0] bias_add_22;
assign bias_add_22 = conv_mac_22 + 5'd12;
logic [31:0] bias_add_23;
assign bias_add_23 = conv_mac_23 + 4'd4;
logic [31:0] bias_add_24;
assign bias_add_24 = conv_mac_24 + 6'd19;
logic [31:0] bias_add_25;
assign bias_add_25 = conv_mac_25 + 5'd11;
logic [31:0] bias_add_26;
assign bias_add_26 = conv_mac_26 + 2'd1;
logic [31:0] bias_add_27;
assign bias_add_27 = conv_mac_27 + 6'd25;
logic [31:0] bias_add_28;
assign bias_add_28 = conv_mac_28 - 4'd5;
logic [31:0] bias_add_29;
assign bias_add_29 = conv_mac_29 + 2'd1;
logic [31:0] bias_add_30;
assign bias_add_30 = conv_mac_30 + 5'd15;
logic [31:0] bias_add_31;
assign bias_add_31 = conv_mac_31 + 3'd3;
logic [31:0] bias_add_32;
assign bias_add_32 = conv_mac_32 + 5'd10;
logic [31:0] bias_add_33;
assign bias_add_33 = conv_mac_33 + 6'd16;
logic [31:0] bias_add_34;
assign bias_add_34 = conv_mac_34 + 5'd11;
logic [31:0] bias_add_35;
assign bias_add_35 = conv_mac_35 + 4'd7;
logic [31:0] bias_add_36;
assign bias_add_36 = conv_mac_36;
logic [31:0] bias_add_37;
assign bias_add_37 = conv_mac_37 + 6'd17;
logic [31:0] bias_add_38;
assign bias_add_38 = conv_mac_38 + 5'd12;
logic [31:0] bias_add_39;
assign bias_add_39 = conv_mac_39 + 5'd10;
logic [31:0] bias_add_40;
assign bias_add_40 = conv_mac_40 + 4'd6;
logic [31:0] bias_add_41;
assign bias_add_41 = conv_mac_41 - 5'd10;
logic [31:0] bias_add_42;
assign bias_add_42 = conv_mac_42 + 5'd15;
logic [31:0] bias_add_43;
assign bias_add_43 = conv_mac_43 + 6'd16;
logic [31:0] bias_add_44;
assign bias_add_44 = conv_mac_44 + 5'd9;
logic [31:0] bias_add_45;
assign bias_add_45 = conv_mac_45 + 4'd4;
logic [31:0] bias_add_46;
assign bias_add_46 = conv_mac_46 + 5'd15;
logic [31:0] bias_add_47;
assign bias_add_47 = conv_mac_47 + 6'd21;
logic [31:0] bias_add_48;
assign bias_add_48 = conv_mac_48 + 5'd15;
logic [31:0] bias_add_49;
assign bias_add_49 = conv_mac_49 + 3'd3;
logic [31:0] bias_add_50;
assign bias_add_50 = conv_mac_50 + 5'd10;
logic [31:0] bias_add_51;
assign bias_add_51 = conv_mac_51 + 4'd6;
logic [31:0] bias_add_52;
assign bias_add_52 = conv_mac_52 + 4'd6;
logic [31:0] bias_add_53;
assign bias_add_53 = conv_mac_53 + 4'd7;
logic [31:0] bias_add_54;
assign bias_add_54 = conv_mac_54 - 3'd3;
logic [31:0] bias_add_55;
assign bias_add_55 = conv_mac_55 + 5'd13;
logic [31:0] bias_add_56;
assign bias_add_56 = conv_mac_56 + 4'd4;
logic [31:0] bias_add_57;
assign bias_add_57 = conv_mac_57 + 6'd20;
logic [31:0] bias_add_58;
assign bias_add_58 = conv_mac_58 + 6'd16;
logic [31:0] bias_add_59;
assign bias_add_59 = conv_mac_59 + 4'd7;
logic [31:0] bias_add_60;
assign bias_add_60 = conv_mac_60 + 6'd17;
logic [31:0] bias_add_61;
assign bias_add_61 = conv_mac_61 + 6'd18;
logic [31:0] bias_add_62;
assign bias_add_62 = conv_mac_62 + 6'd19;
logic [31:0] bias_add_63;
assign bias_add_63 = conv_mac_63 - 4'd4;

logic [7:0] relu_0;
assign relu_0[7:0] = (bias_add_0[31]==0) ? ((bias_add_0<3'd6) ? {{bias_add_0[31],bias_add_0[10:4]}} :'d6) : '0;
logic [7:0] relu_1;
assign relu_1[7:0] = (bias_add_1[31]==0) ? ((bias_add_1<3'd6) ? {{bias_add_1[31],bias_add_1[10:4]}} :'d6) : '0;
logic [7:0] relu_2;
assign relu_2[7:0] = (bias_add_2[31]==0) ? ((bias_add_2<3'd6) ? {{bias_add_2[31],bias_add_2[10:4]}} :'d6) : '0;
logic [7:0] relu_3;
assign relu_3[7:0] = (bias_add_3[31]==0) ? ((bias_add_3<3'd6) ? {{bias_add_3[31],bias_add_3[10:4]}} :'d6) : '0;
logic [7:0] relu_4;
assign relu_4[7:0] = (bias_add_4[31]==0) ? ((bias_add_4<3'd6) ? {{bias_add_4[31],bias_add_4[10:4]}} :'d6) : '0;
logic [7:0] relu_5;
assign relu_5[7:0] = (bias_add_5[31]==0) ? ((bias_add_5<3'd6) ? {{bias_add_5[31],bias_add_5[10:4]}} :'d6) : '0;
logic [7:0] relu_6;
assign relu_6[7:0] = (bias_add_6[31]==0) ? ((bias_add_6<3'd6) ? {{bias_add_6[31],bias_add_6[10:4]}} :'d6) : '0;
logic [7:0] relu_7;
assign relu_7[7:0] = (bias_add_7[31]==0) ? ((bias_add_7<3'd6) ? {{bias_add_7[31],bias_add_7[10:4]}} :'d6) : '0;
logic [7:0] relu_8;
assign relu_8[7:0] = (bias_add_8[31]==0) ? ((bias_add_8<3'd6) ? {{bias_add_8[31],bias_add_8[10:4]}} :'d6) : '0;
logic [7:0] relu_9;
assign relu_9[7:0] = (bias_add_9[31]==0) ? ((bias_add_9<3'd6) ? {{bias_add_9[31],bias_add_9[10:4]}} :'d6) : '0;
logic [7:0] relu_10;
assign relu_10[7:0] = (bias_add_10[31]==0) ? ((bias_add_10<3'd6) ? {{bias_add_10[31],bias_add_10[10:4]}} :'d6) : '0;
logic [7:0] relu_11;
assign relu_11[7:0] = (bias_add_11[31]==0) ? ((bias_add_11<3'd6) ? {{bias_add_11[31],bias_add_11[10:4]}} :'d6) : '0;
logic [7:0] relu_12;
assign relu_12[7:0] = (bias_add_12[31]==0) ? ((bias_add_12<3'd6) ? {{bias_add_12[31],bias_add_12[10:4]}} :'d6) : '0;
logic [7:0] relu_13;
assign relu_13[7:0] = (bias_add_13[31]==0) ? ((bias_add_13<3'd6) ? {{bias_add_13[31],bias_add_13[10:4]}} :'d6) : '0;
logic [7:0] relu_14;
assign relu_14[7:0] = (bias_add_14[31]==0) ? ((bias_add_14<3'd6) ? {{bias_add_14[31],bias_add_14[10:4]}} :'d6) : '0;
logic [7:0] relu_15;
assign relu_15[7:0] = (bias_add_15[31]==0) ? ((bias_add_15<3'd6) ? {{bias_add_15[31],bias_add_15[10:4]}} :'d6) : '0;
logic [7:0] relu_16;
assign relu_16[7:0] = (bias_add_16[31]==0) ? ((bias_add_16<3'd6) ? {{bias_add_16[31],bias_add_16[10:4]}} :'d6) : '0;
logic [7:0] relu_17;
assign relu_17[7:0] = (bias_add_17[31]==0) ? ((bias_add_17<3'd6) ? {{bias_add_17[31],bias_add_17[10:4]}} :'d6) : '0;
logic [7:0] relu_18;
assign relu_18[7:0] = (bias_add_18[31]==0) ? ((bias_add_18<3'd6) ? {{bias_add_18[31],bias_add_18[10:4]}} :'d6) : '0;
logic [7:0] relu_19;
assign relu_19[7:0] = (bias_add_19[31]==0) ? ((bias_add_19<3'd6) ? {{bias_add_19[31],bias_add_19[10:4]}} :'d6) : '0;
logic [7:0] relu_20;
assign relu_20[7:0] = (bias_add_20[31]==0) ? ((bias_add_20<3'd6) ? {{bias_add_20[31],bias_add_20[10:4]}} :'d6) : '0;
logic [7:0] relu_21;
assign relu_21[7:0] = (bias_add_21[31]==0) ? ((bias_add_21<3'd6) ? {{bias_add_21[31],bias_add_21[10:4]}} :'d6) : '0;
logic [7:0] relu_22;
assign relu_22[7:0] = (bias_add_22[31]==0) ? ((bias_add_22<3'd6) ? {{bias_add_22[31],bias_add_22[10:4]}} :'d6) : '0;
logic [7:0] relu_23;
assign relu_23[7:0] = (bias_add_23[31]==0) ? ((bias_add_23<3'd6) ? {{bias_add_23[31],bias_add_23[10:4]}} :'d6) : '0;
logic [7:0] relu_24;
assign relu_24[7:0] = (bias_add_24[31]==0) ? ((bias_add_24<3'd6) ? {{bias_add_24[31],bias_add_24[10:4]}} :'d6) : '0;
logic [7:0] relu_25;
assign relu_25[7:0] = (bias_add_25[31]==0) ? ((bias_add_25<3'd6) ? {{bias_add_25[31],bias_add_25[10:4]}} :'d6) : '0;
logic [7:0] relu_26;
assign relu_26[7:0] = (bias_add_26[31]==0) ? ((bias_add_26<3'd6) ? {{bias_add_26[31],bias_add_26[10:4]}} :'d6) : '0;
logic [7:0] relu_27;
assign relu_27[7:0] = (bias_add_27[31]==0) ? ((bias_add_27<3'd6) ? {{bias_add_27[31],bias_add_27[10:4]}} :'d6) : '0;
logic [7:0] relu_28;
assign relu_28[7:0] = (bias_add_28[31]==0) ? ((bias_add_28<3'd6) ? {{bias_add_28[31],bias_add_28[10:4]}} :'d6) : '0;
logic [7:0] relu_29;
assign relu_29[7:0] = (bias_add_29[31]==0) ? ((bias_add_29<3'd6) ? {{bias_add_29[31],bias_add_29[10:4]}} :'d6) : '0;
logic [7:0] relu_30;
assign relu_30[7:0] = (bias_add_30[31]==0) ? ((bias_add_30<3'd6) ? {{bias_add_30[31],bias_add_30[10:4]}} :'d6) : '0;
logic [7:0] relu_31;
assign relu_31[7:0] = (bias_add_31[31]==0) ? ((bias_add_31<3'd6) ? {{bias_add_31[31],bias_add_31[10:4]}} :'d6) : '0;
logic [7:0] relu_32;
assign relu_32[7:0] = (bias_add_32[31]==0) ? ((bias_add_32<3'd6) ? {{bias_add_32[31],bias_add_32[10:4]}} :'d6) : '0;
logic [7:0] relu_33;
assign relu_33[7:0] = (bias_add_33[31]==0) ? ((bias_add_33<3'd6) ? {{bias_add_33[31],bias_add_33[10:4]}} :'d6) : '0;
logic [7:0] relu_34;
assign relu_34[7:0] = (bias_add_34[31]==0) ? ((bias_add_34<3'd6) ? {{bias_add_34[31],bias_add_34[10:4]}} :'d6) : '0;
logic [7:0] relu_35;
assign relu_35[7:0] = (bias_add_35[31]==0) ? ((bias_add_35<3'd6) ? {{bias_add_35[31],bias_add_35[10:4]}} :'d6) : '0;
logic [7:0] relu_36;
assign relu_36[7:0] = (bias_add_36[31]==0) ? ((bias_add_36<3'd6) ? {{bias_add_36[31],bias_add_36[10:4]}} :'d6) : '0;
logic [7:0] relu_37;
assign relu_37[7:0] = (bias_add_37[31]==0) ? ((bias_add_37<3'd6) ? {{bias_add_37[31],bias_add_37[10:4]}} :'d6) : '0;
logic [7:0] relu_38;
assign relu_38[7:0] = (bias_add_38[31]==0) ? ((bias_add_38<3'd6) ? {{bias_add_38[31],bias_add_38[10:4]}} :'d6) : '0;
logic [7:0] relu_39;
assign relu_39[7:0] = (bias_add_39[31]==0) ? ((bias_add_39<3'd6) ? {{bias_add_39[31],bias_add_39[10:4]}} :'d6) : '0;
logic [7:0] relu_40;
assign relu_40[7:0] = (bias_add_40[31]==0) ? ((bias_add_40<3'd6) ? {{bias_add_40[31],bias_add_40[10:4]}} :'d6) : '0;
logic [7:0] relu_41;
assign relu_41[7:0] = (bias_add_41[31]==0) ? ((bias_add_41<3'd6) ? {{bias_add_41[31],bias_add_41[10:4]}} :'d6) : '0;
logic [7:0] relu_42;
assign relu_42[7:0] = (bias_add_42[31]==0) ? ((bias_add_42<3'd6) ? {{bias_add_42[31],bias_add_42[10:4]}} :'d6) : '0;
logic [7:0] relu_43;
assign relu_43[7:0] = (bias_add_43[31]==0) ? ((bias_add_43<3'd6) ? {{bias_add_43[31],bias_add_43[10:4]}} :'d6) : '0;
logic [7:0] relu_44;
assign relu_44[7:0] = (bias_add_44[31]==0) ? ((bias_add_44<3'd6) ? {{bias_add_44[31],bias_add_44[10:4]}} :'d6) : '0;
logic [7:0] relu_45;
assign relu_45[7:0] = (bias_add_45[31]==0) ? ((bias_add_45<3'd6) ? {{bias_add_45[31],bias_add_45[10:4]}} :'d6) : '0;
logic [7:0] relu_46;
assign relu_46[7:0] = (bias_add_46[31]==0) ? ((bias_add_46<3'd6) ? {{bias_add_46[31],bias_add_46[10:4]}} :'d6) : '0;
logic [7:0] relu_47;
assign relu_47[7:0] = (bias_add_47[31]==0) ? ((bias_add_47<3'd6) ? {{bias_add_47[31],bias_add_47[10:4]}} :'d6) : '0;
logic [7:0] relu_48;
assign relu_48[7:0] = (bias_add_48[31]==0) ? ((bias_add_48<3'd6) ? {{bias_add_48[31],bias_add_48[10:4]}} :'d6) : '0;
logic [7:0] relu_49;
assign relu_49[7:0] = (bias_add_49[31]==0) ? ((bias_add_49<3'd6) ? {{bias_add_49[31],bias_add_49[10:4]}} :'d6) : '0;
logic [7:0] relu_50;
assign relu_50[7:0] = (bias_add_50[31]==0) ? ((bias_add_50<3'd6) ? {{bias_add_50[31],bias_add_50[10:4]}} :'d6) : '0;
logic [7:0] relu_51;
assign relu_51[7:0] = (bias_add_51[31]==0) ? ((bias_add_51<3'd6) ? {{bias_add_51[31],bias_add_51[10:4]}} :'d6) : '0;
logic [7:0] relu_52;
assign relu_52[7:0] = (bias_add_52[31]==0) ? ((bias_add_52<3'd6) ? {{bias_add_52[31],bias_add_52[10:4]}} :'d6) : '0;
logic [7:0] relu_53;
assign relu_53[7:0] = (bias_add_53[31]==0) ? ((bias_add_53<3'd6) ? {{bias_add_53[31],bias_add_53[10:4]}} :'d6) : '0;
logic [7:0] relu_54;
assign relu_54[7:0] = (bias_add_54[31]==0) ? ((bias_add_54<3'd6) ? {{bias_add_54[31],bias_add_54[10:4]}} :'d6) : '0;
logic [7:0] relu_55;
assign relu_55[7:0] = (bias_add_55[31]==0) ? ((bias_add_55<3'd6) ? {{bias_add_55[31],bias_add_55[10:4]}} :'d6) : '0;
logic [7:0] relu_56;
assign relu_56[7:0] = (bias_add_56[31]==0) ? ((bias_add_56<3'd6) ? {{bias_add_56[31],bias_add_56[10:4]}} :'d6) : '0;
logic [7:0] relu_57;
assign relu_57[7:0] = (bias_add_57[31]==0) ? ((bias_add_57<3'd6) ? {{bias_add_57[31],bias_add_57[10:4]}} :'d6) : '0;
logic [7:0] relu_58;
assign relu_58[7:0] = (bias_add_58[31]==0) ? ((bias_add_58<3'd6) ? {{bias_add_58[31],bias_add_58[10:4]}} :'d6) : '0;
logic [7:0] relu_59;
assign relu_59[7:0] = (bias_add_59[31]==0) ? ((bias_add_59<3'd6) ? {{bias_add_59[31],bias_add_59[10:4]}} :'d6) : '0;
logic [7:0] relu_60;
assign relu_60[7:0] = (bias_add_60[31]==0) ? ((bias_add_60<3'd6) ? {{bias_add_60[31],bias_add_60[10:4]}} :'d6) : '0;
logic [7:0] relu_61;
assign relu_61[7:0] = (bias_add_61[31]==0) ? ((bias_add_61<3'd6) ? {{bias_add_61[31],bias_add_61[10:4]}} :'d6) : '0;
logic [7:0] relu_62;
assign relu_62[7:0] = (bias_add_62[31]==0) ? ((bias_add_62<3'd6) ? {{bias_add_62[31],bias_add_62[10:4]}} :'d6) : '0;
logic [7:0] relu_63;
assign relu_63[7:0] = (bias_add_63[31]==0) ? ((bias_add_63<3'd6) ? {{bias_add_63[31],bias_add_63[10:4]}} :'d6) : '0;

assign output_act = {
	relu_63,
	relu_62,
	relu_61,
	relu_60,
	relu_59,
	relu_58,
	relu_57,
	relu_56,
	relu_55,
	relu_54,
	relu_53,
	relu_52,
	relu_51,
	relu_50,
	relu_49,
	relu_48,
	relu_47,
	relu_46,
	relu_45,
	relu_44,
	relu_43,
	relu_42,
	relu_41,
	relu_40,
	relu_39,
	relu_38,
	relu_37,
	relu_36,
	relu_35,
	relu_34,
	relu_33,
	relu_32,
	relu_31,
	relu_30,
	relu_29,
	relu_28,
	relu_27,
	relu_26,
	relu_25,
	relu_24,
	relu_23,
	relu_22,
	relu_21,
	relu_20,
	relu_19,
	relu_18,
	relu_17,
	relu_16,
	relu_15,
	relu_14,
	relu_13,
	relu_12,
	relu_11,
	relu_10,
	relu_9,
	relu_8,
	relu_7,
	relu_6,
	relu_5,
	relu_4,
	relu_3,
	relu_2,
	relu_1,
	relu_0
};

endmodule
module conv8_pw (
    input logic clk,
    input logic rstn,
    input logic valid,
    input logic [512-1:0] input_act,
    output logic [512-1:0] output_act,
    output logic ready
);
logic we;
logic [8:0] zero_number; 
assign zero_number = 9'd0; 
//1
logic [512-1:0] input_act_ff ;
always_ff @(posedge clk) begin
    if (rstn == 0) begin
        input_act_ff <= '0;
      //  ready <= '0;
    end
    else begin
        input_act_ff <= input_act;
     //   ready <= valid;
    end
end
logic [7:0] input_fmap_0;
assign input_fmap_0 = input_act_ff[7:0];
logic [7:0] input_fmap_1;
assign input_fmap_1 = input_act_ff[15:8];
logic [7:0] input_fmap_2;
assign input_fmap_2 = input_act_ff[23:16];
logic [7:0] input_fmap_3;
assign input_fmap_3 = input_act_ff[31:24];
logic [7:0] input_fmap_4;
assign input_fmap_4 = input_act_ff[39:32];
logic [7:0] input_fmap_5;
assign input_fmap_5 = input_act_ff[47:40];
logic [7:0] input_fmap_6;
assign input_fmap_6 = input_act_ff[55:48];
logic [7:0] input_fmap_7;
assign input_fmap_7 = input_act_ff[63:56];
logic [7:0] input_fmap_8;
assign input_fmap_8 = input_act_ff[71:64];
logic [7:0] input_fmap_9;
assign input_fmap_9 = input_act_ff[79:72];
logic [7:0] input_fmap_10;
assign input_fmap_10 = input_act_ff[87:80];
logic [7:0] input_fmap_11;
assign input_fmap_11 = input_act_ff[95:88];
logic [7:0] input_fmap_12;
assign input_fmap_12 = input_act_ff[103:96];
logic [7:0] input_fmap_13;
assign input_fmap_13 = input_act_ff[111:104];
logic [7:0] input_fmap_14;
assign input_fmap_14 = input_act_ff[119:112];
logic [7:0] input_fmap_15;
assign input_fmap_15 = input_act_ff[127:120];
logic [7:0] input_fmap_16;
assign input_fmap_16 = input_act_ff[135:128];
logic [7:0] input_fmap_17;
assign input_fmap_17 = input_act_ff[143:136];
logic [7:0] input_fmap_18;
assign input_fmap_18 = input_act_ff[151:144];
logic [7:0] input_fmap_19;
assign input_fmap_19 = input_act_ff[159:152];
logic [7:0] input_fmap_20;
assign input_fmap_20 = input_act_ff[167:160];
logic [7:0] input_fmap_21;
assign input_fmap_21 = input_act_ff[175:168];
logic [7:0] input_fmap_22;
assign input_fmap_22 = input_act_ff[183:176];
logic [7:0] input_fmap_23;
assign input_fmap_23 = input_act_ff[191:184];
logic [7:0] input_fmap_24;
assign input_fmap_24 = input_act_ff[199:192];
logic [7:0] input_fmap_25;
assign input_fmap_25 = input_act_ff[207:200];
logic [7:0] input_fmap_26;
assign input_fmap_26 = input_act_ff[215:208];
logic [7:0] input_fmap_27;
assign input_fmap_27 = input_act_ff[223:216];
logic [7:0] input_fmap_28;
assign input_fmap_28 = input_act_ff[231:224];
logic [7:0] input_fmap_29;
assign input_fmap_29 = input_act_ff[239:232];
logic [7:0] input_fmap_30;
assign input_fmap_30 = input_act_ff[247:240];
logic [7:0] input_fmap_31;
assign input_fmap_31 = input_act_ff[255:248];
logic [7:0] input_fmap_32;
assign input_fmap_32 = input_act_ff[263:256];
logic [7:0] input_fmap_33;
assign input_fmap_33 = input_act_ff[271:264];
logic [7:0] input_fmap_34;
assign input_fmap_34 = input_act_ff[279:272];
logic [7:0] input_fmap_35;
assign input_fmap_35 = input_act_ff[287:280];
logic [7:0] input_fmap_36;
assign input_fmap_36 = input_act_ff[295:288];
logic [7:0] input_fmap_37;
assign input_fmap_37 = input_act_ff[303:296];
logic [7:0] input_fmap_38;
assign input_fmap_38 = input_act_ff[311:304];
logic [7:0] input_fmap_39;
assign input_fmap_39 = input_act_ff[319:312];
logic [7:0] input_fmap_40;
assign input_fmap_40 = input_act_ff[327:320];
logic [7:0] input_fmap_41;
assign input_fmap_41 = input_act_ff[335:328];
logic [7:0] input_fmap_42;
assign input_fmap_42 = input_act_ff[343:336];
logic [7:0] input_fmap_43;
assign input_fmap_43 = input_act_ff[351:344];
logic [7:0] input_fmap_44;
assign input_fmap_44 = input_act_ff[359:352];
logic [7:0] input_fmap_45;
assign input_fmap_45 = input_act_ff[367:360];
logic [7:0] input_fmap_46;
assign input_fmap_46 = input_act_ff[375:368];
logic [7:0] input_fmap_47;
assign input_fmap_47 = input_act_ff[383:376];
logic [7:0] input_fmap_48;
assign input_fmap_48 = input_act_ff[391:384];
logic [7:0] input_fmap_49;
assign input_fmap_49 = input_act_ff[399:392];
logic [7:0] input_fmap_50;
assign input_fmap_50 = input_act_ff[407:400];
logic [7:0] input_fmap_51;
assign input_fmap_51 = input_act_ff[415:408];
logic [7:0] input_fmap_52;
assign input_fmap_52 = input_act_ff[423:416];
logic [7:0] input_fmap_53;
assign input_fmap_53 = input_act_ff[431:424];
logic [7:0] input_fmap_54;
assign input_fmap_54 = input_act_ff[439:432];
logic [7:0] input_fmap_55;
assign input_fmap_55 = input_act_ff[447:440];
logic [7:0] input_fmap_56;
assign input_fmap_56 = input_act_ff[455:448];
logic [7:0] input_fmap_57;
assign input_fmap_57 = input_act_ff[463:456];
logic [7:0] input_fmap_58;
assign input_fmap_58 = input_act_ff[471:464];
logic [7:0] input_fmap_59;
assign input_fmap_59 = input_act_ff[479:472];
logic [7:0] input_fmap_60;
assign input_fmap_60 = input_act_ff[487:480];
logic [7:0] input_fmap_61;
assign input_fmap_61 = input_act_ff[495:488];
logic [7:0] input_fmap_62;
assign input_fmap_62 = input_act_ff[503:496];
logic [7:0] input_fmap_63;
assign input_fmap_63 = input_act_ff[511:504];

logic signed [31:0] conv_mac_0;
logic signed [63:0] chainout_0_O0; 
logic signed [63:0] O0_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O0(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay(-9'sd2),.bx(input_fmap_3[7:0]),.by(-9'sd1),.cx(input_fmap_5[7:0]),.cy( 9'sd2),.dx(input_fmap_6[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O0_N0_S1),.chainout(chainout_0_O0));
logic signed [63:0] chainout_2_O0; 
logic signed [63:0] O0_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O0(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_7[7:0]),.ay(-9'sd1),.bx(input_fmap_10[7:0]),.by(-9'sd2),.cx(input_fmap_11[7:0]),.cy( 9'sd1),.dx(input_fmap_12[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O0_N2_S1),.chainout(chainout_2_O0));
logic signed [63:0] chainout_4_O0; 
logic signed [63:0] O0_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O0(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_13[7:0]),.ay( 9'sd1),.bx(input_fmap_14[7:0]),.by(-9'sd1),.cx(input_fmap_17[7:0]),.cy(-9'sd2),.dx(input_fmap_18[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O0_N4_S1),.chainout(chainout_4_O0));
logic signed [63:0] chainout_6_O0; 
logic signed [63:0] O0_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O0(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_20[7:0]),.ay( 9'sd2),.bx(input_fmap_21[7:0]),.by( 9'sd1),.cx(input_fmap_23[7:0]),.cy( 9'sd1),.dx(input_fmap_25[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O0_N6_S1),.chainout(chainout_6_O0));
logic signed [63:0] chainout_8_O0; 
logic signed [63:0] O0_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O0(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_26[7:0]),.ay(-9'sd1),.bx(input_fmap_27[7:0]),.by( 9'sd1),.cx(input_fmap_28[7:0]),.cy( 9'sd1),.dx(input_fmap_29[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O0_N8_S1),.chainout(chainout_8_O0));
logic signed [63:0] chainout_10_O0; 
logic signed [63:0] O0_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O0(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_30[7:0]),.ay(-9'sd2),.bx(input_fmap_32[7:0]),.by( 9'sd1),.cx(input_fmap_34[7:0]),.cy( 9'sd1),.dx(input_fmap_35[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O0_N10_S1),.chainout(chainout_10_O0));
logic signed [63:0] chainout_12_O0; 
logic signed [63:0] O0_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O0(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_36[7:0]),.ay(-9'sd1),.bx(input_fmap_37[7:0]),.by(-9'sd2),.cx(input_fmap_38[7:0]),.cy( 9'sd1),.dx(input_fmap_39[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O0_N12_S1),.chainout(chainout_12_O0));
logic signed [63:0] chainout_14_O0; 
logic signed [63:0] O0_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O0(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_42[7:0]),.ay(-9'sd1),.bx(input_fmap_43[7:0]),.by(-9'sd1),.cx(input_fmap_44[7:0]),.cy(-9'sd1),.dx(input_fmap_46[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O0_N14_S1),.chainout(chainout_14_O0));
logic signed [63:0] chainout_16_O0; 
logic signed [63:0] O0_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O0(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_47[7:0]),.ay(-9'sd1),.bx(input_fmap_48[7:0]),.by(-9'sd2),.cx(input_fmap_50[7:0]),.cy(-9'sd1),.dx(input_fmap_51[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O0_N16_S1),.chainout(chainout_16_O0));
logic signed [63:0] chainout_18_O0; 
logic signed [63:0] O0_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O0(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_52[7:0]),.ay( 9'sd1),.bx(input_fmap_54[7:0]),.by(-9'sd1),.cx(input_fmap_56[7:0]),.cy( 9'sd4),.dx(input_fmap_58[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O0_N18_S1),.chainout(chainout_18_O0));
logic signed [63:0] chainout_20_O0; 
logic signed [63:0] O0_N20_S1; 
 int_sop_4_wrapper int_sop_4_inst_20_O0(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_59[7:0]),.ay( 9'sd1),.bx(input_fmap_62[7:0]),.by(-9'sd1),.cx(input_fmap_63[7:0]),.cy(-9'sd1),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O0_N20_S1),.chainout(chainout_20_O0));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O0_N0_S2;		always @(posedge clk) O0_N0_S2 <=     O0_N0_S1  +  O0_N2_S1 ;
 logic signed [21:0] O0_N2_S2;		always @(posedge clk) O0_N2_S2 <=     O0_N4_S1  +  O0_N6_S1 ;
 logic signed [21:0] O0_N4_S2;		always @(posedge clk) O0_N4_S2 <=     O0_N8_S1  +  O0_N10_S1 ;
 logic signed [21:0] O0_N6_S2;		always @(posedge clk) O0_N6_S2 <=     O0_N12_S1  +  O0_N14_S1 ;
 logic signed [21:0] O0_N8_S2;		always @(posedge clk) O0_N8_S2 <=     O0_N16_S1  +  O0_N18_S1 ;
 logic signed [21:0] O0_N10_S2;		always @(posedge clk) O0_N10_S2 <=     O0_N20_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O0_N0_S3;		always @(posedge clk) O0_N0_S3 <=     O0_N0_S2  +  O0_N2_S2 ;
 logic signed [22:0] O0_N2_S3;		always @(posedge clk) O0_N2_S3 <=     O0_N4_S2  +  O0_N6_S2 ;
 logic signed [22:0] O0_N4_S3;		always @(posedge clk) O0_N4_S3 <=     O0_N8_S2  +  O0_N10_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O0_N0_S4;		always @(posedge clk) O0_N0_S4 <=     O0_N0_S3  +  O0_N2_S3 ;
 logic signed [23:0] O0_N2_S4;		always @(posedge clk) O0_N2_S4 <=     O0_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O0_N0_S5;		always @(posedge clk) O0_N0_S5 <=     O0_N0_S4  +  O0_N2_S4 ;
 assign conv_mac_0 = O0_N0_S5;

logic signed [31:0] conv_mac_1;
logic signed [63:0] chainout_0_O1; 
logic signed [63:0] O1_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O1(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay( 9'sd1),.bx(input_fmap_2[7:0]),.by(-9'sd3),.cx(input_fmap_4[7:0]),.cy( 9'sd1),.dx(input_fmap_5[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O1_N0_S1),.chainout(chainout_0_O1));
logic signed [63:0] chainout_2_O1; 
logic signed [63:0] O1_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O1(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_6[7:0]),.ay( 9'sd1),.bx(input_fmap_7[7:0]),.by(-9'sd1),.cx(input_fmap_8[7:0]),.cy(-9'sd3),.dx(input_fmap_11[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O1_N2_S1),.chainout(chainout_2_O1));
logic signed [63:0] chainout_4_O1; 
logic signed [63:0] O1_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O1(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_14[7:0]),.ay(-9'sd1),.bx(input_fmap_17[7:0]),.by(-9'sd2),.cx(input_fmap_18[7:0]),.cy(-9'sd1),.dx(input_fmap_19[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O1_N4_S1),.chainout(chainout_4_O1));
logic signed [63:0] chainout_6_O1; 
logic signed [63:0] O1_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O1(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_20[7:0]),.ay(-9'sd1),.bx(input_fmap_21[7:0]),.by( 9'sd2),.cx(input_fmap_24[7:0]),.cy(-9'sd1),.dx(input_fmap_25[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O1_N6_S1),.chainout(chainout_6_O1));
logic signed [63:0] chainout_8_O1; 
logic signed [63:0] O1_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O1(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_29[7:0]),.ay( 9'sd1),.bx(input_fmap_33[7:0]),.by( 9'sd2),.cx(input_fmap_34[7:0]),.cy(-9'sd1),.dx(input_fmap_35[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O1_N8_S1),.chainout(chainout_8_O1));
logic signed [63:0] chainout_10_O1; 
logic signed [63:0] O1_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O1(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_37[7:0]),.ay(-9'sd1),.bx(input_fmap_41[7:0]),.by(-9'sd1),.cx(input_fmap_42[7:0]),.cy(-9'sd1),.dx(input_fmap_45[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O1_N10_S1),.chainout(chainout_10_O1));
logic signed [63:0] chainout_12_O1; 
logic signed [63:0] O1_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O1(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_46[7:0]),.ay( 9'sd1),.bx(input_fmap_47[7:0]),.by( 9'sd4),.cx(input_fmap_48[7:0]),.cy( 9'sd2),.dx(input_fmap_49[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O1_N12_S1),.chainout(chainout_12_O1));
logic signed [63:0] chainout_14_O1; 
logic signed [63:0] O1_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O1(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_50[7:0]),.ay( 9'sd1),.bx(input_fmap_51[7:0]),.by(-9'sd2),.cx(input_fmap_52[7:0]),.cy(-9'sd1),.dx(input_fmap_54[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O1_N14_S1),.chainout(chainout_14_O1));
logic signed [63:0] chainout_16_O1; 
logic signed [63:0] O1_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O1(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_58[7:0]),.ay( 9'sd2),.bx(input_fmap_59[7:0]),.by( 9'sd1),.cx(input_fmap_60[7:0]),.cy( 9'sd1),.dx(input_fmap_62[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O1_N16_S1),.chainout(chainout_16_O1));
logic signed [63:0] chainout_18_O1; 
logic signed [63:0] O1_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O1(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_63[7:0]),.ay( 9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O1_N18_S1),.chainout(chainout_18_O1));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O1_N0_S2;		always @(posedge clk) O1_N0_S2 <=     O1_N0_S1  +  O1_N2_S1 ;
 logic signed [21:0] O1_N2_S2;		always @(posedge clk) O1_N2_S2 <=     O1_N4_S1  +  O1_N6_S1 ;
 logic signed [21:0] O1_N4_S2;		always @(posedge clk) O1_N4_S2 <=     O1_N8_S1  +  O1_N10_S1 ;
 logic signed [21:0] O1_N6_S2;		always @(posedge clk) O1_N6_S2 <=     O1_N12_S1  +  O1_N14_S1 ;
 logic signed [21:0] O1_N8_S2;		always @(posedge clk) O1_N8_S2 <=     O1_N16_S1  +  O1_N18_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O1_N0_S3;		always @(posedge clk) O1_N0_S3 <=     O1_N0_S2  +  O1_N2_S2 ;
 logic signed [22:0] O1_N2_S3;		always @(posedge clk) O1_N2_S3 <=     O1_N4_S2  +  O1_N6_S2 ;
 logic signed [22:0] O1_N4_S3;		always @(posedge clk) O1_N4_S3 <=     O1_N8_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O1_N0_S4;		always @(posedge clk) O1_N0_S4 <=     O1_N0_S3  +  O1_N2_S3 ;
 logic signed [23:0] O1_N2_S4;		always @(posedge clk) O1_N2_S4 <=     O1_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O1_N0_S5;		always @(posedge clk) O1_N0_S5 <=     O1_N0_S4  +  O1_N2_S4 ;
 assign conv_mac_1 = O1_N0_S5;

logic signed [31:0] conv_mac_2;
logic signed [63:0] chainout_0_O2; 
logic signed [63:0] O2_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O2(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd2),.bx(input_fmap_1[7:0]),.by( 9'sd1),.cx(input_fmap_2[7:0]),.cy(-9'sd1),.dx(input_fmap_5[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O2_N0_S1),.chainout(chainout_0_O2));
logic signed [63:0] chainout_2_O2; 
logic signed [63:0] O2_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O2(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_6[7:0]),.ay(-9'sd1),.bx(input_fmap_7[7:0]),.by( 9'sd1),.cx(input_fmap_9[7:0]),.cy( 9'sd1),.dx(input_fmap_10[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O2_N2_S1),.chainout(chainout_2_O2));
logic signed [63:0] chainout_4_O2; 
logic signed [63:0] O2_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O2(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_11[7:0]),.ay(-9'sd1),.bx(input_fmap_12[7:0]),.by( 9'sd1),.cx(input_fmap_15[7:0]),.cy( 9'sd1),.dx(input_fmap_16[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O2_N4_S1),.chainout(chainout_4_O2));
logic signed [63:0] chainout_6_O2; 
logic signed [63:0] O2_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O2(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_19[7:0]),.ay( 9'sd1),.bx(input_fmap_22[7:0]),.by(-9'sd1),.cx(input_fmap_23[7:0]),.cy( 9'sd1),.dx(input_fmap_24[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O2_N6_S1),.chainout(chainout_6_O2));
logic signed [63:0] chainout_8_O2; 
logic signed [63:0] O2_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O2(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_26[7:0]),.ay( 9'sd1),.bx(input_fmap_27[7:0]),.by(-9'sd1),.cx(input_fmap_28[7:0]),.cy( 9'sd1),.dx(input_fmap_30[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O2_N8_S1),.chainout(chainout_8_O2));
logic signed [63:0] chainout_10_O2; 
logic signed [63:0] O2_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O2(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_31[7:0]),.ay( 9'sd1),.bx(input_fmap_32[7:0]),.by(-9'sd1),.cx(input_fmap_33[7:0]),.cy( 9'sd1),.dx(input_fmap_35[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O2_N10_S1),.chainout(chainout_10_O2));
logic signed [63:0] chainout_12_O2; 
logic signed [63:0] O2_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O2(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_36[7:0]),.ay( 9'sd1),.bx(input_fmap_37[7:0]),.by( 9'sd1),.cx(input_fmap_38[7:0]),.cy( 9'sd1),.dx(input_fmap_39[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O2_N12_S1),.chainout(chainout_12_O2));
logic signed [63:0] chainout_14_O2; 
logic signed [63:0] O2_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O2(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_41[7:0]),.ay( 9'sd1),.bx(input_fmap_43[7:0]),.by( 9'sd1),.cx(input_fmap_45[7:0]),.cy( 9'sd1),.dx(input_fmap_46[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O2_N14_S1),.chainout(chainout_14_O2));
logic signed [63:0] chainout_16_O2; 
logic signed [63:0] O2_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O2(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_48[7:0]),.ay( 9'sd1),.bx(input_fmap_52[7:0]),.by(-9'sd1),.cx(input_fmap_54[7:0]),.cy( 9'sd1),.dx(input_fmap_57[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O2_N16_S1),.chainout(chainout_16_O2));
logic signed [63:0] chainout_18_O2; 
logic signed [63:0] O2_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O2(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_58[7:0]),.ay( 9'sd4),.bx(input_fmap_59[7:0]),.by( 9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O2_N18_S1),.chainout(chainout_18_O2));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O2_N0_S2;		always @(posedge clk) O2_N0_S2 <=     O2_N0_S1  +  O2_N2_S1 ;
 logic signed [21:0] O2_N2_S2;		always @(posedge clk) O2_N2_S2 <=     O2_N4_S1  +  O2_N6_S1 ;
 logic signed [21:0] O2_N4_S2;		always @(posedge clk) O2_N4_S2 <=     O2_N8_S1  +  O2_N10_S1 ;
 logic signed [21:0] O2_N6_S2;		always @(posedge clk) O2_N6_S2 <=     O2_N12_S1  +  O2_N14_S1 ;
 logic signed [21:0] O2_N8_S2;		always @(posedge clk) O2_N8_S2 <=     O2_N16_S1  +  O2_N18_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O2_N0_S3;		always @(posedge clk) O2_N0_S3 <=     O2_N0_S2  +  O2_N2_S2 ;
 logic signed [22:0] O2_N2_S3;		always @(posedge clk) O2_N2_S3 <=     O2_N4_S2  +  O2_N6_S2 ;
 logic signed [22:0] O2_N4_S3;		always @(posedge clk) O2_N4_S3 <=     O2_N8_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O2_N0_S4;		always @(posedge clk) O2_N0_S4 <=     O2_N0_S3  +  O2_N2_S3 ;
 logic signed [23:0] O2_N2_S4;		always @(posedge clk) O2_N2_S4 <=     O2_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O2_N0_S5;		always @(posedge clk) O2_N0_S5 <=     O2_N0_S4  +  O2_N2_S4 ;
 assign conv_mac_2 = O2_N0_S5;

logic signed [31:0] conv_mac_3;
logic signed [63:0] chainout_0_O3; 
logic signed [63:0] O3_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O3(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_2[7:0]),.ay( 9'sd1),.bx(input_fmap_3[7:0]),.by(-9'sd1),.cx(input_fmap_4[7:0]),.cy(-9'sd1),.dx(input_fmap_5[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O3_N0_S1),.chainout(chainout_0_O3));
logic signed [63:0] chainout_2_O3; 
logic signed [63:0] O3_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O3(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_11[7:0]),.ay(-9'sd1),.bx(input_fmap_13[7:0]),.by( 9'sd1),.cx(input_fmap_19[7:0]),.cy(-9'sd1),.dx(input_fmap_22[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O3_N2_S1),.chainout(chainout_2_O3));
logic signed [63:0] chainout_4_O3; 
logic signed [63:0] O3_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O3(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_25[7:0]),.ay( 9'sd1),.bx(input_fmap_29[7:0]),.by(-9'sd2),.cx(input_fmap_30[7:0]),.cy(-9'sd1),.dx(input_fmap_34[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O3_N4_S1),.chainout(chainout_4_O3));
logic signed [63:0] chainout_6_O3; 
logic signed [63:0] O3_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O3(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_35[7:0]),.ay(-9'sd1),.bx(input_fmap_39[7:0]),.by(-9'sd1),.cx(input_fmap_40[7:0]),.cy( 9'sd1),.dx(input_fmap_43[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O3_N6_S1),.chainout(chainout_6_O3));
logic signed [63:0] chainout_8_O3; 
logic signed [63:0] O3_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O3(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_48[7:0]),.ay(-9'sd1),.bx(input_fmap_49[7:0]),.by(-9'sd1),.cx(input_fmap_50[7:0]),.cy( 9'sd1),.dx(input_fmap_57[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O3_N8_S1),.chainout(chainout_8_O3));
logic signed [63:0] chainout_10_O3; 
logic signed [63:0] O3_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O3(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_60[7:0]),.ay( 9'sd1),.bx(input_fmap_63[7:0]),.by( 9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O3_N10_S1),.chainout(chainout_10_O3));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O3_N0_S2;		always @(posedge clk) O3_N0_S2 <=     O3_N0_S1  +  O3_N2_S1 ;
 logic signed [21:0] O3_N2_S2;		always @(posedge clk) O3_N2_S2 <=     O3_N4_S1  +  O3_N6_S1 ;
 logic signed [21:0] O3_N4_S2;		always @(posedge clk) O3_N4_S2 <=     O3_N8_S1  +  O3_N10_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O3_N0_S3;		always @(posedge clk) O3_N0_S3 <=     O3_N0_S2  +  O3_N2_S2 ;
 logic signed [22:0] O3_N2_S3;		always @(posedge clk) O3_N2_S3 <=     O3_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O3_N0_S4;		always @(posedge clk) O3_N0_S4 <=     O3_N0_S3  +  O3_N2_S3 ;
 assign conv_mac_3 = O3_N0_S4;

logic signed [31:0] conv_mac_4;
logic signed [63:0] chainout_0_O4; 
logic signed [63:0] O4_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O4(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay(-9'sd1),.bx(input_fmap_4[7:0]),.by( 9'sd1),.cx(input_fmap_5[7:0]),.cy(-9'sd1),.dx(input_fmap_10[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O4_N0_S1),.chainout(chainout_0_O4));
logic signed [63:0] chainout_2_O4; 
logic signed [63:0] O4_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O4(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_12[7:0]),.ay(-9'sd1),.bx(input_fmap_13[7:0]),.by( 9'sd1),.cx(input_fmap_20[7:0]),.cy(-9'sd1),.dx(input_fmap_24[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O4_N2_S1),.chainout(chainout_2_O4));
logic signed [63:0] chainout_4_O4; 
logic signed [63:0] O4_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O4(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_25[7:0]),.ay(-9'sd1),.bx(input_fmap_27[7:0]),.by(-9'sd1),.cx(input_fmap_28[7:0]),.cy( 9'sd1),.dx(input_fmap_30[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O4_N4_S1),.chainout(chainout_4_O4));
logic signed [63:0] chainout_6_O4; 
logic signed [63:0] O4_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O4(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_31[7:0]),.ay( 9'sd1),.bx(input_fmap_32[7:0]),.by(-9'sd1),.cx(input_fmap_33[7:0]),.cy(-9'sd2),.dx(input_fmap_34[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O4_N6_S1),.chainout(chainout_6_O4));
logic signed [63:0] chainout_8_O4; 
logic signed [63:0] O4_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O4(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_36[7:0]),.ay(-9'sd1),.bx(input_fmap_38[7:0]),.by(-9'sd1),.cx(input_fmap_40[7:0]),.cy(-9'sd2),.dx(input_fmap_43[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O4_N8_S1),.chainout(chainout_8_O4));
logic signed [63:0] chainout_10_O4; 
logic signed [63:0] O4_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O4(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_46[7:0]),.ay(-9'sd2),.bx(input_fmap_47[7:0]),.by( 9'sd1),.cx(input_fmap_49[7:0]),.cy( 9'sd1),.dx(input_fmap_51[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O4_N10_S1),.chainout(chainout_10_O4));
logic signed [63:0] chainout_12_O4; 
logic signed [63:0] O4_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O4(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_54[7:0]),.ay( 9'sd1),.bx(input_fmap_55[7:0]),.by( 9'sd2),.cx(input_fmap_56[7:0]),.cy( 9'sd1),.dx(input_fmap_57[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O4_N12_S1),.chainout(chainout_12_O4));
logic signed [63:0] chainout_14_O4; 
logic signed [63:0] O4_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O4(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_59[7:0]),.ay(-9'sd1),.bx(input_fmap_60[7:0]),.by(-9'sd1),.cx(input_fmap_61[7:0]),.cy( 9'sd2),.dx(input_fmap_62[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O4_N14_S1),.chainout(chainout_14_O4));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O4_N0_S2;		always @(posedge clk) O4_N0_S2 <=     O4_N0_S1  +  O4_N2_S1 ;
 logic signed [21:0] O4_N2_S2;		always @(posedge clk) O4_N2_S2 <=     O4_N4_S1  +  O4_N6_S1 ;
 logic signed [21:0] O4_N4_S2;		always @(posedge clk) O4_N4_S2 <=     O4_N8_S1  +  O4_N10_S1 ;
 logic signed [21:0] O4_N6_S2;		always @(posedge clk) O4_N6_S2 <=     O4_N12_S1  +  O4_N14_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O4_N0_S3;		always @(posedge clk) O4_N0_S3 <=     O4_N0_S2  +  O4_N2_S2 ;
 logic signed [22:0] O4_N2_S3;		always @(posedge clk) O4_N2_S3 <=     O4_N4_S2  +  O4_N6_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O4_N0_S4;		always @(posedge clk) O4_N0_S4 <=     O4_N0_S3  +  O4_N2_S3 ;
 assign conv_mac_4 = O4_N0_S4;

logic signed [31:0] conv_mac_5;
logic signed [63:0] chainout_0_O5; 
logic signed [63:0] O5_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O5(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd1),.bx(input_fmap_2[7:0]),.by( 9'sd1),.cx(input_fmap_10[7:0]),.cy(-9'sd1),.dx(input_fmap_15[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O5_N0_S1),.chainout(chainout_0_O5));
logic signed [63:0] chainout_2_O5; 
logic signed [63:0] O5_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O5(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_19[7:0]),.ay( 9'sd2),.bx(input_fmap_20[7:0]),.by( 9'sd1),.cx(input_fmap_21[7:0]),.cy( 9'sd1),.dx(input_fmap_25[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O5_N2_S1),.chainout(chainout_2_O5));
logic signed [63:0] chainout_4_O5; 
logic signed [63:0] O5_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O5(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_29[7:0]),.ay(-9'sd1),.bx(input_fmap_34[7:0]),.by( 9'sd1),.cx(input_fmap_35[7:0]),.cy(-9'sd1),.dx(input_fmap_38[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O5_N4_S1),.chainout(chainout_4_O5));
logic signed [63:0] chainout_6_O5; 
logic signed [63:0] O5_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O5(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_40[7:0]),.ay( 9'sd1),.bx(input_fmap_56[7:0]),.by( 9'sd1),.cx(input_fmap_57[7:0]),.cy(-9'sd1),.dx(input_fmap_58[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O5_N6_S1),.chainout(chainout_6_O5));
logic signed [63:0] chainout_8_O5; 
logic signed [63:0] O5_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O5(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_60[7:0]),.ay(-9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O5_N8_S1),.chainout(chainout_8_O5));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O5_N0_S2;		always @(posedge clk) O5_N0_S2 <=     O5_N0_S1  +  O5_N2_S1 ;
 logic signed [21:0] O5_N2_S2;		always @(posedge clk) O5_N2_S2 <=     O5_N4_S1  +  O5_N6_S1 ;
 logic signed [21:0] O5_N4_S2;		always @(posedge clk) O5_N4_S2 <=     O5_N8_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O5_N0_S3;		always @(posedge clk) O5_N0_S3 <=     O5_N0_S2  +  O5_N2_S2 ;
 logic signed [22:0] O5_N2_S3;		always @(posedge clk) O5_N2_S3 <=     O5_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O5_N0_S4;		always @(posedge clk) O5_N0_S4 <=     O5_N0_S3  +  O5_N2_S3 ;
 assign conv_mac_5 = O5_N0_S4;

logic signed [31:0] conv_mac_6;
logic signed [63:0] chainout_0_O6; 
logic signed [63:0] O6_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O6(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_2[7:0]),.ay( 9'sd1),.bx(input_fmap_3[7:0]),.by( 9'sd2),.cx(input_fmap_6[7:0]),.cy( 9'sd1),.dx(input_fmap_8[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O6_N0_S1),.chainout(chainout_0_O6));
logic signed [63:0] chainout_2_O6; 
logic signed [63:0] O6_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O6(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_9[7:0]),.ay(-9'sd1),.bx(input_fmap_10[7:0]),.by( 9'sd1),.cx(input_fmap_12[7:0]),.cy( 9'sd1),.dx(input_fmap_14[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O6_N2_S1),.chainout(chainout_2_O6));
logic signed [63:0] chainout_4_O6; 
logic signed [63:0] O6_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O6(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_15[7:0]),.ay(-9'sd1),.bx(input_fmap_18[7:0]),.by(-9'sd1),.cx(input_fmap_19[7:0]),.cy( 9'sd2),.dx(input_fmap_21[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O6_N4_S1),.chainout(chainout_4_O6));
logic signed [63:0] chainout_6_O6; 
logic signed [63:0] O6_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O6(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_25[7:0]),.ay(-9'sd1),.bx(input_fmap_26[7:0]),.by( 9'sd2),.cx(input_fmap_27[7:0]),.cy(-9'sd1),.dx(input_fmap_29[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O6_N6_S1),.chainout(chainout_6_O6));
logic signed [63:0] chainout_8_O6; 
logic signed [63:0] O6_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O6(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_30[7:0]),.ay(-9'sd2),.bx(input_fmap_31[7:0]),.by( 9'sd1),.cx(input_fmap_35[7:0]),.cy(-9'sd1),.dx(input_fmap_36[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O6_N8_S1),.chainout(chainout_8_O6));
logic signed [63:0] chainout_10_O6; 
logic signed [63:0] O6_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O6(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_37[7:0]),.ay(-9'sd1),.bx(input_fmap_38[7:0]),.by(-9'sd1),.cx(input_fmap_40[7:0]),.cy( 9'sd1),.dx(input_fmap_43[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O6_N10_S1),.chainout(chainout_10_O6));
logic signed [63:0] chainout_12_O6; 
logic signed [63:0] O6_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O6(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_44[7:0]),.ay(-9'sd1),.bx(input_fmap_45[7:0]),.by( 9'sd1),.cx(input_fmap_47[7:0]),.cy(-9'sd1),.dx(input_fmap_48[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O6_N12_S1),.chainout(chainout_12_O6));
logic signed [63:0] chainout_14_O6; 
logic signed [63:0] O6_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O6(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_50[7:0]),.ay( 9'sd1),.bx(input_fmap_52[7:0]),.by( 9'sd1),.cx(input_fmap_54[7:0]),.cy( 9'sd2),.dx(input_fmap_57[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O6_N14_S1),.chainout(chainout_14_O6));
logic signed [63:0] chainout_16_O6; 
logic signed [63:0] O6_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O6(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_58[7:0]),.ay(-9'sd1),.bx(input_fmap_59[7:0]),.by( 9'sd1),.cx(input_fmap_60[7:0]),.cy( 9'sd2),.dx(input_fmap_61[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O6_N16_S1),.chainout(chainout_16_O6));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O6_N0_S2;		always @(posedge clk) O6_N0_S2 <=     O6_N0_S1  +  O6_N2_S1 ;
 logic signed [21:0] O6_N2_S2;		always @(posedge clk) O6_N2_S2 <=     O6_N4_S1  +  O6_N6_S1 ;
 logic signed [21:0] O6_N4_S2;		always @(posedge clk) O6_N4_S2 <=     O6_N8_S1  +  O6_N10_S1 ;
 logic signed [21:0] O6_N6_S2;		always @(posedge clk) O6_N6_S2 <=     O6_N12_S1  +  O6_N14_S1 ;
 logic signed [21:0] O6_N8_S2;		always @(posedge clk) O6_N8_S2 <=     O6_N16_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O6_N0_S3;		always @(posedge clk) O6_N0_S3 <=     O6_N0_S2  +  O6_N2_S2 ;
 logic signed [22:0] O6_N2_S3;		always @(posedge clk) O6_N2_S3 <=     O6_N4_S2  +  O6_N6_S2 ;
 logic signed [22:0] O6_N4_S3;		always @(posedge clk) O6_N4_S3 <=     O6_N8_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O6_N0_S4;		always @(posedge clk) O6_N0_S4 <=     O6_N0_S3  +  O6_N2_S3 ;
 logic signed [23:0] O6_N2_S4;		always @(posedge clk) O6_N2_S4 <=     O6_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O6_N0_S5;		always @(posedge clk) O6_N0_S5 <=     O6_N0_S4  +  O6_N2_S4 ;
 assign conv_mac_6 = O6_N0_S5;

logic signed [31:0] conv_mac_7;
logic signed [63:0] chainout_0_O7; 
logic signed [63:0] O7_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O7(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay(-9'sd1),.bx(input_fmap_2[7:0]),.by( 9'sd1),.cx(input_fmap_4[7:0]),.cy( 9'sd1),.dx(input_fmap_8[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O7_N0_S1),.chainout(chainout_0_O7));
logic signed [63:0] chainout_2_O7; 
logic signed [63:0] O7_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O7(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_10[7:0]),.ay( 9'sd2),.bx(input_fmap_13[7:0]),.by( 9'sd1),.cx(input_fmap_15[7:0]),.cy(-9'sd2),.dx(input_fmap_17[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O7_N2_S1),.chainout(chainout_2_O7));
logic signed [63:0] chainout_4_O7; 
logic signed [63:0] O7_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O7(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_20[7:0]),.ay( 9'sd1),.bx(input_fmap_21[7:0]),.by(-9'sd1),.cx(input_fmap_22[7:0]),.cy(-9'sd1),.dx(input_fmap_24[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O7_N4_S1),.chainout(chainout_4_O7));
logic signed [63:0] chainout_6_O7; 
logic signed [63:0] O7_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O7(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_27[7:0]),.ay(-9'sd1),.bx(input_fmap_28[7:0]),.by( 9'sd1),.cx(input_fmap_32[7:0]),.cy( 9'sd1),.dx(input_fmap_33[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O7_N6_S1),.chainout(chainout_6_O7));
logic signed [63:0] chainout_8_O7; 
logic signed [63:0] O7_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O7(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_34[7:0]),.ay( 9'sd1),.bx(input_fmap_35[7:0]),.by(-9'sd1),.cx(input_fmap_38[7:0]),.cy( 9'sd1),.dx(input_fmap_39[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O7_N8_S1),.chainout(chainout_8_O7));
logic signed [63:0] chainout_10_O7; 
logic signed [63:0] O7_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O7(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_44[7:0]),.ay(-9'sd1),.bx(input_fmap_46[7:0]),.by(-9'sd1),.cx(input_fmap_47[7:0]),.cy( 9'sd1),.dx(input_fmap_48[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O7_N10_S1),.chainout(chainout_10_O7));
logic signed [63:0] chainout_12_O7; 
logic signed [63:0] O7_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O7(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_55[7:0]),.ay( 9'sd1),.bx(input_fmap_57[7:0]),.by(-9'sd2),.cx(input_fmap_58[7:0]),.cy(-9'sd1),.dx(input_fmap_60[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O7_N12_S1),.chainout(chainout_12_O7));
logic signed [63:0] chainout_14_O7; 
logic signed [63:0] O7_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O7(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_61[7:0]),.ay( 9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O7_N14_S1),.chainout(chainout_14_O7));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O7_N0_S2;		always @(posedge clk) O7_N0_S2 <=     O7_N0_S1  +  O7_N2_S1 ;
 logic signed [21:0] O7_N2_S2;		always @(posedge clk) O7_N2_S2 <=     O7_N4_S1  +  O7_N6_S1 ;
 logic signed [21:0] O7_N4_S2;		always @(posedge clk) O7_N4_S2 <=     O7_N8_S1  +  O7_N10_S1 ;
 logic signed [21:0] O7_N6_S2;		always @(posedge clk) O7_N6_S2 <=     O7_N12_S1  +  O7_N14_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O7_N0_S3;		always @(posedge clk) O7_N0_S3 <=     O7_N0_S2  +  O7_N2_S2 ;
 logic signed [22:0] O7_N2_S3;		always @(posedge clk) O7_N2_S3 <=     O7_N4_S2  +  O7_N6_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O7_N0_S4;		always @(posedge clk) O7_N0_S4 <=     O7_N0_S3  +  O7_N2_S3 ;
 assign conv_mac_7 = O7_N0_S4;

logic signed [31:0] conv_mac_8;
logic signed [63:0] chainout_0_O8; 
logic signed [63:0] O8_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O8(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd1),.bx(input_fmap_1[7:0]),.by( 9'sd1),.cx(input_fmap_2[7:0]),.cy( 9'sd2),.dx(input_fmap_5[7:0]),.dy( 9'sd3),.chainin(63'd0),.result(O8_N0_S1),.chainout(chainout_0_O8));
logic signed [63:0] chainout_2_O8; 
logic signed [63:0] O8_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O8(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_8[7:0]),.ay( 9'sd1),.bx(input_fmap_9[7:0]),.by( 9'sd1),.cx(input_fmap_15[7:0]),.cy( 9'sd1),.dx(input_fmap_17[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O8_N2_S1),.chainout(chainout_2_O8));
logic signed [63:0] chainout_4_O8; 
logic signed [63:0] O8_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O8(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_18[7:0]),.ay(-9'sd1),.bx(input_fmap_20[7:0]),.by( 9'sd1),.cx(input_fmap_22[7:0]),.cy( 9'sd1),.dx(input_fmap_23[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O8_N4_S1),.chainout(chainout_4_O8));
logic signed [63:0] chainout_6_O8; 
logic signed [63:0] O8_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O8(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_26[7:0]),.ay( 9'sd1),.bx(input_fmap_27[7:0]),.by( 9'sd1),.cx(input_fmap_32[7:0]),.cy( 9'sd1),.dx(input_fmap_35[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O8_N6_S1),.chainout(chainout_6_O8));
logic signed [63:0] chainout_8_O8; 
logic signed [63:0] O8_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O8(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_37[7:0]),.ay( 9'sd1),.bx(input_fmap_41[7:0]),.by( 9'sd1),.cx(input_fmap_42[7:0]),.cy(-9'sd1),.dx(input_fmap_44[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O8_N8_S1),.chainout(chainout_8_O8));
logic signed [63:0] chainout_10_O8; 
logic signed [63:0] O8_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O8(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_48[7:0]),.ay(-9'sd1),.bx(input_fmap_51[7:0]),.by(-9'sd1),.cx(input_fmap_53[7:0]),.cy( 9'sd1),.dx(input_fmap_54[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O8_N10_S1),.chainout(chainout_10_O8));
logic signed [63:0] chainout_12_O8; 
logic signed [63:0] O8_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O8(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_57[7:0]),.ay( 9'sd1),.bx(input_fmap_61[7:0]),.by(-9'sd1),.cx(input_fmap_63[7:0]),.cy(-9'sd1),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O8_N12_S1),.chainout(chainout_12_O8));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O8_N0_S2;		always @(posedge clk) O8_N0_S2 <=     O8_N0_S1  +  O8_N2_S1 ;
 logic signed [21:0] O8_N2_S2;		always @(posedge clk) O8_N2_S2 <=     O8_N4_S1  +  O8_N6_S1 ;
 logic signed [21:0] O8_N4_S2;		always @(posedge clk) O8_N4_S2 <=     O8_N8_S1  +  O8_N10_S1 ;
 logic signed [21:0] O8_N6_S2;		always @(posedge clk) O8_N6_S2 <=     O8_N12_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O8_N0_S3;		always @(posedge clk) O8_N0_S3 <=     O8_N0_S2  +  O8_N2_S2 ;
 logic signed [22:0] O8_N2_S3;		always @(posedge clk) O8_N2_S3 <=     O8_N4_S2  +  O8_N6_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O8_N0_S4;		always @(posedge clk) O8_N0_S4 <=     O8_N0_S3  +  O8_N2_S3 ;
 assign conv_mac_8 = O8_N0_S4;

logic signed [31:0] conv_mac_9;
logic signed [63:0] chainout_0_O9; 
logic signed [63:0] O9_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O9(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_2[7:0]),.ay( 9'sd1),.bx(input_fmap_5[7:0]),.by(-9'sd1),.cx(input_fmap_13[7:0]),.cy(-9'sd1),.dx(input_fmap_16[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O9_N0_S1),.chainout(chainout_0_O9));
logic signed [63:0] chainout_2_O9; 
logic signed [63:0] O9_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O9(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_19[7:0]),.ay( 9'sd1),.bx(input_fmap_26[7:0]),.by( 9'sd1),.cx(input_fmap_27[7:0]),.cy( 9'sd1),.dx(input_fmap_33[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O9_N2_S1),.chainout(chainout_2_O9));
logic signed [63:0] chainout_4_O9; 
logic signed [63:0] O9_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O9(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_34[7:0]),.ay(-9'sd1),.bx(input_fmap_37[7:0]),.by( 9'sd1),.cx(input_fmap_39[7:0]),.cy(-9'sd1),.dx(input_fmap_41[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O9_N4_S1),.chainout(chainout_4_O9));
logic signed [63:0] chainout_6_O9; 
logic signed [63:0] O9_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O9(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_48[7:0]),.ay(-9'sd1),.bx(input_fmap_49[7:0]),.by(-9'sd1),.cx(input_fmap_51[7:0]),.cy(-9'sd1),.dx(input_fmap_54[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O9_N6_S1),.chainout(chainout_6_O9));
logic signed [63:0] chainout_8_O9; 
logic signed [63:0] O9_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O9(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_55[7:0]),.ay(-9'sd1),.bx(input_fmap_56[7:0]),.by(-9'sd1),.cx(input_fmap_57[7:0]),.cy( 9'sd1),.dx(input_fmap_58[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O9_N8_S1),.chainout(chainout_8_O9));
logic signed [63:0] chainout_10_O9; 
logic signed [63:0] O9_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O9(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_60[7:0]),.ay( 9'sd1),.bx(input_fmap_61[7:0]),.by( 9'sd1),.cx(input_fmap_63[7:0]),.cy( 9'sd1),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O9_N10_S1),.chainout(chainout_10_O9));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O9_N0_S2;		always @(posedge clk) O9_N0_S2 <=     O9_N0_S1  +  O9_N2_S1 ;
 logic signed [21:0] O9_N2_S2;		always @(posedge clk) O9_N2_S2 <=     O9_N4_S1  +  O9_N6_S1 ;
 logic signed [21:0] O9_N4_S2;		always @(posedge clk) O9_N4_S2 <=     O9_N8_S1  +  O9_N10_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O9_N0_S3;		always @(posedge clk) O9_N0_S3 <=     O9_N0_S2  +  O9_N2_S2 ;
 logic signed [22:0] O9_N2_S3;		always @(posedge clk) O9_N2_S3 <=     O9_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O9_N0_S4;		always @(posedge clk) O9_N0_S4 <=     O9_N0_S3  +  O9_N2_S3 ;
 assign conv_mac_9 = O9_N0_S4;

logic signed [31:0] conv_mac_10;
logic signed [63:0] chainout_0_O10; 
logic signed [63:0] O10_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O10(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd1),.bx(input_fmap_1[7:0]),.by(-9'sd2),.cx(input_fmap_2[7:0]),.cy(-9'sd3),.dx(input_fmap_3[7:0]),.dy(-9'sd3),.chainin(63'd0),.result(O10_N0_S1),.chainout(chainout_0_O10));
logic signed [63:0] chainout_2_O10; 
logic signed [63:0] O10_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O10(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_4[7:0]),.ay( 9'sd1),.bx(input_fmap_6[7:0]),.by(-9'sd1),.cx(input_fmap_7[7:0]),.cy( 9'sd3),.dx(input_fmap_8[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O10_N2_S1),.chainout(chainout_2_O10));
logic signed [63:0] chainout_4_O10; 
logic signed [63:0] O10_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O10(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_10[7:0]),.ay(-9'sd2),.bx(input_fmap_11[7:0]),.by( 9'sd2),.cx(input_fmap_12[7:0]),.cy(-9'sd1),.dx(input_fmap_13[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O10_N4_S1),.chainout(chainout_4_O10));
logic signed [63:0] chainout_6_O10; 
logic signed [63:0] O10_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O10(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_14[7:0]),.ay( 9'sd1),.bx(input_fmap_15[7:0]),.by(-9'sd1),.cx(input_fmap_16[7:0]),.cy( 9'sd1),.dx(input_fmap_17[7:0]),.dy(-9'sd3),.chainin(63'd0),.result(O10_N6_S1),.chainout(chainout_6_O10));
logic signed [63:0] chainout_8_O10; 
logic signed [63:0] O10_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O10(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_18[7:0]),.ay( 9'sd1),.bx(input_fmap_19[7:0]),.by( 9'sd3),.cx(input_fmap_22[7:0]),.cy(-9'sd3),.dx(input_fmap_23[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O10_N8_S1),.chainout(chainout_8_O10));
logic signed [63:0] chainout_10_O10; 
logic signed [63:0] O10_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O10(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_24[7:0]),.ay(-9'sd3),.bx(input_fmap_27[7:0]),.by( 9'sd2),.cx(input_fmap_28[7:0]),.cy( 9'sd1),.dx(input_fmap_29[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O10_N10_S1),.chainout(chainout_10_O10));
logic signed [63:0] chainout_12_O10; 
logic signed [63:0] O10_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O10(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_30[7:0]),.ay(-9'sd1),.bx(input_fmap_31[7:0]),.by(-9'sd1),.cx(input_fmap_32[7:0]),.cy(-9'sd1),.dx(input_fmap_33[7:0]),.dy(-9'sd3),.chainin(63'd0),.result(O10_N12_S1),.chainout(chainout_12_O10));
logic signed [63:0] chainout_14_O10; 
logic signed [63:0] O10_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O10(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_36[7:0]),.ay(-9'sd1),.bx(input_fmap_37[7:0]),.by( 9'sd2),.cx(input_fmap_38[7:0]),.cy( 9'sd1),.dx(input_fmap_39[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O10_N14_S1),.chainout(chainout_14_O10));
logic signed [63:0] chainout_16_O10; 
logic signed [63:0] O10_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O10(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_40[7:0]),.ay( 9'sd3),.bx(input_fmap_41[7:0]),.by( 9'sd1),.cx(input_fmap_42[7:0]),.cy( 9'sd1),.dx(input_fmap_44[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O10_N16_S1),.chainout(chainout_16_O10));
logic signed [63:0] chainout_18_O10; 
logic signed [63:0] O10_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O10(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_46[7:0]),.ay( 9'sd3),.bx(input_fmap_47[7:0]),.by( 9'sd2),.cx(input_fmap_48[7:0]),.cy(-9'sd2),.dx(input_fmap_49[7:0]),.dy( 9'sd3),.chainin(63'd0),.result(O10_N18_S1),.chainout(chainout_18_O10));
logic signed [63:0] chainout_20_O10; 
logic signed [63:0] O10_N20_S1; 
 int_sop_4_wrapper int_sop_4_inst_20_O10(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_50[7:0]),.ay(-9'sd1),.bx(input_fmap_51[7:0]),.by( 9'sd1),.cx(input_fmap_52[7:0]),.cy( 9'sd1),.dx(input_fmap_53[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O10_N20_S1),.chainout(chainout_20_O10));
logic signed [63:0] chainout_22_O10; 
logic signed [63:0] O10_N22_S1; 
 int_sop_4_wrapper int_sop_4_inst_22_O10(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_55[7:0]),.ay( 9'sd1),.bx(input_fmap_56[7:0]),.by(-9'sd1),.cx(input_fmap_57[7:0]),.cy(-9'sd1),.dx(input_fmap_58[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O10_N22_S1),.chainout(chainout_22_O10));
logic signed [63:0] chainout_24_O10; 
logic signed [63:0] O10_N24_S1; 
 int_sop_4_wrapper int_sop_4_inst_24_O10(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_62[7:0]),.ay( 9'sd1),.bx(input_fmap_63[7:0]),.by(-9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O10_N24_S1),.chainout(chainout_24_O10));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O10_N0_S2;		always @(posedge clk) O10_N0_S2 <=     O10_N0_S1  +  O10_N2_S1 ;
 logic signed [21:0] O10_N2_S2;		always @(posedge clk) O10_N2_S2 <=     O10_N4_S1  +  O10_N6_S1 ;
 logic signed [21:0] O10_N4_S2;		always @(posedge clk) O10_N4_S2 <=     O10_N8_S1  +  O10_N10_S1 ;
 logic signed [21:0] O10_N6_S2;		always @(posedge clk) O10_N6_S2 <=     O10_N12_S1  +  O10_N14_S1 ;
 logic signed [21:0] O10_N8_S2;		always @(posedge clk) O10_N8_S2 <=     O10_N16_S1  +  O10_N18_S1 ;
 logic signed [21:0] O10_N10_S2;		always @(posedge clk) O10_N10_S2 <=     O10_N20_S1  +  O10_N22_S1 ;
 logic signed [21:0] O10_N12_S2;		always @(posedge clk) O10_N12_S2 <=     O10_N24_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O10_N0_S3;		always @(posedge clk) O10_N0_S3 <=     O10_N0_S2  +  O10_N2_S2 ;
 logic signed [22:0] O10_N2_S3;		always @(posedge clk) O10_N2_S3 <=     O10_N4_S2  +  O10_N6_S2 ;
 logic signed [22:0] O10_N4_S3;		always @(posedge clk) O10_N4_S3 <=     O10_N8_S2  +  O10_N10_S2 ;
 logic signed [22:0] O10_N6_S3;		always @(posedge clk) O10_N6_S3 <=     O10_N12_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O10_N0_S4;		always @(posedge clk) O10_N0_S4 <=     O10_N0_S3  +  O10_N2_S3 ;
 logic signed [23:0] O10_N2_S4;		always @(posedge clk) O10_N2_S4 <=     O10_N4_S3  +  O10_N6_S3 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O10_N0_S5;		always @(posedge clk) O10_N0_S5 <=     O10_N0_S4  +  O10_N2_S4 ;
 assign conv_mac_10 = O10_N0_S5;

logic signed [31:0] conv_mac_11;
logic signed [63:0] chainout_0_O11; 
logic signed [63:0] O11_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O11(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd1),.bx(input_fmap_1[7:0]),.by( 9'sd1),.cx(input_fmap_5[7:0]),.cy(-9'sd1),.dx(input_fmap_7[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O11_N0_S1),.chainout(chainout_0_O11));
logic signed [63:0] chainout_2_O11; 
logic signed [63:0] O11_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O11(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_8[7:0]),.ay(-9'sd1),.bx(input_fmap_12[7:0]),.by(-9'sd1),.cx(input_fmap_13[7:0]),.cy(-9'sd1),.dx(input_fmap_14[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O11_N2_S1),.chainout(chainout_2_O11));
logic signed [63:0] chainout_4_O11; 
logic signed [63:0] O11_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O11(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_17[7:0]),.ay( 9'sd1),.bx(input_fmap_21[7:0]),.by( 9'sd1),.cx(input_fmap_23[7:0]),.cy(-9'sd1),.dx(input_fmap_25[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O11_N4_S1),.chainout(chainout_4_O11));
logic signed [63:0] chainout_6_O11; 
logic signed [63:0] O11_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O11(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_26[7:0]),.ay(-9'sd1),.bx(input_fmap_28[7:0]),.by(-9'sd1),.cx(input_fmap_30[7:0]),.cy(-9'sd1),.dx(input_fmap_36[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O11_N6_S1),.chainout(chainout_6_O11));
logic signed [63:0] chainout_8_O11; 
logic signed [63:0] O11_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O11(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_38[7:0]),.ay(-9'sd1),.bx(input_fmap_40[7:0]),.by( 9'sd2),.cx(input_fmap_42[7:0]),.cy( 9'sd1),.dx(input_fmap_45[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O11_N8_S1),.chainout(chainout_8_O11));
logic signed [63:0] chainout_10_O11; 
logic signed [63:0] O11_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O11(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_46[7:0]),.ay(-9'sd1),.bx(input_fmap_47[7:0]),.by( 9'sd1),.cx(input_fmap_48[7:0]),.cy( 9'sd1),.dx(input_fmap_51[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O11_N10_S1),.chainout(chainout_10_O11));
logic signed [63:0] chainout_12_O11; 
logic signed [63:0] O11_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O11(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_54[7:0]),.ay( 9'sd1),.bx(input_fmap_55[7:0]),.by(-9'sd1),.cx(input_fmap_56[7:0]),.cy(-9'sd1),.dx(input_fmap_57[7:0]),.dy( 9'sd4),.chainin(63'd0),.result(O11_N12_S1),.chainout(chainout_12_O11));
logic signed [63:0] chainout_14_O11; 
logic signed [63:0] O11_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O11(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_59[7:0]),.ay(-9'sd1),.bx(input_fmap_61[7:0]),.by( 9'sd2),.cx(input_fmap_63[7:0]),.cy(-9'sd1),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O11_N14_S1),.chainout(chainout_14_O11));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O11_N0_S2;		always @(posedge clk) O11_N0_S2 <=     O11_N0_S1  +  O11_N2_S1 ;
 logic signed [21:0] O11_N2_S2;		always @(posedge clk) O11_N2_S2 <=     O11_N4_S1  +  O11_N6_S1 ;
 logic signed [21:0] O11_N4_S2;		always @(posedge clk) O11_N4_S2 <=     O11_N8_S1  +  O11_N10_S1 ;
 logic signed [21:0] O11_N6_S2;		always @(posedge clk) O11_N6_S2 <=     O11_N12_S1  +  O11_N14_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O11_N0_S3;		always @(posedge clk) O11_N0_S3 <=     O11_N0_S2  +  O11_N2_S2 ;
 logic signed [22:0] O11_N2_S3;		always @(posedge clk) O11_N2_S3 <=     O11_N4_S2  +  O11_N6_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O11_N0_S4;		always @(posedge clk) O11_N0_S4 <=     O11_N0_S3  +  O11_N2_S3 ;
 assign conv_mac_11 = O11_N0_S4;

logic signed [31:0] conv_mac_12;
logic signed [63:0] chainout_0_O12; 
logic signed [63:0] O12_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O12(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd1),.bx(input_fmap_5[7:0]),.by( 9'sd1),.cx(input_fmap_7[7:0]),.cy( 9'sd2),.dx(input_fmap_8[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O12_N0_S1),.chainout(chainout_0_O12));
logic signed [63:0] chainout_2_O12; 
logic signed [63:0] O12_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O12(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_11[7:0]),.ay(-9'sd1),.bx(input_fmap_15[7:0]),.by(-9'sd1),.cx(input_fmap_18[7:0]),.cy(-9'sd1),.dx(input_fmap_19[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O12_N2_S1),.chainout(chainout_2_O12));
logic signed [63:0] chainout_4_O12; 
logic signed [63:0] O12_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O12(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_20[7:0]),.ay(-9'sd1),.bx(input_fmap_21[7:0]),.by(-9'sd1),.cx(input_fmap_23[7:0]),.cy( 9'sd1),.dx(input_fmap_24[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O12_N4_S1),.chainout(chainout_4_O12));
logic signed [63:0] chainout_6_O12; 
logic signed [63:0] O12_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O12(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_26[7:0]),.ay( 9'sd2),.bx(input_fmap_27[7:0]),.by(-9'sd1),.cx(input_fmap_29[7:0]),.cy(-9'sd1),.dx(input_fmap_33[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O12_N6_S1),.chainout(chainout_6_O12));
logic signed [63:0] chainout_8_O12; 
logic signed [63:0] O12_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O12(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_36[7:0]),.ay(-9'sd1),.bx(input_fmap_41[7:0]),.by( 9'sd1),.cx(input_fmap_42[7:0]),.cy(-9'sd1),.dx(input_fmap_45[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O12_N8_S1),.chainout(chainout_8_O12));
logic signed [63:0] chainout_10_O12; 
logic signed [63:0] O12_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O12(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_47[7:0]),.ay(-9'sd1),.bx(input_fmap_50[7:0]),.by( 9'sd1),.cx(input_fmap_52[7:0]),.cy( 9'sd1),.dx(input_fmap_53[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O12_N10_S1),.chainout(chainout_10_O12));
logic signed [63:0] chainout_12_O12; 
logic signed [63:0] O12_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O12(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_54[7:0]),.ay( 9'sd1),.bx(input_fmap_57[7:0]),.by( 9'sd2),.cx(input_fmap_60[7:0]),.cy( 9'sd1),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O12_N12_S1),.chainout(chainout_12_O12));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O12_N0_S2;		always @(posedge clk) O12_N0_S2 <=     O12_N0_S1  +  O12_N2_S1 ;
 logic signed [21:0] O12_N2_S2;		always @(posedge clk) O12_N2_S2 <=     O12_N4_S1  +  O12_N6_S1 ;
 logic signed [21:0] O12_N4_S2;		always @(posedge clk) O12_N4_S2 <=     O12_N8_S1  +  O12_N10_S1 ;
 logic signed [21:0] O12_N6_S2;		always @(posedge clk) O12_N6_S2 <=     O12_N12_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O12_N0_S3;		always @(posedge clk) O12_N0_S3 <=     O12_N0_S2  +  O12_N2_S2 ;
 logic signed [22:0] O12_N2_S3;		always @(posedge clk) O12_N2_S3 <=     O12_N4_S2  +  O12_N6_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O12_N0_S4;		always @(posedge clk) O12_N0_S4 <=     O12_N0_S3  +  O12_N2_S3 ;
 assign conv_mac_12 = O12_N0_S4;

logic signed [31:0] conv_mac_13;
logic signed [63:0] chainout_0_O13; 
logic signed [63:0] O13_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O13(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_3[7:0]),.ay( 9'sd1),.bx(input_fmap_4[7:0]),.by( 9'sd2),.cx(input_fmap_6[7:0]),.cy(-9'sd1),.dx(input_fmap_7[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O13_N0_S1),.chainout(chainout_0_O13));
logic signed [63:0] chainout_2_O13; 
logic signed [63:0] O13_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O13(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_8[7:0]),.ay( 9'sd1),.bx(input_fmap_10[7:0]),.by(-9'sd2),.cx(input_fmap_11[7:0]),.cy( 9'sd1),.dx(input_fmap_12[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O13_N2_S1),.chainout(chainout_2_O13));
logic signed [63:0] chainout_4_O13; 
logic signed [63:0] O13_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O13(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_13[7:0]),.ay( 9'sd1),.bx(input_fmap_14[7:0]),.by( 9'sd1),.cx(input_fmap_16[7:0]),.cy( 9'sd3),.dx(input_fmap_19[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O13_N4_S1),.chainout(chainout_4_O13));
logic signed [63:0] chainout_6_O13; 
logic signed [63:0] O13_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O13(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_21[7:0]),.ay(-9'sd1),.bx(input_fmap_22[7:0]),.by( 9'sd1),.cx(input_fmap_23[7:0]),.cy( 9'sd1),.dx(input_fmap_24[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O13_N6_S1),.chainout(chainout_6_O13));
logic signed [63:0] chainout_8_O13; 
logic signed [63:0] O13_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O13(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_31[7:0]),.ay(-9'sd1),.bx(input_fmap_33[7:0]),.by( 9'sd1),.cx(input_fmap_35[7:0]),.cy(-9'sd1),.dx(input_fmap_37[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O13_N8_S1),.chainout(chainout_8_O13));
logic signed [63:0] chainout_10_O13; 
logic signed [63:0] O13_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O13(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_39[7:0]),.ay(-9'sd1),.bx(input_fmap_41[7:0]),.by( 9'sd1),.cx(input_fmap_43[7:0]),.cy( 9'sd1),.dx(input_fmap_44[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O13_N10_S1),.chainout(chainout_10_O13));
logic signed [63:0] chainout_12_O13; 
logic signed [63:0] O13_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O13(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_47[7:0]),.ay(-9'sd1),.bx(input_fmap_49[7:0]),.by( 9'sd1),.cx(input_fmap_53[7:0]),.cy(-9'sd1),.dx(input_fmap_55[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O13_N12_S1),.chainout(chainout_12_O13));
logic signed [63:0] chainout_14_O13; 
logic signed [63:0] O13_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O13(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_56[7:0]),.ay( 9'sd1),.bx(input_fmap_57[7:0]),.by( 9'sd1),.cx(input_fmap_58[7:0]),.cy(-9'sd1),.dx(input_fmap_59[7:0]),.dy( 9'sd3),.chainin(63'd0),.result(O13_N14_S1),.chainout(chainout_14_O13));
logic signed [63:0] chainout_16_O13; 
logic signed [63:0] O13_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O13(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_60[7:0]),.ay(-9'sd1),.bx(input_fmap_63[7:0]),.by(-9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O13_N16_S1),.chainout(chainout_16_O13));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O13_N0_S2;		always @(posedge clk) O13_N0_S2 <=     O13_N0_S1  +  O13_N2_S1 ;
 logic signed [21:0] O13_N2_S2;		always @(posedge clk) O13_N2_S2 <=     O13_N4_S1  +  O13_N6_S1 ;
 logic signed [21:0] O13_N4_S2;		always @(posedge clk) O13_N4_S2 <=     O13_N8_S1  +  O13_N10_S1 ;
 logic signed [21:0] O13_N6_S2;		always @(posedge clk) O13_N6_S2 <=     O13_N12_S1  +  O13_N14_S1 ;
 logic signed [21:0] O13_N8_S2;		always @(posedge clk) O13_N8_S2 <=     O13_N16_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O13_N0_S3;		always @(posedge clk) O13_N0_S3 <=     O13_N0_S2  +  O13_N2_S2 ;
 logic signed [22:0] O13_N2_S3;		always @(posedge clk) O13_N2_S3 <=     O13_N4_S2  +  O13_N6_S2 ;
 logic signed [22:0] O13_N4_S3;		always @(posedge clk) O13_N4_S3 <=     O13_N8_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O13_N0_S4;		always @(posedge clk) O13_N0_S4 <=     O13_N0_S3  +  O13_N2_S3 ;
 logic signed [23:0] O13_N2_S4;		always @(posedge clk) O13_N2_S4 <=     O13_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O13_N0_S5;		always @(posedge clk) O13_N0_S5 <=     O13_N0_S4  +  O13_N2_S4 ;
 assign conv_mac_13 = O13_N0_S5;

logic signed [31:0] conv_mac_14;
logic signed [63:0] chainout_0_O14; 
logic signed [63:0] O14_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O14(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay(-9'sd2),.bx(input_fmap_2[7:0]),.by(-9'sd2),.cx(input_fmap_3[7:0]),.cy( 9'sd1),.dx(input_fmap_7[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O14_N0_S1),.chainout(chainout_0_O14));
logic signed [63:0] chainout_2_O14; 
logic signed [63:0] O14_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O14(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_8[7:0]),.ay(-9'sd2),.bx(input_fmap_10[7:0]),.by(-9'sd2),.cx(input_fmap_12[7:0]),.cy( 9'sd1),.dx(input_fmap_14[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O14_N2_S1),.chainout(chainout_2_O14));
logic signed [63:0] chainout_4_O14; 
logic signed [63:0] O14_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O14(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_15[7:0]),.ay( 9'sd1),.bx(input_fmap_16[7:0]),.by(-9'sd1),.cx(input_fmap_17[7:0]),.cy(-9'sd1),.dx(input_fmap_18[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O14_N4_S1),.chainout(chainout_4_O14));
logic signed [63:0] chainout_6_O14; 
logic signed [63:0] O14_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O14(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_19[7:0]),.ay(-9'sd2),.bx(input_fmap_22[7:0]),.by( 9'sd2),.cx(input_fmap_23[7:0]),.cy( 9'sd1),.dx(input_fmap_25[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O14_N6_S1),.chainout(chainout_6_O14));
logic signed [63:0] chainout_8_O14; 
logic signed [63:0] O14_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O14(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_26[7:0]),.ay( 9'sd1),.bx(input_fmap_27[7:0]),.by(-9'sd1),.cx(input_fmap_28[7:0]),.cy(-9'sd2),.dx(input_fmap_30[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O14_N8_S1),.chainout(chainout_8_O14));
logic signed [63:0] chainout_10_O14; 
logic signed [63:0] O14_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O14(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_31[7:0]),.ay( 9'sd1),.bx(input_fmap_35[7:0]),.by(-9'sd1),.cx(input_fmap_37[7:0]),.cy( 9'sd1),.dx(input_fmap_38[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O14_N10_S1),.chainout(chainout_10_O14));
logic signed [63:0] chainout_12_O14; 
logic signed [63:0] O14_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O14(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_40[7:0]),.ay(-9'sd1),.bx(input_fmap_42[7:0]),.by( 9'sd1),.cx(input_fmap_43[7:0]),.cy( 9'sd1),.dx(input_fmap_47[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O14_N12_S1),.chainout(chainout_12_O14));
logic signed [63:0] chainout_14_O14; 
logic signed [63:0] O14_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O14(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_50[7:0]),.ay( 9'sd1),.bx(input_fmap_51[7:0]),.by(-9'sd1),.cx(input_fmap_52[7:0]),.cy(-9'sd1),.dx(input_fmap_53[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O14_N14_S1),.chainout(chainout_14_O14));
logic signed [63:0] chainout_16_O14; 
logic signed [63:0] O14_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O14(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_54[7:0]),.ay( 9'sd1),.bx(input_fmap_58[7:0]),.by(-9'sd1),.cx(input_fmap_59[7:0]),.cy(-9'sd1),.dx(input_fmap_60[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O14_N16_S1),.chainout(chainout_16_O14));
logic signed [63:0] chainout_18_O14; 
logic signed [63:0] O14_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O14(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_62[7:0]),.ay(-9'sd1),.bx(input_fmap_63[7:0]),.by(-9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O14_N18_S1),.chainout(chainout_18_O14));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O14_N0_S2;		always @(posedge clk) O14_N0_S2 <=     O14_N0_S1  +  O14_N2_S1 ;
 logic signed [21:0] O14_N2_S2;		always @(posedge clk) O14_N2_S2 <=     O14_N4_S1  +  O14_N6_S1 ;
 logic signed [21:0] O14_N4_S2;		always @(posedge clk) O14_N4_S2 <=     O14_N8_S1  +  O14_N10_S1 ;
 logic signed [21:0] O14_N6_S2;		always @(posedge clk) O14_N6_S2 <=     O14_N12_S1  +  O14_N14_S1 ;
 logic signed [21:0] O14_N8_S2;		always @(posedge clk) O14_N8_S2 <=     O14_N16_S1  +  O14_N18_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O14_N0_S3;		always @(posedge clk) O14_N0_S3 <=     O14_N0_S2  +  O14_N2_S2 ;
 logic signed [22:0] O14_N2_S3;		always @(posedge clk) O14_N2_S3 <=     O14_N4_S2  +  O14_N6_S2 ;
 logic signed [22:0] O14_N4_S3;		always @(posedge clk) O14_N4_S3 <=     O14_N8_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O14_N0_S4;		always @(posedge clk) O14_N0_S4 <=     O14_N0_S3  +  O14_N2_S3 ;
 logic signed [23:0] O14_N2_S4;		always @(posedge clk) O14_N2_S4 <=     O14_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O14_N0_S5;		always @(posedge clk) O14_N0_S5 <=     O14_N0_S4  +  O14_N2_S4 ;
 assign conv_mac_14 = O14_N0_S5;

logic signed [31:0] conv_mac_15;
logic signed [63:0] chainout_0_O15; 
logic signed [63:0] O15_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O15(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_5[7:0]),.ay( 9'sd1),.bx(input_fmap_8[7:0]),.by( 9'sd1),.cx(input_fmap_11[7:0]),.cy(-9'sd1),.dx(input_fmap_13[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O15_N0_S1),.chainout(chainout_0_O15));
logic signed [63:0] chainout_2_O15; 
logic signed [63:0] O15_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O15(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_22[7:0]),.ay(-9'sd1),.bx(input_fmap_23[7:0]),.by(-9'sd1),.cx(input_fmap_24[7:0]),.cy(-9'sd1),.dx(input_fmap_34[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O15_N2_S1),.chainout(chainout_2_O15));
logic signed [63:0] chainout_4_O15; 
logic signed [63:0] O15_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O15(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_37[7:0]),.ay( 9'sd1),.bx(input_fmap_38[7:0]),.by(-9'sd1),.cx(input_fmap_39[7:0]),.cy( 9'sd1),.dx(input_fmap_40[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O15_N4_S1),.chainout(chainout_4_O15));
logic signed [63:0] chainout_6_O15; 
logic signed [63:0] O15_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O15(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_42[7:0]),.ay(-9'sd1),.bx(input_fmap_43[7:0]),.by( 9'sd1),.cx(input_fmap_45[7:0]),.cy( 9'sd1),.dx(input_fmap_46[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O15_N6_S1),.chainout(chainout_6_O15));
logic signed [63:0] chainout_8_O15; 
logic signed [63:0] O15_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O15(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_47[7:0]),.ay( 9'sd1),.bx(input_fmap_53[7:0]),.by( 9'sd1),.cx(input_fmap_57[7:0]),.cy( 9'sd1),.dx(input_fmap_60[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O15_N8_S1),.chainout(chainout_8_O15));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O15_N0_S2;		always @(posedge clk) O15_N0_S2 <=     O15_N0_S1  +  O15_N2_S1 ;
 logic signed [21:0] O15_N2_S2;		always @(posedge clk) O15_N2_S2 <=     O15_N4_S1  +  O15_N6_S1 ;
 logic signed [21:0] O15_N4_S2;		always @(posedge clk) O15_N4_S2 <=     O15_N8_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O15_N0_S3;		always @(posedge clk) O15_N0_S3 <=     O15_N0_S2  +  O15_N2_S2 ;
 logic signed [22:0] O15_N2_S3;		always @(posedge clk) O15_N2_S3 <=     O15_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O15_N0_S4;		always @(posedge clk) O15_N0_S4 <=     O15_N0_S3  +  O15_N2_S3 ;
 assign conv_mac_15 = O15_N0_S4;

logic signed [31:0] conv_mac_16;
logic signed [63:0] chainout_0_O16; 
logic signed [63:0] O16_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O16(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd1),.bx(input_fmap_1[7:0]),.by( 9'sd4),.cx(input_fmap_2[7:0]),.cy(-9'sd1),.dx(input_fmap_4[7:0]),.dy( 9'sd3),.chainin(63'd0),.result(O16_N0_S1),.chainout(chainout_0_O16));
logic signed [63:0] chainout_2_O16; 
logic signed [63:0] O16_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O16(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_5[7:0]),.ay(-9'sd4),.bx(input_fmap_8[7:0]),.by( 9'sd1),.cx(input_fmap_9[7:0]),.cy( 9'sd1),.dx(input_fmap_10[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O16_N2_S1),.chainout(chainout_2_O16));
logic signed [63:0] chainout_4_O16; 
logic signed [63:0] O16_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O16(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_11[7:0]),.ay( 9'sd1),.bx(input_fmap_12[7:0]),.by(-9'sd1),.cx(input_fmap_18[7:0]),.cy(-9'sd3),.dx(input_fmap_19[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O16_N4_S1),.chainout(chainout_4_O16));
logic signed [63:0] chainout_6_O16; 
logic signed [63:0] O16_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O16(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_20[7:0]),.ay(-9'sd2),.bx(input_fmap_21[7:0]),.by(-9'sd1),.cx(input_fmap_23[7:0]),.cy( 9'sd1),.dx(input_fmap_25[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O16_N6_S1),.chainout(chainout_6_O16));
logic signed [63:0] chainout_8_O16; 
logic signed [63:0] O16_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O16(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_26[7:0]),.ay( 9'sd2),.bx(input_fmap_28[7:0]),.by( 9'sd1),.cx(input_fmap_29[7:0]),.cy(-9'sd1),.dx(input_fmap_30[7:0]),.dy( 9'sd3),.chainin(63'd0),.result(O16_N8_S1),.chainout(chainout_8_O16));
logic signed [63:0] chainout_10_O16; 
logic signed [63:0] O16_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O16(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_31[7:0]),.ay( 9'sd2),.bx(input_fmap_33[7:0]),.by( 9'sd2),.cx(input_fmap_34[7:0]),.cy(-9'sd1),.dx(input_fmap_35[7:0]),.dy(-9'sd3),.chainin(63'd0),.result(O16_N10_S1),.chainout(chainout_10_O16));
logic signed [63:0] chainout_12_O16; 
logic signed [63:0] O16_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O16(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_36[7:0]),.ay( 9'sd2),.bx(input_fmap_37[7:0]),.by( 9'sd2),.cx(input_fmap_38[7:0]),.cy( 9'sd2),.dx(input_fmap_39[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O16_N12_S1),.chainout(chainout_12_O16));
logic signed [63:0] chainout_14_O16; 
logic signed [63:0] O16_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O16(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_40[7:0]),.ay(-9'sd1),.bx(input_fmap_42[7:0]),.by(-9'sd1),.cx(input_fmap_43[7:0]),.cy(-9'sd1),.dx(input_fmap_44[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O16_N14_S1),.chainout(chainout_14_O16));
logic signed [63:0] chainout_16_O16; 
logic signed [63:0] O16_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O16(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_45[7:0]),.ay( 9'sd1),.bx(input_fmap_46[7:0]),.by(-9'sd1),.cx(input_fmap_48[7:0]),.cy( 9'sd1),.dx(input_fmap_49[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O16_N16_S1),.chainout(chainout_16_O16));
logic signed [63:0] chainout_18_O16; 
logic signed [63:0] O16_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O16(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_50[7:0]),.ay( 9'sd1),.bx(input_fmap_51[7:0]),.by(-9'sd1),.cx(input_fmap_53[7:0]),.cy(-9'sd3),.dx(input_fmap_54[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O16_N18_S1),.chainout(chainout_18_O16));
logic signed [63:0] chainout_20_O16; 
logic signed [63:0] O16_N20_S1; 
 int_sop_4_wrapper int_sop_4_inst_20_O16(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_56[7:0]),.ay( 9'sd3),.bx(input_fmap_58[7:0]),.by( 9'sd2),.cx(input_fmap_59[7:0]),.cy(-9'sd1),.dx(input_fmap_60[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O16_N20_S1),.chainout(chainout_20_O16));
logic signed [63:0] chainout_22_O16; 
logic signed [63:0] O16_N22_S1; 
 int_sop_4_wrapper int_sop_4_inst_22_O16(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_61[7:0]),.ay(-9'sd1),.bx(input_fmap_62[7:0]),.by(-9'sd2),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O16_N22_S1),.chainout(chainout_22_O16));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O16_N0_S2;		always @(posedge clk) O16_N0_S2 <=     O16_N0_S1  +  O16_N2_S1 ;
 logic signed [21:0] O16_N2_S2;		always @(posedge clk) O16_N2_S2 <=     O16_N4_S1  +  O16_N6_S1 ;
 logic signed [21:0] O16_N4_S2;		always @(posedge clk) O16_N4_S2 <=     O16_N8_S1  +  O16_N10_S1 ;
 logic signed [21:0] O16_N6_S2;		always @(posedge clk) O16_N6_S2 <=     O16_N12_S1  +  O16_N14_S1 ;
 logic signed [21:0] O16_N8_S2;		always @(posedge clk) O16_N8_S2 <=     O16_N16_S1  +  O16_N18_S1 ;
 logic signed [21:0] O16_N10_S2;		always @(posedge clk) O16_N10_S2 <=     O16_N20_S1  +  O16_N22_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O16_N0_S3;		always @(posedge clk) O16_N0_S3 <=     O16_N0_S2  +  O16_N2_S2 ;
 logic signed [22:0] O16_N2_S3;		always @(posedge clk) O16_N2_S3 <=     O16_N4_S2  +  O16_N6_S2 ;
 logic signed [22:0] O16_N4_S3;		always @(posedge clk) O16_N4_S3 <=     O16_N8_S2  +  O16_N10_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O16_N0_S4;		always @(posedge clk) O16_N0_S4 <=     O16_N0_S3  +  O16_N2_S3 ;
 logic signed [23:0] O16_N2_S4;		always @(posedge clk) O16_N2_S4 <=     O16_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O16_N0_S5;		always @(posedge clk) O16_N0_S5 <=     O16_N0_S4  +  O16_N2_S4 ;
 assign conv_mac_16 = O16_N0_S5;

logic signed [31:0] conv_mac_17;
logic signed [63:0] chainout_0_O17; 
logic signed [63:0] O17_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O17(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_8[7:0]),.ay(-9'sd1),.bx(input_fmap_12[7:0]),.by( 9'sd1),.cx(input_fmap_19[7:0]),.cy(-9'sd1),.dx(input_fmap_20[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O17_N0_S1),.chainout(chainout_0_O17));
logic signed [63:0] chainout_2_O17; 
logic signed [63:0] O17_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O17(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_22[7:0]),.ay( 9'sd1),.bx(input_fmap_23[7:0]),.by(-9'sd1),.cx(input_fmap_34[7:0]),.cy( 9'sd1),.dx(input_fmap_38[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O17_N2_S1),.chainout(chainout_2_O17));
logic signed [63:0] chainout_4_O17; 
logic signed [63:0] O17_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O17(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_40[7:0]),.ay( 9'sd1),.bx(input_fmap_43[7:0]),.by( 9'sd1),.cx(input_fmap_44[7:0]),.cy(-9'sd1),.dx(input_fmap_46[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O17_N4_S1),.chainout(chainout_4_O17));
logic signed [63:0] chainout_6_O17; 
logic signed [63:0] O17_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O17(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_47[7:0]),.ay( 9'sd1),.bx(input_fmap_50[7:0]),.by( 9'sd1),.cx(input_fmap_51[7:0]),.cy( 9'sd1),.dx(input_fmap_54[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O17_N6_S1),.chainout(chainout_6_O17));
logic signed [63:0] chainout_8_O17; 
logic signed [63:0] O17_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O17(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_58[7:0]),.ay(-9'sd1),.bx(input_fmap_60[7:0]),.by(-9'sd1),.cx(input_fmap_62[7:0]),.cy(-9'sd1),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O17_N8_S1),.chainout(chainout_8_O17));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O17_N0_S2;		always @(posedge clk) O17_N0_S2 <=     O17_N0_S1  +  O17_N2_S1 ;
 logic signed [21:0] O17_N2_S2;		always @(posedge clk) O17_N2_S2 <=     O17_N4_S1  +  O17_N6_S1 ;
 logic signed [21:0] O17_N4_S2;		always @(posedge clk) O17_N4_S2 <=     O17_N8_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O17_N0_S3;		always @(posedge clk) O17_N0_S3 <=     O17_N0_S2  +  O17_N2_S2 ;
 logic signed [22:0] O17_N2_S3;		always @(posedge clk) O17_N2_S3 <=     O17_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O17_N0_S4;		always @(posedge clk) O17_N0_S4 <=     O17_N0_S3  +  O17_N2_S3 ;
 assign conv_mac_17 = O17_N0_S4;

logic signed [31:0] conv_mac_18;
logic signed [63:0] chainout_0_O18; 
logic signed [63:0] O18_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O18(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd1),.bx(input_fmap_1[7:0]),.by(-9'sd1),.cx(input_fmap_3[7:0]),.cy(-9'sd1),.dx(input_fmap_6[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O18_N0_S1),.chainout(chainout_0_O18));
logic signed [63:0] chainout_2_O18; 
logic signed [63:0] O18_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O18(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_7[7:0]),.ay( 9'sd1),.bx(input_fmap_8[7:0]),.by(-9'sd1),.cx(input_fmap_10[7:0]),.cy(-9'sd2),.dx(input_fmap_11[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O18_N2_S1),.chainout(chainout_2_O18));
logic signed [63:0] chainout_4_O18; 
logic signed [63:0] O18_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O18(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_12[7:0]),.ay( 9'sd1),.bx(input_fmap_13[7:0]),.by( 9'sd1),.cx(input_fmap_14[7:0]),.cy(-9'sd2),.dx(input_fmap_15[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O18_N4_S1),.chainout(chainout_4_O18));
logic signed [63:0] chainout_6_O18; 
logic signed [63:0] O18_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O18(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_16[7:0]),.ay(-9'sd1),.bx(input_fmap_18[7:0]),.by(-9'sd1),.cx(input_fmap_19[7:0]),.cy(-9'sd2),.dx(input_fmap_20[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O18_N6_S1),.chainout(chainout_6_O18));
logic signed [63:0] chainout_8_O18; 
logic signed [63:0] O18_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O18(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_21[7:0]),.ay( 9'sd4),.bx(input_fmap_22[7:0]),.by(-9'sd1),.cx(input_fmap_23[7:0]),.cy( 9'sd1),.dx(input_fmap_24[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O18_N8_S1),.chainout(chainout_8_O18));
logic signed [63:0] chainout_10_O18; 
logic signed [63:0] O18_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O18(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_26[7:0]),.ay( 9'sd1),.bx(input_fmap_27[7:0]),.by(-9'sd1),.cx(input_fmap_28[7:0]),.cy(-9'sd1),.dx(input_fmap_29[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O18_N10_S1),.chainout(chainout_10_O18));
logic signed [63:0] chainout_12_O18; 
logic signed [63:0] O18_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O18(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_31[7:0]),.ay(-9'sd1),.bx(input_fmap_32[7:0]),.by(-9'sd1),.cx(input_fmap_37[7:0]),.cy( 9'sd1),.dx(input_fmap_39[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O18_N12_S1),.chainout(chainout_12_O18));
logic signed [63:0] chainout_14_O18; 
logic signed [63:0] O18_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O18(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_40[7:0]),.ay( 9'sd1),.bx(input_fmap_41[7:0]),.by( 9'sd3),.cx(input_fmap_44[7:0]),.cy(-9'sd1),.dx(input_fmap_45[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O18_N14_S1),.chainout(chainout_14_O18));
logic signed [63:0] chainout_16_O18; 
logic signed [63:0] O18_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O18(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_47[7:0]),.ay(-9'sd2),.bx(input_fmap_48[7:0]),.by( 9'sd1),.cx(input_fmap_49[7:0]),.cy( 9'sd1),.dx(input_fmap_50[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O18_N16_S1),.chainout(chainout_16_O18));
logic signed [63:0] chainout_18_O18; 
logic signed [63:0] O18_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O18(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_51[7:0]),.ay( 9'sd2),.bx(input_fmap_54[7:0]),.by(-9'sd1),.cx(input_fmap_58[7:0]),.cy(-9'sd1),.dx(input_fmap_59[7:0]),.dy( 9'sd3),.chainin(63'd0),.result(O18_N18_S1),.chainout(chainout_18_O18));
logic signed [63:0] chainout_20_O18; 
logic signed [63:0] O18_N20_S1; 
 int_sop_4_wrapper int_sop_4_inst_20_O18(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_61[7:0]),.ay( 9'sd2),.bx(input_fmap_62[7:0]),.by(-9'sd1),.cx(input_fmap_63[7:0]),.cy(-9'sd1),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O18_N20_S1),.chainout(chainout_20_O18));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O18_N0_S2;		always @(posedge clk) O18_N0_S2 <=     O18_N0_S1  +  O18_N2_S1 ;
 logic signed [21:0] O18_N2_S2;		always @(posedge clk) O18_N2_S2 <=     O18_N4_S1  +  O18_N6_S1 ;
 logic signed [21:0] O18_N4_S2;		always @(posedge clk) O18_N4_S2 <=     O18_N8_S1  +  O18_N10_S1 ;
 logic signed [21:0] O18_N6_S2;		always @(posedge clk) O18_N6_S2 <=     O18_N12_S1  +  O18_N14_S1 ;
 logic signed [21:0] O18_N8_S2;		always @(posedge clk) O18_N8_S2 <=     O18_N16_S1  +  O18_N18_S1 ;
 logic signed [21:0] O18_N10_S2;		always @(posedge clk) O18_N10_S2 <=     O18_N20_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O18_N0_S3;		always @(posedge clk) O18_N0_S3 <=     O18_N0_S2  +  O18_N2_S2 ;
 logic signed [22:0] O18_N2_S3;		always @(posedge clk) O18_N2_S3 <=     O18_N4_S2  +  O18_N6_S2 ;
 logic signed [22:0] O18_N4_S3;		always @(posedge clk) O18_N4_S3 <=     O18_N8_S2  +  O18_N10_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O18_N0_S4;		always @(posedge clk) O18_N0_S4 <=     O18_N0_S3  +  O18_N2_S3 ;
 logic signed [23:0] O18_N2_S4;		always @(posedge clk) O18_N2_S4 <=     O18_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O18_N0_S5;		always @(posedge clk) O18_N0_S5 <=     O18_N0_S4  +  O18_N2_S4 ;
 assign conv_mac_18 = O18_N0_S5;

logic signed [31:0] conv_mac_19;
logic signed [63:0] chainout_0_O19; 
logic signed [63:0] O19_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O19(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay( 9'sd2),.bx(input_fmap_2[7:0]),.by( 9'sd1),.cx(input_fmap_4[7:0]),.cy(-9'sd2),.dx(input_fmap_7[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O19_N0_S1),.chainout(chainout_0_O19));
logic signed [63:0] chainout_2_O19; 
logic signed [63:0] O19_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O19(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_8[7:0]),.ay(-9'sd1),.bx(input_fmap_9[7:0]),.by( 9'sd1),.cx(input_fmap_12[7:0]),.cy( 9'sd1),.dx(input_fmap_16[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O19_N2_S1),.chainout(chainout_2_O19));
logic signed [63:0] chainout_4_O19; 
logic signed [63:0] O19_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O19(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_18[7:0]),.ay(-9'sd1),.bx(input_fmap_21[7:0]),.by( 9'sd1),.cx(input_fmap_24[7:0]),.cy(-9'sd1),.dx(input_fmap_27[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O19_N4_S1),.chainout(chainout_4_O19));
logic signed [63:0] chainout_6_O19; 
logic signed [63:0] O19_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O19(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_34[7:0]),.ay(-9'sd1),.bx(input_fmap_35[7:0]),.by(-9'sd1),.cx(input_fmap_37[7:0]),.cy(-9'sd1),.dx(input_fmap_39[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O19_N6_S1),.chainout(chainout_6_O19));
logic signed [63:0] chainout_8_O19; 
logic signed [63:0] O19_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O19(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_40[7:0]),.ay( 9'sd1),.bx(input_fmap_48[7:0]),.by(-9'sd1),.cx(input_fmap_52[7:0]),.cy( 9'sd1),.dx(input_fmap_53[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O19_N8_S1),.chainout(chainout_8_O19));
logic signed [63:0] chainout_10_O19; 
logic signed [63:0] O19_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O19(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_59[7:0]),.ay(-9'sd2),.bx(input_fmap_61[7:0]),.by( 9'sd1),.cx(input_fmap_62[7:0]),.cy( 9'sd1),.dx(input_fmap_63[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O19_N10_S1),.chainout(chainout_10_O19));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O19_N0_S2;		always @(posedge clk) O19_N0_S2 <=     O19_N0_S1  +  O19_N2_S1 ;
 logic signed [21:0] O19_N2_S2;		always @(posedge clk) O19_N2_S2 <=     O19_N4_S1  +  O19_N6_S1 ;
 logic signed [21:0] O19_N4_S2;		always @(posedge clk) O19_N4_S2 <=     O19_N8_S1  +  O19_N10_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O19_N0_S3;		always @(posedge clk) O19_N0_S3 <=     O19_N0_S2  +  O19_N2_S2 ;
 logic signed [22:0] O19_N2_S3;		always @(posedge clk) O19_N2_S3 <=     O19_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O19_N0_S4;		always @(posedge clk) O19_N0_S4 <=     O19_N0_S3  +  O19_N2_S3 ;
 assign conv_mac_19 = O19_N0_S4;

logic signed [31:0] conv_mac_20;
logic signed [63:0] chainout_0_O20; 
logic signed [63:0] O20_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O20(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay(-9'sd1),.bx(input_fmap_2[7:0]),.by( 9'sd1),.cx(input_fmap_3[7:0]),.cy( 9'sd1),.dx(input_fmap_5[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O20_N0_S1),.chainout(chainout_0_O20));
logic signed [63:0] chainout_2_O20; 
logic signed [63:0] O20_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O20(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_7[7:0]),.ay( 9'sd1),.bx(input_fmap_8[7:0]),.by( 9'sd1),.cx(input_fmap_9[7:0]),.cy( 9'sd3),.dx(input_fmap_11[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O20_N2_S1),.chainout(chainout_2_O20));
logic signed [63:0] chainout_4_O20; 
logic signed [63:0] O20_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O20(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_14[7:0]),.ay( 9'sd1),.bx(input_fmap_15[7:0]),.by(-9'sd1),.cx(input_fmap_16[7:0]),.cy( 9'sd1),.dx(input_fmap_19[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O20_N4_S1),.chainout(chainout_4_O20));
logic signed [63:0] chainout_6_O20; 
logic signed [63:0] O20_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O20(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_20[7:0]),.ay( 9'sd1),.bx(input_fmap_21[7:0]),.by( 9'sd1),.cx(input_fmap_23[7:0]),.cy(-9'sd1),.dx(input_fmap_25[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O20_N6_S1),.chainout(chainout_6_O20));
logic signed [63:0] chainout_8_O20; 
logic signed [63:0] O20_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O20(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_27[7:0]),.ay(-9'sd1),.bx(input_fmap_28[7:0]),.by(-9'sd2),.cx(input_fmap_29[7:0]),.cy(-9'sd1),.dx(input_fmap_30[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O20_N8_S1),.chainout(chainout_8_O20));
logic signed [63:0] chainout_10_O20; 
logic signed [63:0] O20_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O20(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_32[7:0]),.ay( 9'sd1),.bx(input_fmap_33[7:0]),.by( 9'sd2),.cx(input_fmap_34[7:0]),.cy(-9'sd1),.dx(input_fmap_35[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O20_N10_S1),.chainout(chainout_10_O20));
logic signed [63:0] chainout_12_O20; 
logic signed [63:0] O20_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O20(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_38[7:0]),.ay( 9'sd2),.bx(input_fmap_40[7:0]),.by( 9'sd1),.cx(input_fmap_42[7:0]),.cy( 9'sd2),.dx(input_fmap_43[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O20_N12_S1),.chainout(chainout_12_O20));
logic signed [63:0] chainout_14_O20; 
logic signed [63:0] O20_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O20(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_45[7:0]),.ay(-9'sd1),.bx(input_fmap_46[7:0]),.by( 9'sd1),.cx(input_fmap_47[7:0]),.cy(-9'sd1),.dx(input_fmap_50[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O20_N14_S1),.chainout(chainout_14_O20));
logic signed [63:0] chainout_16_O20; 
logic signed [63:0] O20_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O20(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_52[7:0]),.ay(-9'sd2),.bx(input_fmap_53[7:0]),.by( 9'sd2),.cx(input_fmap_54[7:0]),.cy(-9'sd1),.dx(input_fmap_56[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O20_N16_S1),.chainout(chainout_16_O20));
logic signed [63:0] chainout_18_O20; 
logic signed [63:0] O20_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O20(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_57[7:0]),.ay( 9'sd1),.bx(input_fmap_58[7:0]),.by(-9'sd1),.cx(input_fmap_59[7:0]),.cy( 9'sd1),.dx(input_fmap_61[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O20_N18_S1),.chainout(chainout_18_O20));
logic signed [63:0] chainout_20_O20; 
logic signed [63:0] O20_N20_S1; 
 int_sop_4_wrapper int_sop_4_inst_20_O20(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_62[7:0]),.ay( 9'sd2),.bx(input_fmap_63[7:0]),.by(-9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O20_N20_S1),.chainout(chainout_20_O20));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O20_N0_S2;		always @(posedge clk) O20_N0_S2 <=     O20_N0_S1  +  O20_N2_S1 ;
 logic signed [21:0] O20_N2_S2;		always @(posedge clk) O20_N2_S2 <=     O20_N4_S1  +  O20_N6_S1 ;
 logic signed [21:0] O20_N4_S2;		always @(posedge clk) O20_N4_S2 <=     O20_N8_S1  +  O20_N10_S1 ;
 logic signed [21:0] O20_N6_S2;		always @(posedge clk) O20_N6_S2 <=     O20_N12_S1  +  O20_N14_S1 ;
 logic signed [21:0] O20_N8_S2;		always @(posedge clk) O20_N8_S2 <=     O20_N16_S1  +  O20_N18_S1 ;
 logic signed [21:0] O20_N10_S2;		always @(posedge clk) O20_N10_S2 <=     O20_N20_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O20_N0_S3;		always @(posedge clk) O20_N0_S3 <=     O20_N0_S2  +  O20_N2_S2 ;
 logic signed [22:0] O20_N2_S3;		always @(posedge clk) O20_N2_S3 <=     O20_N4_S2  +  O20_N6_S2 ;
 logic signed [22:0] O20_N4_S3;		always @(posedge clk) O20_N4_S3 <=     O20_N8_S2  +  O20_N10_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O20_N0_S4;		always @(posedge clk) O20_N0_S4 <=     O20_N0_S3  +  O20_N2_S3 ;
 logic signed [23:0] O20_N2_S4;		always @(posedge clk) O20_N2_S4 <=     O20_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O20_N0_S5;		always @(posedge clk) O20_N0_S5 <=     O20_N0_S4  +  O20_N2_S4 ;
 assign conv_mac_20 = O20_N0_S5;

logic signed [31:0] conv_mac_21;
logic signed [63:0] chainout_0_O21; 
logic signed [63:0] O21_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O21(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd1),.bx(input_fmap_2[7:0]),.by(-9'sd1),.cx(input_fmap_3[7:0]),.cy( 9'sd1),.dx(input_fmap_4[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O21_N0_S1),.chainout(chainout_0_O21));
logic signed [63:0] chainout_2_O21; 
logic signed [63:0] O21_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O21(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_5[7:0]),.ay( 9'sd1),.bx(input_fmap_8[7:0]),.by(-9'sd1),.cx(input_fmap_9[7:0]),.cy( 9'sd1),.dx(input_fmap_10[7:0]),.dy(-9'sd3),.chainin(63'd0),.result(O21_N2_S1),.chainout(chainout_2_O21));
logic signed [63:0] chainout_4_O21; 
logic signed [63:0] O21_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O21(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_11[7:0]),.ay( 9'sd1),.bx(input_fmap_12[7:0]),.by(-9'sd4),.cx(input_fmap_13[7:0]),.cy(-9'sd1),.dx(input_fmap_14[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O21_N4_S1),.chainout(chainout_4_O21));
logic signed [63:0] chainout_6_O21; 
logic signed [63:0] O21_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O21(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_15[7:0]),.ay(-9'sd1),.bx(input_fmap_17[7:0]),.by(-9'sd1),.cx(input_fmap_18[7:0]),.cy(-9'sd1),.dx(input_fmap_19[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O21_N6_S1),.chainout(chainout_6_O21));
logic signed [63:0] chainout_8_O21; 
logic signed [63:0] O21_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O21(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_20[7:0]),.ay( 9'sd1),.bx(input_fmap_21[7:0]),.by(-9'sd1),.cx(input_fmap_22[7:0]),.cy( 9'sd2),.dx(input_fmap_24[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O21_N8_S1),.chainout(chainout_8_O21));
logic signed [63:0] chainout_10_O21; 
logic signed [63:0] O21_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O21(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_25[7:0]),.ay( 9'sd1),.bx(input_fmap_26[7:0]),.by( 9'sd1),.cx(input_fmap_28[7:0]),.cy( 9'sd1),.dx(input_fmap_29[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O21_N10_S1),.chainout(chainout_10_O21));
logic signed [63:0] chainout_12_O21; 
logic signed [63:0] O21_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O21(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_31[7:0]),.ay( 9'sd3),.bx(input_fmap_33[7:0]),.by(-9'sd2),.cx(input_fmap_34[7:0]),.cy(-9'sd1),.dx(input_fmap_35[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O21_N12_S1),.chainout(chainout_12_O21));
logic signed [63:0] chainout_14_O21; 
logic signed [63:0] O21_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O21(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_36[7:0]),.ay( 9'sd1),.bx(input_fmap_37[7:0]),.by(-9'sd1),.cx(input_fmap_38[7:0]),.cy( 9'sd2),.dx(input_fmap_40[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O21_N14_S1),.chainout(chainout_14_O21));
logic signed [63:0] chainout_16_O21; 
logic signed [63:0] O21_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O21(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_41[7:0]),.ay(-9'sd1),.bx(input_fmap_44[7:0]),.by( 9'sd1),.cx(input_fmap_45[7:0]),.cy( 9'sd1),.dx(input_fmap_46[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O21_N16_S1),.chainout(chainout_16_O21));
logic signed [63:0] chainout_18_O21; 
logic signed [63:0] O21_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O21(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_47[7:0]),.ay( 9'sd1),.bx(input_fmap_48[7:0]),.by( 9'sd1),.cx(input_fmap_50[7:0]),.cy( 9'sd2),.dx(input_fmap_54[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O21_N18_S1),.chainout(chainout_18_O21));
logic signed [63:0] chainout_20_O21; 
logic signed [63:0] O21_N20_S1; 
 int_sop_4_wrapper int_sop_4_inst_20_O21(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_56[7:0]),.ay( 9'sd2),.bx(input_fmap_57[7:0]),.by(-9'sd1),.cx(input_fmap_59[7:0]),.cy(-9'sd1),.dx(input_fmap_60[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O21_N20_S1),.chainout(chainout_20_O21));
logic signed [63:0] chainout_22_O21; 
logic signed [63:0] O21_N22_S1; 
 int_sop_4_wrapper int_sop_4_inst_22_O21(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_63[7:0]),.ay(-9'sd3),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O21_N22_S1),.chainout(chainout_22_O21));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O21_N0_S2;		always @(posedge clk) O21_N0_S2 <=     O21_N0_S1  +  O21_N2_S1 ;
 logic signed [21:0] O21_N2_S2;		always @(posedge clk) O21_N2_S2 <=     O21_N4_S1  +  O21_N6_S1 ;
 logic signed [21:0] O21_N4_S2;		always @(posedge clk) O21_N4_S2 <=     O21_N8_S1  +  O21_N10_S1 ;
 logic signed [21:0] O21_N6_S2;		always @(posedge clk) O21_N6_S2 <=     O21_N12_S1  +  O21_N14_S1 ;
 logic signed [21:0] O21_N8_S2;		always @(posedge clk) O21_N8_S2 <=     O21_N16_S1  +  O21_N18_S1 ;
 logic signed [21:0] O21_N10_S2;		always @(posedge clk) O21_N10_S2 <=     O21_N20_S1  +  O21_N22_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O21_N0_S3;		always @(posedge clk) O21_N0_S3 <=     O21_N0_S2  +  O21_N2_S2 ;
 logic signed [22:0] O21_N2_S3;		always @(posedge clk) O21_N2_S3 <=     O21_N4_S2  +  O21_N6_S2 ;
 logic signed [22:0] O21_N4_S3;		always @(posedge clk) O21_N4_S3 <=     O21_N8_S2  +  O21_N10_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O21_N0_S4;		always @(posedge clk) O21_N0_S4 <=     O21_N0_S3  +  O21_N2_S3 ;
 logic signed [23:0] O21_N2_S4;		always @(posedge clk) O21_N2_S4 <=     O21_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O21_N0_S5;		always @(posedge clk) O21_N0_S5 <=     O21_N0_S4  +  O21_N2_S4 ;
 assign conv_mac_21 = O21_N0_S5;

logic signed [31:0] conv_mac_22;
logic signed [63:0] chainout_0_O22; 
logic signed [63:0] O22_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O22(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd1),.bx(input_fmap_1[7:0]),.by( 9'sd1),.cx(input_fmap_5[7:0]),.cy(-9'sd1),.dx(input_fmap_6[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O22_N0_S1),.chainout(chainout_0_O22));
logic signed [63:0] chainout_2_O22; 
logic signed [63:0] O22_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O22(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_10[7:0]),.ay( 9'sd1),.bx(input_fmap_12[7:0]),.by( 9'sd1),.cx(input_fmap_14[7:0]),.cy( 9'sd1),.dx(input_fmap_15[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O22_N2_S1),.chainout(chainout_2_O22));
logic signed [63:0] chainout_4_O22; 
logic signed [63:0] O22_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O22(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_16[7:0]),.ay(-9'sd1),.bx(input_fmap_17[7:0]),.by(-9'sd1),.cx(input_fmap_18[7:0]),.cy( 9'sd2),.dx(input_fmap_21[7:0]),.dy( 9'sd3),.chainin(63'd0),.result(O22_N4_S1),.chainout(chainout_4_O22));
logic signed [63:0] chainout_6_O22; 
logic signed [63:0] O22_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O22(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_24[7:0]),.ay( 9'sd1),.bx(input_fmap_25[7:0]),.by(-9'sd1),.cx(input_fmap_26[7:0]),.cy(-9'sd1),.dx(input_fmap_28[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O22_N6_S1),.chainout(chainout_6_O22));
logic signed [63:0] chainout_8_O22; 
logic signed [63:0] O22_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O22(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_29[7:0]),.ay( 9'sd1),.bx(input_fmap_30[7:0]),.by( 9'sd1),.cx(input_fmap_31[7:0]),.cy(-9'sd1),.dx(input_fmap_33[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O22_N8_S1),.chainout(chainout_8_O22));
logic signed [63:0] chainout_10_O22; 
logic signed [63:0] O22_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O22(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_35[7:0]),.ay(-9'sd1),.bx(input_fmap_36[7:0]),.by(-9'sd1),.cx(input_fmap_37[7:0]),.cy(-9'sd1),.dx(input_fmap_39[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O22_N10_S1),.chainout(chainout_10_O22));
logic signed [63:0] chainout_12_O22; 
logic signed [63:0] O22_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O22(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_41[7:0]),.ay( 9'sd1),.bx(input_fmap_42[7:0]),.by( 9'sd1),.cx(input_fmap_45[7:0]),.cy(-9'sd1),.dx(input_fmap_46[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O22_N12_S1),.chainout(chainout_12_O22));
logic signed [63:0] chainout_14_O22; 
logic signed [63:0] O22_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O22(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_47[7:0]),.ay(-9'sd1),.bx(input_fmap_50[7:0]),.by(-9'sd1),.cx(input_fmap_51[7:0]),.cy(-9'sd2),.dx(input_fmap_56[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O22_N14_S1),.chainout(chainout_14_O22));
logic signed [63:0] chainout_16_O22; 
logic signed [63:0] O22_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O22(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_57[7:0]),.ay( 9'sd1),.bx(input_fmap_58[7:0]),.by( 9'sd1),.cx(input_fmap_61[7:0]),.cy( 9'sd2),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O22_N16_S1),.chainout(chainout_16_O22));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O22_N0_S2;		always @(posedge clk) O22_N0_S2 <=     O22_N0_S1  +  O22_N2_S1 ;
 logic signed [21:0] O22_N2_S2;		always @(posedge clk) O22_N2_S2 <=     O22_N4_S1  +  O22_N6_S1 ;
 logic signed [21:0] O22_N4_S2;		always @(posedge clk) O22_N4_S2 <=     O22_N8_S1  +  O22_N10_S1 ;
 logic signed [21:0] O22_N6_S2;		always @(posedge clk) O22_N6_S2 <=     O22_N12_S1  +  O22_N14_S1 ;
 logic signed [21:0] O22_N8_S2;		always @(posedge clk) O22_N8_S2 <=     O22_N16_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O22_N0_S3;		always @(posedge clk) O22_N0_S3 <=     O22_N0_S2  +  O22_N2_S2 ;
 logic signed [22:0] O22_N2_S3;		always @(posedge clk) O22_N2_S3 <=     O22_N4_S2  +  O22_N6_S2 ;
 logic signed [22:0] O22_N4_S3;		always @(posedge clk) O22_N4_S3 <=     O22_N8_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O22_N0_S4;		always @(posedge clk) O22_N0_S4 <=     O22_N0_S3  +  O22_N2_S3 ;
 logic signed [23:0] O22_N2_S4;		always @(posedge clk) O22_N2_S4 <=     O22_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O22_N0_S5;		always @(posedge clk) O22_N0_S5 <=     O22_N0_S4  +  O22_N2_S4 ;
 assign conv_mac_22 = O22_N0_S5;

logic signed [31:0] conv_mac_23;
logic signed [63:0] chainout_0_O23; 
logic signed [63:0] O23_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O23(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay( 9'sd2),.bx(input_fmap_2[7:0]),.by( 9'sd1),.cx(input_fmap_3[7:0]),.cy(-9'sd1),.dx(input_fmap_4[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O23_N0_S1),.chainout(chainout_0_O23));
logic signed [63:0] chainout_2_O23; 
logic signed [63:0] O23_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O23(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_6[7:0]),.ay(-9'sd1),.bx(input_fmap_7[7:0]),.by(-9'sd1),.cx(input_fmap_10[7:0]),.cy( 9'sd1),.dx(input_fmap_12[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O23_N2_S1),.chainout(chainout_2_O23));
logic signed [63:0] chainout_4_O23; 
logic signed [63:0] O23_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O23(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_14[7:0]),.ay(-9'sd1),.bx(input_fmap_15[7:0]),.by(-9'sd1),.cx(input_fmap_16[7:0]),.cy( 9'sd1),.dx(input_fmap_19[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O23_N4_S1),.chainout(chainout_4_O23));
logic signed [63:0] chainout_6_O23; 
logic signed [63:0] O23_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O23(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_23[7:0]),.ay( 9'sd1),.bx(input_fmap_25[7:0]),.by( 9'sd1),.cx(input_fmap_29[7:0]),.cy(-9'sd1),.dx(input_fmap_30[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O23_N6_S1),.chainout(chainout_6_O23));
logic signed [63:0] chainout_8_O23; 
logic signed [63:0] O23_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O23(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_34[7:0]),.ay( 9'sd1),.bx(input_fmap_37[7:0]),.by(-9'sd1),.cx(input_fmap_39[7:0]),.cy(-9'sd1),.dx(input_fmap_40[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O23_N8_S1),.chainout(chainout_8_O23));
logic signed [63:0] chainout_10_O23; 
logic signed [63:0] O23_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O23(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_41[7:0]),.ay(-9'sd1),.bx(input_fmap_44[7:0]),.by(-9'sd1),.cx(input_fmap_45[7:0]),.cy( 9'sd1),.dx(input_fmap_48[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O23_N10_S1),.chainout(chainout_10_O23));
logic signed [63:0] chainout_12_O23; 
logic signed [63:0] O23_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O23(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_50[7:0]),.ay( 9'sd1),.bx(input_fmap_52[7:0]),.by(-9'sd1),.cx(input_fmap_53[7:0]),.cy( 9'sd1),.dx(input_fmap_56[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O23_N12_S1),.chainout(chainout_12_O23));
logic signed [63:0] chainout_14_O23; 
logic signed [63:0] O23_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O23(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_57[7:0]),.ay( 9'sd1),.bx(input_fmap_58[7:0]),.by(-9'sd1),.cx(input_fmap_59[7:0]),.cy(-9'sd1),.dx(input_fmap_61[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O23_N14_S1),.chainout(chainout_14_O23));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O23_N0_S2;		always @(posedge clk) O23_N0_S2 <=     O23_N0_S1  +  O23_N2_S1 ;
 logic signed [21:0] O23_N2_S2;		always @(posedge clk) O23_N2_S2 <=     O23_N4_S1  +  O23_N6_S1 ;
 logic signed [21:0] O23_N4_S2;		always @(posedge clk) O23_N4_S2 <=     O23_N8_S1  +  O23_N10_S1 ;
 logic signed [21:0] O23_N6_S2;		always @(posedge clk) O23_N6_S2 <=     O23_N12_S1  +  O23_N14_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O23_N0_S3;		always @(posedge clk) O23_N0_S3 <=     O23_N0_S2  +  O23_N2_S2 ;
 logic signed [22:0] O23_N2_S3;		always @(posedge clk) O23_N2_S3 <=     O23_N4_S2  +  O23_N6_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O23_N0_S4;		always @(posedge clk) O23_N0_S4 <=     O23_N0_S3  +  O23_N2_S3 ;
 assign conv_mac_23 = O23_N0_S4;

logic signed [31:0] conv_mac_24;
logic signed [63:0] chainout_0_O24; 
logic signed [63:0] O24_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O24(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_5[7:0]),.ay( 9'sd1),.bx(input_fmap_7[7:0]),.by( 9'sd1),.cx(input_fmap_10[7:0]),.cy( 9'sd1),.dx(input_fmap_15[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O24_N0_S1),.chainout(chainout_0_O24));
logic signed [63:0] chainout_2_O24; 
logic signed [63:0] O24_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O24(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_16[7:0]),.ay( 9'sd1),.bx(input_fmap_18[7:0]),.by( 9'sd2),.cx(input_fmap_21[7:0]),.cy( 9'sd1),.dx(input_fmap_24[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O24_N2_S1),.chainout(chainout_2_O24));
logic signed [63:0] chainout_4_O24; 
logic signed [63:0] O24_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O24(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_26[7:0]),.ay( 9'sd1),.bx(input_fmap_31[7:0]),.by( 9'sd1),.cx(input_fmap_34[7:0]),.cy(-9'sd1),.dx(input_fmap_35[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O24_N4_S1),.chainout(chainout_4_O24));
logic signed [63:0] chainout_6_O24; 
logic signed [63:0] O24_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O24(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_41[7:0]),.ay( 9'sd1),.bx(input_fmap_45[7:0]),.by(-9'sd1),.cx(input_fmap_59[7:0]),.cy(-9'sd1),.dx(input_fmap_61[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O24_N6_S1),.chainout(chainout_6_O24));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O24_N0_S2;		always @(posedge clk) O24_N0_S2 <=     O24_N0_S1  +  O24_N2_S1 ;
 logic signed [21:0] O24_N2_S2;		always @(posedge clk) O24_N2_S2 <=     O24_N4_S1  +  O24_N6_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O24_N0_S3;		always @(posedge clk) O24_N0_S3 <=     O24_N0_S2  +  O24_N2_S2 ;
 assign conv_mac_24 = O24_N0_S3;

logic signed [31:0] conv_mac_25;
logic signed [63:0] chainout_0_O25; 
logic signed [63:0] O25_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O25(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd1),.bx(input_fmap_1[7:0]),.by(-9'sd1),.cx(input_fmap_2[7:0]),.cy(-9'sd2),.dx(input_fmap_5[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O25_N0_S1),.chainout(chainout_0_O25));
logic signed [63:0] chainout_2_O25; 
logic signed [63:0] O25_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O25(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_6[7:0]),.ay(-9'sd2),.bx(input_fmap_8[7:0]),.by(-9'sd3),.cx(input_fmap_9[7:0]),.cy( 9'sd5),.dx(input_fmap_10[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O25_N2_S1),.chainout(chainout_2_O25));
logic signed [63:0] chainout_4_O25; 
logic signed [63:0] O25_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O25(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_13[7:0]),.ay( 9'sd1),.bx(input_fmap_14[7:0]),.by(-9'sd1),.cx(input_fmap_15[7:0]),.cy( 9'sd1),.dx(input_fmap_17[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O25_N4_S1),.chainout(chainout_4_O25));
logic signed [63:0] chainout_6_O25; 
logic signed [63:0] O25_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O25(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_21[7:0]),.ay(-9'sd1),.bx(input_fmap_23[7:0]),.by(-9'sd1),.cx(input_fmap_25[7:0]),.cy(-9'sd1),.dx(input_fmap_26[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O25_N6_S1),.chainout(chainout_6_O25));
logic signed [63:0] chainout_8_O25; 
logic signed [63:0] O25_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O25(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_27[7:0]),.ay( 9'sd1),.bx(input_fmap_28[7:0]),.by(-9'sd1),.cx(input_fmap_29[7:0]),.cy( 9'sd1),.dx(input_fmap_30[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O25_N8_S1),.chainout(chainout_8_O25));
logic signed [63:0] chainout_10_O25; 
logic signed [63:0] O25_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O25(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_34[7:0]),.ay( 9'sd1),.bx(input_fmap_36[7:0]),.by( 9'sd1),.cx(input_fmap_37[7:0]),.cy(-9'sd3),.dx(input_fmap_41[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O25_N10_S1),.chainout(chainout_10_O25));
logic signed [63:0] chainout_12_O25; 
logic signed [63:0] O25_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O25(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_44[7:0]),.ay( 9'sd1),.bx(input_fmap_46[7:0]),.by(-9'sd2),.cx(input_fmap_47[7:0]),.cy( 9'sd1),.dx(input_fmap_51[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O25_N12_S1),.chainout(chainout_12_O25));
logic signed [63:0] chainout_14_O25; 
logic signed [63:0] O25_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O25(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_52[7:0]),.ay(-9'sd1),.bx(input_fmap_53[7:0]),.by( 9'sd1),.cx(input_fmap_54[7:0]),.cy(-9'sd1),.dx(input_fmap_55[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O25_N14_S1),.chainout(chainout_14_O25));
logic signed [63:0] chainout_16_O25; 
logic signed [63:0] O25_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O25(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_57[7:0]),.ay(-9'sd1),.bx(input_fmap_58[7:0]),.by( 9'sd2),.cx(input_fmap_59[7:0]),.cy(-9'sd1),.dx(input_fmap_63[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O25_N16_S1),.chainout(chainout_16_O25));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O25_N0_S2;		always @(posedge clk) O25_N0_S2 <=     O25_N0_S1  +  O25_N2_S1 ;
 logic signed [21:0] O25_N2_S2;		always @(posedge clk) O25_N2_S2 <=     O25_N4_S1  +  O25_N6_S1 ;
 logic signed [21:0] O25_N4_S2;		always @(posedge clk) O25_N4_S2 <=     O25_N8_S1  +  O25_N10_S1 ;
 logic signed [21:0] O25_N6_S2;		always @(posedge clk) O25_N6_S2 <=     O25_N12_S1  +  O25_N14_S1 ;
 logic signed [21:0] O25_N8_S2;		always @(posedge clk) O25_N8_S2 <=     O25_N16_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O25_N0_S3;		always @(posedge clk) O25_N0_S3 <=     O25_N0_S2  +  O25_N2_S2 ;
 logic signed [22:0] O25_N2_S3;		always @(posedge clk) O25_N2_S3 <=     O25_N4_S2  +  O25_N6_S2 ;
 logic signed [22:0] O25_N4_S3;		always @(posedge clk) O25_N4_S3 <=     O25_N8_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O25_N0_S4;		always @(posedge clk) O25_N0_S4 <=     O25_N0_S3  +  O25_N2_S3 ;
 logic signed [23:0] O25_N2_S4;		always @(posedge clk) O25_N2_S4 <=     O25_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O25_N0_S5;		always @(posedge clk) O25_N0_S5 <=     O25_N0_S4  +  O25_N2_S4 ;
 assign conv_mac_25 = O25_N0_S5;

logic signed [31:0] conv_mac_26;
logic signed [63:0] chainout_0_O26; 
logic signed [63:0] O26_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O26(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay(-9'sd1),.bx(input_fmap_3[7:0]),.by( 9'sd1),.cx(input_fmap_5[7:0]),.cy(-9'sd1),.dx(input_fmap_6[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O26_N0_S1),.chainout(chainout_0_O26));
logic signed [63:0] chainout_2_O26; 
logic signed [63:0] O26_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O26(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_9[7:0]),.ay(-9'sd1),.bx(input_fmap_10[7:0]),.by( 9'sd1),.cx(input_fmap_11[7:0]),.cy( 9'sd2),.dx(input_fmap_12[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O26_N2_S1),.chainout(chainout_2_O26));
logic signed [63:0] chainout_4_O26; 
logic signed [63:0] O26_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O26(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_13[7:0]),.ay(-9'sd1),.bx(input_fmap_14[7:0]),.by( 9'sd1),.cx(input_fmap_16[7:0]),.cy( 9'sd1),.dx(input_fmap_17[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O26_N4_S1),.chainout(chainout_4_O26));
logic signed [63:0] chainout_6_O26; 
logic signed [63:0] O26_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O26(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_20[7:0]),.ay(-9'sd1),.bx(input_fmap_21[7:0]),.by(-9'sd1),.cx(input_fmap_23[7:0]),.cy( 9'sd1),.dx(input_fmap_25[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O26_N6_S1),.chainout(chainout_6_O26));
logic signed [63:0] chainout_8_O26; 
logic signed [63:0] O26_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O26(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_29[7:0]),.ay(-9'sd1),.bx(input_fmap_30[7:0]),.by(-9'sd1),.cx(input_fmap_31[7:0]),.cy(-9'sd1),.dx(input_fmap_34[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O26_N8_S1),.chainout(chainout_8_O26));
logic signed [63:0] chainout_10_O26; 
logic signed [63:0] O26_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O26(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_35[7:0]),.ay(-9'sd2),.bx(input_fmap_39[7:0]),.by( 9'sd2),.cx(input_fmap_40[7:0]),.cy( 9'sd1),.dx(input_fmap_42[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O26_N10_S1),.chainout(chainout_10_O26));
logic signed [63:0] chainout_12_O26; 
logic signed [63:0] O26_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O26(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_43[7:0]),.ay( 9'sd1),.bx(input_fmap_44[7:0]),.by(-9'sd1),.cx(input_fmap_45[7:0]),.cy(-9'sd1),.dx(input_fmap_47[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O26_N12_S1),.chainout(chainout_12_O26));
logic signed [63:0] chainout_14_O26; 
logic signed [63:0] O26_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O26(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_50[7:0]),.ay(-9'sd1),.bx(input_fmap_52[7:0]),.by( 9'sd1),.cx(input_fmap_53[7:0]),.cy( 9'sd1),.dx(input_fmap_56[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O26_N14_S1),.chainout(chainout_14_O26));
logic signed [63:0] chainout_16_O26; 
logic signed [63:0] O26_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O26(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_57[7:0]),.ay(-9'sd1),.bx(input_fmap_60[7:0]),.by( 9'sd1),.cx(input_fmap_61[7:0]),.cy(-9'sd1),.dx(input_fmap_62[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O26_N16_S1),.chainout(chainout_16_O26));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O26_N0_S2;		always @(posedge clk) O26_N0_S2 <=     O26_N0_S1  +  O26_N2_S1 ;
 logic signed [21:0] O26_N2_S2;		always @(posedge clk) O26_N2_S2 <=     O26_N4_S1  +  O26_N6_S1 ;
 logic signed [21:0] O26_N4_S2;		always @(posedge clk) O26_N4_S2 <=     O26_N8_S1  +  O26_N10_S1 ;
 logic signed [21:0] O26_N6_S2;		always @(posedge clk) O26_N6_S2 <=     O26_N12_S1  +  O26_N14_S1 ;
 logic signed [21:0] O26_N8_S2;		always @(posedge clk) O26_N8_S2 <=     O26_N16_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O26_N0_S3;		always @(posedge clk) O26_N0_S3 <=     O26_N0_S2  +  O26_N2_S2 ;
 logic signed [22:0] O26_N2_S3;		always @(posedge clk) O26_N2_S3 <=     O26_N4_S2  +  O26_N6_S2 ;
 logic signed [22:0] O26_N4_S3;		always @(posedge clk) O26_N4_S3 <=     O26_N8_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O26_N0_S4;		always @(posedge clk) O26_N0_S4 <=     O26_N0_S3  +  O26_N2_S3 ;
 logic signed [23:0] O26_N2_S4;		always @(posedge clk) O26_N2_S4 <=     O26_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O26_N0_S5;		always @(posedge clk) O26_N0_S5 <=     O26_N0_S4  +  O26_N2_S4 ;
 assign conv_mac_26 = O26_N0_S5;

logic signed [31:0] conv_mac_27;
logic signed [63:0] chainout_0_O27; 
logic signed [63:0] O27_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O27(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay(-9'sd1),.bx(input_fmap_9[7:0]),.by(-9'sd1),.cx(input_fmap_11[7:0]),.cy( 9'sd1),.dx(input_fmap_24[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O27_N0_S1),.chainout(chainout_0_O27));
logic signed [63:0] chainout_2_O27; 
logic signed [63:0] O27_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O27(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_27[7:0]),.ay( 9'sd1),.bx(input_fmap_28[7:0]),.by( 9'sd1),.cx(input_fmap_32[7:0]),.cy(-9'sd1),.dx(input_fmap_33[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O27_N2_S1),.chainout(chainout_2_O27));
logic signed [63:0] chainout_4_O27; 
logic signed [63:0] O27_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O27(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_38[7:0]),.ay(-9'sd1),.bx(input_fmap_39[7:0]),.by( 9'sd1),.cx(input_fmap_42[7:0]),.cy(-9'sd1),.dx(input_fmap_46[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O27_N4_S1),.chainout(chainout_4_O27));
logic signed [63:0] chainout_6_O27; 
logic signed [63:0] O27_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O27(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_50[7:0]),.ay(-9'sd1),.bx(input_fmap_52[7:0]),.by( 9'sd1),.cx(input_fmap_55[7:0]),.cy(-9'sd1),.dx(input_fmap_57[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O27_N6_S1),.chainout(chainout_6_O27));
logic signed [63:0] chainout_8_O27; 
logic signed [63:0] O27_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O27(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_58[7:0]),.ay(-9'sd1),.bx(input_fmap_61[7:0]),.by( 9'sd1),.cx(input_fmap_63[7:0]),.cy(-9'sd1),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O27_N8_S1),.chainout(chainout_8_O27));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O27_N0_S2;		always @(posedge clk) O27_N0_S2 <=     O27_N0_S1  +  O27_N2_S1 ;
 logic signed [21:0] O27_N2_S2;		always @(posedge clk) O27_N2_S2 <=     O27_N4_S1  +  O27_N6_S1 ;
 logic signed [21:0] O27_N4_S2;		always @(posedge clk) O27_N4_S2 <=     O27_N8_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O27_N0_S3;		always @(posedge clk) O27_N0_S3 <=     O27_N0_S2  +  O27_N2_S2 ;
 logic signed [22:0] O27_N2_S3;		always @(posedge clk) O27_N2_S3 <=     O27_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O27_N0_S4;		always @(posedge clk) O27_N0_S4 <=     O27_N0_S3  +  O27_N2_S3 ;
 assign conv_mac_27 = O27_N0_S4;

logic signed [31:0] conv_mac_28;
logic signed [63:0] chainout_0_O28; 
logic signed [63:0] O28_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O28(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd1),.bx(input_fmap_2[7:0]),.by( 9'sd1),.cx(input_fmap_3[7:0]),.cy( 9'sd1),.dx(input_fmap_4[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O28_N0_S1),.chainout(chainout_0_O28));
logic signed [63:0] chainout_2_O28; 
logic signed [63:0] O28_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O28(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_5[7:0]),.ay( 9'sd2),.bx(input_fmap_6[7:0]),.by(-9'sd1),.cx(input_fmap_7[7:0]),.cy( 9'sd2),.dx(input_fmap_8[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O28_N2_S1),.chainout(chainout_2_O28));
logic signed [63:0] chainout_4_O28; 
logic signed [63:0] O28_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O28(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_11[7:0]),.ay( 9'sd1),.bx(input_fmap_12[7:0]),.by(-9'sd1),.cx(input_fmap_14[7:0]),.cy(-9'sd2),.dx(input_fmap_15[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O28_N4_S1),.chainout(chainout_4_O28));
logic signed [63:0] chainout_6_O28; 
logic signed [63:0] O28_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O28(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_19[7:0]),.ay(-9'sd1),.bx(input_fmap_20[7:0]),.by(-9'sd1),.cx(input_fmap_21[7:0]),.cy(-9'sd1),.dx(input_fmap_23[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O28_N6_S1),.chainout(chainout_6_O28));
logic signed [63:0] chainout_8_O28; 
logic signed [63:0] O28_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O28(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_27[7:0]),.ay(-9'sd1),.bx(input_fmap_28[7:0]),.by( 9'sd2),.cx(input_fmap_29[7:0]),.cy(-9'sd1),.dx(input_fmap_31[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O28_N8_S1),.chainout(chainout_8_O28));
logic signed [63:0] chainout_10_O28; 
logic signed [63:0] O28_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O28(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_33[7:0]),.ay( 9'sd2),.bx(input_fmap_36[7:0]),.by( 9'sd1),.cx(input_fmap_39[7:0]),.cy(-9'sd1),.dx(input_fmap_41[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O28_N10_S1),.chainout(chainout_10_O28));
logic signed [63:0] chainout_12_O28; 
logic signed [63:0] O28_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O28(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_42[7:0]),.ay(-9'sd1),.bx(input_fmap_43[7:0]),.by(-9'sd1),.cx(input_fmap_44[7:0]),.cy( 9'sd1),.dx(input_fmap_45[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O28_N12_S1),.chainout(chainout_12_O28));
logic signed [63:0] chainout_14_O28; 
logic signed [63:0] O28_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O28(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_47[7:0]),.ay(-9'sd2),.bx(input_fmap_48[7:0]),.by(-9'sd1),.cx(input_fmap_49[7:0]),.cy( 9'sd1),.dx(input_fmap_50[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O28_N14_S1),.chainout(chainout_14_O28));
logic signed [63:0] chainout_16_O28; 
logic signed [63:0] O28_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O28(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_51[7:0]),.ay(-9'sd1),.bx(input_fmap_52[7:0]),.by(-9'sd1),.cx(input_fmap_53[7:0]),.cy(-9'sd1),.dx(input_fmap_54[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O28_N16_S1),.chainout(chainout_16_O28));
logic signed [63:0] chainout_18_O28; 
logic signed [63:0] O28_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O28(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_56[7:0]),.ay( 9'sd1),.bx(input_fmap_57[7:0]),.by( 9'sd1),.cx(input_fmap_58[7:0]),.cy(-9'sd1),.dx(input_fmap_59[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O28_N18_S1),.chainout(chainout_18_O28));
logic signed [63:0] chainout_20_O28; 
logic signed [63:0] O28_N20_S1; 
 int_sop_4_wrapper int_sop_4_inst_20_O28(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_60[7:0]),.ay(-9'sd1),.bx(input_fmap_63[7:0]),.by( 9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O28_N20_S1),.chainout(chainout_20_O28));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O28_N0_S2;		always @(posedge clk) O28_N0_S2 <=     O28_N0_S1  +  O28_N2_S1 ;
 logic signed [21:0] O28_N2_S2;		always @(posedge clk) O28_N2_S2 <=     O28_N4_S1  +  O28_N6_S1 ;
 logic signed [21:0] O28_N4_S2;		always @(posedge clk) O28_N4_S2 <=     O28_N8_S1  +  O28_N10_S1 ;
 logic signed [21:0] O28_N6_S2;		always @(posedge clk) O28_N6_S2 <=     O28_N12_S1  +  O28_N14_S1 ;
 logic signed [21:0] O28_N8_S2;		always @(posedge clk) O28_N8_S2 <=     O28_N16_S1  +  O28_N18_S1 ;
 logic signed [21:0] O28_N10_S2;		always @(posedge clk) O28_N10_S2 <=     O28_N20_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O28_N0_S3;		always @(posedge clk) O28_N0_S3 <=     O28_N0_S2  +  O28_N2_S2 ;
 logic signed [22:0] O28_N2_S3;		always @(posedge clk) O28_N2_S3 <=     O28_N4_S2  +  O28_N6_S2 ;
 logic signed [22:0] O28_N4_S3;		always @(posedge clk) O28_N4_S3 <=     O28_N8_S2  +  O28_N10_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O28_N0_S4;		always @(posedge clk) O28_N0_S4 <=     O28_N0_S3  +  O28_N2_S3 ;
 logic signed [23:0] O28_N2_S4;		always @(posedge clk) O28_N2_S4 <=     O28_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O28_N0_S5;		always @(posedge clk) O28_N0_S5 <=     O28_N0_S4  +  O28_N2_S4 ;
 assign conv_mac_28 = O28_N0_S5;

logic signed [31:0] conv_mac_29;
logic signed [63:0] chainout_0_O29; 
logic signed [63:0] O29_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O29(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_2[7:0]),.ay( 9'sd2),.bx(input_fmap_4[7:0]),.by( 9'sd2),.cx(input_fmap_6[7:0]),.cy( 9'sd1),.dx(input_fmap_8[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O29_N0_S1),.chainout(chainout_0_O29));
logic signed [63:0] chainout_2_O29; 
logic signed [63:0] O29_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O29(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_9[7:0]),.ay( 9'sd1),.bx(input_fmap_12[7:0]),.by(-9'sd1),.cx(input_fmap_14[7:0]),.cy( 9'sd1),.dx(input_fmap_16[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O29_N2_S1),.chainout(chainout_2_O29));
logic signed [63:0] chainout_4_O29; 
logic signed [63:0] O29_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O29(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_17[7:0]),.ay(-9'sd1),.bx(input_fmap_18[7:0]),.by( 9'sd5),.cx(input_fmap_19[7:0]),.cy( 9'sd1),.dx(input_fmap_21[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O29_N4_S1),.chainout(chainout_4_O29));
logic signed [63:0] chainout_6_O29; 
logic signed [63:0] O29_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O29(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_22[7:0]),.ay( 9'sd1),.bx(input_fmap_25[7:0]),.by( 9'sd1),.cx(input_fmap_27[7:0]),.cy( 9'sd1),.dx(input_fmap_28[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O29_N6_S1),.chainout(chainout_6_O29));
logic signed [63:0] chainout_8_O29; 
logic signed [63:0] O29_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O29(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_32[7:0]),.ay( 9'sd1),.bx(input_fmap_35[7:0]),.by(-9'sd1),.cx(input_fmap_36[7:0]),.cy(-9'sd1),.dx(input_fmap_40[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O29_N8_S1),.chainout(chainout_8_O29));
logic signed [63:0] chainout_10_O29; 
logic signed [63:0] O29_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O29(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_44[7:0]),.ay(-9'sd1),.bx(input_fmap_48[7:0]),.by(-9'sd1),.cx(input_fmap_49[7:0]),.cy( 9'sd1),.dx(input_fmap_55[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O29_N10_S1),.chainout(chainout_10_O29));
logic signed [63:0] chainout_12_O29; 
logic signed [63:0] O29_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O29(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_58[7:0]),.ay( 9'sd2),.bx(input_fmap_59[7:0]),.by( 9'sd1),.cx(input_fmap_60[7:0]),.cy(-9'sd1),.dx(input_fmap_62[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O29_N12_S1),.chainout(chainout_12_O29));
logic signed [63:0] chainout_14_O29; 
logic signed [63:0] O29_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O29(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_63[7:0]),.ay(-9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O29_N14_S1),.chainout(chainout_14_O29));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O29_N0_S2;		always @(posedge clk) O29_N0_S2 <=     O29_N0_S1  +  O29_N2_S1 ;
 logic signed [21:0] O29_N2_S2;		always @(posedge clk) O29_N2_S2 <=     O29_N4_S1  +  O29_N6_S1 ;
 logic signed [21:0] O29_N4_S2;		always @(posedge clk) O29_N4_S2 <=     O29_N8_S1  +  O29_N10_S1 ;
 logic signed [21:0] O29_N6_S2;		always @(posedge clk) O29_N6_S2 <=     O29_N12_S1  +  O29_N14_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O29_N0_S3;		always @(posedge clk) O29_N0_S3 <=     O29_N0_S2  +  O29_N2_S2 ;
 logic signed [22:0] O29_N2_S3;		always @(posedge clk) O29_N2_S3 <=     O29_N4_S2  +  O29_N6_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O29_N0_S4;		always @(posedge clk) O29_N0_S4 <=     O29_N0_S3  +  O29_N2_S3 ;
 assign conv_mac_29 = O29_N0_S4;

logic signed [31:0] conv_mac_30;
logic signed [63:0] chainout_0_O30; 
logic signed [63:0] O30_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O30(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_3[7:0]),.ay( 9'sd1),.bx(input_fmap_5[7:0]),.by(-9'sd1),.cx(input_fmap_9[7:0]),.cy( 9'sd1),.dx(input_fmap_10[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O30_N0_S1),.chainout(chainout_0_O30));
logic signed [63:0] chainout_2_O30; 
logic signed [63:0] O30_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O30(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_11[7:0]),.ay( 9'sd1),.bx(input_fmap_12[7:0]),.by(-9'sd1),.cx(input_fmap_13[7:0]),.cy(-9'sd1),.dx(input_fmap_15[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O30_N2_S1),.chainout(chainout_2_O30));
logic signed [63:0] chainout_4_O30; 
logic signed [63:0] O30_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O30(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_19[7:0]),.ay( 9'sd2),.bx(input_fmap_22[7:0]),.by( 9'sd1),.cx(input_fmap_25[7:0]),.cy(-9'sd1),.dx(input_fmap_30[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O30_N4_S1),.chainout(chainout_4_O30));
logic signed [63:0] chainout_6_O30; 
logic signed [63:0] O30_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O30(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_32[7:0]),.ay( 9'sd1),.bx(input_fmap_33[7:0]),.by(-9'sd1),.cx(input_fmap_36[7:0]),.cy( 9'sd2),.dx(input_fmap_41[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O30_N6_S1),.chainout(chainout_6_O30));
logic signed [63:0] chainout_8_O30; 
logic signed [63:0] O30_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O30(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_47[7:0]),.ay(-9'sd1),.bx(input_fmap_50[7:0]),.by(-9'sd1),.cx(input_fmap_51[7:0]),.cy(-9'sd1),.dx(input_fmap_54[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O30_N8_S1),.chainout(chainout_8_O30));
logic signed [63:0] chainout_10_O30; 
logic signed [63:0] O30_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O30(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_56[7:0]),.ay(-9'sd1),.bx(input_fmap_59[7:0]),.by(-9'sd1),.cx(input_fmap_61[7:0]),.cy( 9'sd1),.dx(input_fmap_62[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O30_N10_S1),.chainout(chainout_10_O30));
logic signed [63:0] chainout_12_O30; 
logic signed [63:0] O30_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O30(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_63[7:0]),.ay(-9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O30_N12_S1),.chainout(chainout_12_O30));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O30_N0_S2;		always @(posedge clk) O30_N0_S2 <=     O30_N0_S1  +  O30_N2_S1 ;
 logic signed [21:0] O30_N2_S2;		always @(posedge clk) O30_N2_S2 <=     O30_N4_S1  +  O30_N6_S1 ;
 logic signed [21:0] O30_N4_S2;		always @(posedge clk) O30_N4_S2 <=     O30_N8_S1  +  O30_N10_S1 ;
 logic signed [21:0] O30_N6_S2;		always @(posedge clk) O30_N6_S2 <=     O30_N12_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O30_N0_S3;		always @(posedge clk) O30_N0_S3 <=     O30_N0_S2  +  O30_N2_S2 ;
 logic signed [22:0] O30_N2_S3;		always @(posedge clk) O30_N2_S3 <=     O30_N4_S2  +  O30_N6_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O30_N0_S4;		always @(posedge clk) O30_N0_S4 <=     O30_N0_S3  +  O30_N2_S3 ;
 assign conv_mac_30 = O30_N0_S4;

logic signed [31:0] conv_mac_31;
logic signed [63:0] chainout_0_O31; 
logic signed [63:0] O31_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O31(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_3[7:0]),.ay( 9'sd1),.bx(input_fmap_4[7:0]),.by( 9'sd1),.cx(input_fmap_5[7:0]),.cy( 9'sd1),.dx(input_fmap_10[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O31_N0_S1),.chainout(chainout_0_O31));
logic signed [63:0] chainout_2_O31; 
logic signed [63:0] O31_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O31(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_11[7:0]),.ay( 9'sd1),.bx(input_fmap_16[7:0]),.by( 9'sd1),.cx(input_fmap_18[7:0]),.cy( 9'sd1),.dx(input_fmap_19[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O31_N2_S1),.chainout(chainout_2_O31));
logic signed [63:0] chainout_4_O31; 
logic signed [63:0] O31_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O31(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_21[7:0]),.ay(-9'sd1),.bx(input_fmap_27[7:0]),.by(-9'sd1),.cx(input_fmap_29[7:0]),.cy( 9'sd1),.dx(input_fmap_30[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O31_N4_S1),.chainout(chainout_4_O31));
logic signed [63:0] chainout_6_O31; 
logic signed [63:0] O31_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O31(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_31[7:0]),.ay( 9'sd1),.bx(input_fmap_33[7:0]),.by( 9'sd1),.cx(input_fmap_34[7:0]),.cy( 9'sd1),.dx(input_fmap_37[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O31_N6_S1),.chainout(chainout_6_O31));
logic signed [63:0] chainout_8_O31; 
logic signed [63:0] O31_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O31(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_44[7:0]),.ay(-9'sd1),.bx(input_fmap_48[7:0]),.by( 9'sd1),.cx(input_fmap_49[7:0]),.cy( 9'sd1),.dx(input_fmap_50[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O31_N8_S1),.chainout(chainout_8_O31));
logic signed [63:0] chainout_10_O31; 
logic signed [63:0] O31_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O31(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_54[7:0]),.ay(-9'sd1),.bx(input_fmap_55[7:0]),.by( 9'sd1),.cx(input_fmap_57[7:0]),.cy( 9'sd1),.dx(input_fmap_58[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O31_N10_S1),.chainout(chainout_10_O31));
logic signed [63:0] chainout_12_O31; 
logic signed [63:0] O31_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O31(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_59[7:0]),.ay( 9'sd2),.bx(input_fmap_61[7:0]),.by(-9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O31_N12_S1),.chainout(chainout_12_O31));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O31_N0_S2;		always @(posedge clk) O31_N0_S2 <=     O31_N0_S1  +  O31_N2_S1 ;
 logic signed [21:0] O31_N2_S2;		always @(posedge clk) O31_N2_S2 <=     O31_N4_S1  +  O31_N6_S1 ;
 logic signed [21:0] O31_N4_S2;		always @(posedge clk) O31_N4_S2 <=     O31_N8_S1  +  O31_N10_S1 ;
 logic signed [21:0] O31_N6_S2;		always @(posedge clk) O31_N6_S2 <=     O31_N12_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O31_N0_S3;		always @(posedge clk) O31_N0_S3 <=     O31_N0_S2  +  O31_N2_S2 ;
 logic signed [22:0] O31_N2_S3;		always @(posedge clk) O31_N2_S3 <=     O31_N4_S2  +  O31_N6_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O31_N0_S4;		always @(posedge clk) O31_N0_S4 <=     O31_N0_S3  +  O31_N2_S3 ;
 assign conv_mac_31 = O31_N0_S4;

logic signed [31:0] conv_mac_32;
logic signed [63:0] chainout_0_O32; 
logic signed [63:0] O32_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O32(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd1),.bx(input_fmap_2[7:0]),.by(-9'sd2),.cx(input_fmap_4[7:0]),.cy(-9'sd1),.dx(input_fmap_7[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O32_N0_S1),.chainout(chainout_0_O32));
logic signed [63:0] chainout_2_O32; 
logic signed [63:0] O32_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O32(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_8[7:0]),.ay(-9'sd3),.bx(input_fmap_9[7:0]),.by(-9'sd1),.cx(input_fmap_10[7:0]),.cy( 9'sd1),.dx(input_fmap_11[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O32_N2_S1),.chainout(chainout_2_O32));
logic signed [63:0] chainout_4_O32; 
logic signed [63:0] O32_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O32(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_13[7:0]),.ay( 9'sd1),.bx(input_fmap_14[7:0]),.by( 9'sd4),.cx(input_fmap_16[7:0]),.cy(-9'sd1),.dx(input_fmap_17[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O32_N4_S1),.chainout(chainout_4_O32));
logic signed [63:0] chainout_6_O32; 
logic signed [63:0] O32_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O32(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_18[7:0]),.ay(-9'sd1),.bx(input_fmap_21[7:0]),.by(-9'sd2),.cx(input_fmap_22[7:0]),.cy( 9'sd1),.dx(input_fmap_23[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O32_N6_S1),.chainout(chainout_6_O32));
logic signed [63:0] chainout_8_O32; 
logic signed [63:0] O32_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O32(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_25[7:0]),.ay(-9'sd2),.bx(input_fmap_27[7:0]),.by( 9'sd1),.cx(input_fmap_28[7:0]),.cy(-9'sd1),.dx(input_fmap_29[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O32_N8_S1),.chainout(chainout_8_O32));
logic signed [63:0] chainout_10_O32; 
logic signed [63:0] O32_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O32(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_30[7:0]),.ay(-9'sd1),.bx(input_fmap_35[7:0]),.by(-9'sd2),.cx(input_fmap_37[7:0]),.cy( 9'sd1),.dx(input_fmap_38[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O32_N10_S1),.chainout(chainout_10_O32));
logic signed [63:0] chainout_12_O32; 
logic signed [63:0] O32_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O32(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_39[7:0]),.ay(-9'sd1),.bx(input_fmap_40[7:0]),.by(-9'sd1),.cx(input_fmap_41[7:0]),.cy( 9'sd1),.dx(input_fmap_43[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O32_N12_S1),.chainout(chainout_12_O32));
logic signed [63:0] chainout_14_O32; 
logic signed [63:0] O32_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O32(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_44[7:0]),.ay( 9'sd1),.bx(input_fmap_45[7:0]),.by( 9'sd1),.cx(input_fmap_46[7:0]),.cy(-9'sd1),.dx(input_fmap_47[7:0]),.dy( 9'sd3),.chainin(63'd0),.result(O32_N14_S1),.chainout(chainout_14_O32));
logic signed [63:0] chainout_16_O32; 
logic signed [63:0] O32_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O32(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_48[7:0]),.ay(-9'sd1),.bx(input_fmap_49[7:0]),.by( 9'sd2),.cx(input_fmap_50[7:0]),.cy(-9'sd2),.dx(input_fmap_51[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O32_N16_S1),.chainout(chainout_16_O32));
logic signed [63:0] chainout_18_O32; 
logic signed [63:0] O32_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O32(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_52[7:0]),.ay( 9'sd1),.bx(input_fmap_53[7:0]),.by(-9'sd1),.cx(input_fmap_55[7:0]),.cy(-9'sd2),.dx(input_fmap_57[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O32_N18_S1),.chainout(chainout_18_O32));
logic signed [63:0] chainout_20_O32; 
logic signed [63:0] O32_N20_S1; 
 int_sop_4_wrapper int_sop_4_inst_20_O32(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_58[7:0]),.ay( 9'sd2),.bx(input_fmap_59[7:0]),.by( 9'sd3),.cx(input_fmap_61[7:0]),.cy(-9'sd1),.dx(input_fmap_62[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O32_N20_S1),.chainout(chainout_20_O32));
logic signed [63:0] chainout_22_O32; 
logic signed [63:0] O32_N22_S1; 
 int_sop_4_wrapper int_sop_4_inst_22_O32(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_63[7:0]),.ay(-9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O32_N22_S1),.chainout(chainout_22_O32));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O32_N0_S2;		always @(posedge clk) O32_N0_S2 <=     O32_N0_S1  +  O32_N2_S1 ;
 logic signed [21:0] O32_N2_S2;		always @(posedge clk) O32_N2_S2 <=     O32_N4_S1  +  O32_N6_S1 ;
 logic signed [21:0] O32_N4_S2;		always @(posedge clk) O32_N4_S2 <=     O32_N8_S1  +  O32_N10_S1 ;
 logic signed [21:0] O32_N6_S2;		always @(posedge clk) O32_N6_S2 <=     O32_N12_S1  +  O32_N14_S1 ;
 logic signed [21:0] O32_N8_S2;		always @(posedge clk) O32_N8_S2 <=     O32_N16_S1  +  O32_N18_S1 ;
 logic signed [21:0] O32_N10_S2;		always @(posedge clk) O32_N10_S2 <=     O32_N20_S1  +  O32_N22_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O32_N0_S3;		always @(posedge clk) O32_N0_S3 <=     O32_N0_S2  +  O32_N2_S2 ;
 logic signed [22:0] O32_N2_S3;		always @(posedge clk) O32_N2_S3 <=     O32_N4_S2  +  O32_N6_S2 ;
 logic signed [22:0] O32_N4_S3;		always @(posedge clk) O32_N4_S3 <=     O32_N8_S2  +  O32_N10_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O32_N0_S4;		always @(posedge clk) O32_N0_S4 <=     O32_N0_S3  +  O32_N2_S3 ;
 logic signed [23:0] O32_N2_S4;		always @(posedge clk) O32_N2_S4 <=     O32_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O32_N0_S5;		always @(posedge clk) O32_N0_S5 <=     O32_N0_S4  +  O32_N2_S4 ;
 assign conv_mac_32 = O32_N0_S5;

logic signed [31:0] conv_mac_33;
logic signed [63:0] chainout_0_O33; 
logic signed [63:0] O33_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O33(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd1),.bx(input_fmap_1[7:0]),.by(-9'sd1),.cx(input_fmap_3[7:0]),.cy(-9'sd1),.dx(input_fmap_4[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O33_N0_S1),.chainout(chainout_0_O33));
logic signed [63:0] chainout_2_O33; 
logic signed [63:0] O33_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O33(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_6[7:0]),.ay( 9'sd1),.bx(input_fmap_11[7:0]),.by( 9'sd1),.cx(input_fmap_13[7:0]),.cy(-9'sd1),.dx(input_fmap_14[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O33_N2_S1),.chainout(chainout_2_O33));
logic signed [63:0] chainout_4_O33; 
logic signed [63:0] O33_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O33(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_21[7:0]),.ay( 9'sd1),.bx(input_fmap_22[7:0]),.by(-9'sd2),.cx(input_fmap_24[7:0]),.cy(-9'sd2),.dx(input_fmap_26[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O33_N4_S1),.chainout(chainout_4_O33));
logic signed [63:0] chainout_6_O33; 
logic signed [63:0] O33_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O33(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_27[7:0]),.ay(-9'sd1),.bx(input_fmap_31[7:0]),.by(-9'sd2),.cx(input_fmap_33[7:0]),.cy(-9'sd1),.dx(input_fmap_34[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O33_N6_S1),.chainout(chainout_6_O33));
logic signed [63:0] chainout_8_O33; 
logic signed [63:0] O33_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O33(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_35[7:0]),.ay(-9'sd1),.bx(input_fmap_37[7:0]),.by(-9'sd1),.cx(input_fmap_38[7:0]),.cy(-9'sd2),.dx(input_fmap_39[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O33_N8_S1),.chainout(chainout_8_O33));
logic signed [63:0] chainout_10_O33; 
logic signed [63:0] O33_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O33(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_40[7:0]),.ay( 9'sd1),.bx(input_fmap_41[7:0]),.by(-9'sd1),.cx(input_fmap_42[7:0]),.cy( 9'sd2),.dx(input_fmap_43[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O33_N10_S1),.chainout(chainout_10_O33));
logic signed [63:0] chainout_12_O33; 
logic signed [63:0] O33_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O33(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_44[7:0]),.ay( 9'sd1),.bx(input_fmap_45[7:0]),.by( 9'sd1),.cx(input_fmap_46[7:0]),.cy( 9'sd1),.dx(input_fmap_47[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O33_N12_S1),.chainout(chainout_12_O33));
logic signed [63:0] chainout_14_O33; 
logic signed [63:0] O33_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O33(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_49[7:0]),.ay( 9'sd1),.bx(input_fmap_51[7:0]),.by(-9'sd1),.cx(input_fmap_53[7:0]),.cy(-9'sd1),.dx(input_fmap_54[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O33_N14_S1),.chainout(chainout_14_O33));
logic signed [63:0] chainout_16_O33; 
logic signed [63:0] O33_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O33(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_55[7:0]),.ay( 9'sd2),.bx(input_fmap_59[7:0]),.by(-9'sd1),.cx(input_fmap_60[7:0]),.cy(-9'sd1),.dx(input_fmap_61[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O33_N16_S1),.chainout(chainout_16_O33));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O33_N0_S2;		always @(posedge clk) O33_N0_S2 <=     O33_N0_S1  +  O33_N2_S1 ;
 logic signed [21:0] O33_N2_S2;		always @(posedge clk) O33_N2_S2 <=     O33_N4_S1  +  O33_N6_S1 ;
 logic signed [21:0] O33_N4_S2;		always @(posedge clk) O33_N4_S2 <=     O33_N8_S1  +  O33_N10_S1 ;
 logic signed [21:0] O33_N6_S2;		always @(posedge clk) O33_N6_S2 <=     O33_N12_S1  +  O33_N14_S1 ;
 logic signed [21:0] O33_N8_S2;		always @(posedge clk) O33_N8_S2 <=     O33_N16_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O33_N0_S3;		always @(posedge clk) O33_N0_S3 <=     O33_N0_S2  +  O33_N2_S2 ;
 logic signed [22:0] O33_N2_S3;		always @(posedge clk) O33_N2_S3 <=     O33_N4_S2  +  O33_N6_S2 ;
 logic signed [22:0] O33_N4_S3;		always @(posedge clk) O33_N4_S3 <=     O33_N8_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O33_N0_S4;		always @(posedge clk) O33_N0_S4 <=     O33_N0_S3  +  O33_N2_S3 ;
 logic signed [23:0] O33_N2_S4;		always @(posedge clk) O33_N2_S4 <=     O33_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O33_N0_S5;		always @(posedge clk) O33_N0_S5 <=     O33_N0_S4  +  O33_N2_S4 ;
 assign conv_mac_33 = O33_N0_S5;

logic signed [31:0] conv_mac_34;
logic signed [63:0] chainout_0_O34; 
logic signed [63:0] O34_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O34(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd1),.bx(input_fmap_1[7:0]),.by( 9'sd1),.cx(input_fmap_6[7:0]),.cy(-9'sd1),.dx(input_fmap_11[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O34_N0_S1),.chainout(chainout_0_O34));
logic signed [63:0] chainout_2_O34; 
logic signed [63:0] O34_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O34(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_14[7:0]),.ay(-9'sd1),.bx(input_fmap_17[7:0]),.by(-9'sd2),.cx(input_fmap_18[7:0]),.cy( 9'sd1),.dx(input_fmap_19[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O34_N2_S1),.chainout(chainout_2_O34));
logic signed [63:0] chainout_4_O34; 
logic signed [63:0] O34_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O34(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_22[7:0]),.ay( 9'sd1),.bx(input_fmap_23[7:0]),.by(-9'sd1),.cx(input_fmap_25[7:0]),.cy( 9'sd1),.dx(input_fmap_26[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O34_N4_S1),.chainout(chainout_4_O34));
logic signed [63:0] chainout_6_O34; 
logic signed [63:0] O34_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O34(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_29[7:0]),.ay(-9'sd1),.bx(input_fmap_30[7:0]),.by(-9'sd1),.cx(input_fmap_33[7:0]),.cy( 9'sd1),.dx(input_fmap_35[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O34_N6_S1),.chainout(chainout_6_O34));
logic signed [63:0] chainout_8_O34; 
logic signed [63:0] O34_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O34(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_36[7:0]),.ay( 9'sd1),.bx(input_fmap_37[7:0]),.by( 9'sd1),.cx(input_fmap_39[7:0]),.cy(-9'sd2),.dx(input_fmap_40[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O34_N8_S1),.chainout(chainout_8_O34));
logic signed [63:0] chainout_10_O34; 
logic signed [63:0] O34_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O34(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_41[7:0]),.ay(-9'sd1),.bx(input_fmap_42[7:0]),.by(-9'sd2),.cx(input_fmap_43[7:0]),.cy(-9'sd1),.dx(input_fmap_44[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O34_N10_S1),.chainout(chainout_10_O34));
logic signed [63:0] chainout_12_O34; 
logic signed [63:0] O34_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O34(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_45[7:0]),.ay( 9'sd3),.bx(input_fmap_46[7:0]),.by( 9'sd1),.cx(input_fmap_47[7:0]),.cy(-9'sd1),.dx(input_fmap_48[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O34_N12_S1),.chainout(chainout_12_O34));
logic signed [63:0] chainout_14_O34; 
logic signed [63:0] O34_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O34(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_49[7:0]),.ay(-9'sd1),.bx(input_fmap_50[7:0]),.by(-9'sd1),.cx(input_fmap_53[7:0]),.cy( 9'sd1),.dx(input_fmap_57[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O34_N14_S1),.chainout(chainout_14_O34));
logic signed [63:0] chainout_16_O34; 
logic signed [63:0] O34_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O34(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_58[7:0]),.ay( 9'sd2),.bx(input_fmap_59[7:0]),.by( 9'sd1),.cx(input_fmap_62[7:0]),.cy( 9'sd3),.dx(input_fmap_63[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O34_N16_S1),.chainout(chainout_16_O34));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O34_N0_S2;		always @(posedge clk) O34_N0_S2 <=     O34_N0_S1  +  O34_N2_S1 ;
 logic signed [21:0] O34_N2_S2;		always @(posedge clk) O34_N2_S2 <=     O34_N4_S1  +  O34_N6_S1 ;
 logic signed [21:0] O34_N4_S2;		always @(posedge clk) O34_N4_S2 <=     O34_N8_S1  +  O34_N10_S1 ;
 logic signed [21:0] O34_N6_S2;		always @(posedge clk) O34_N6_S2 <=     O34_N12_S1  +  O34_N14_S1 ;
 logic signed [21:0] O34_N8_S2;		always @(posedge clk) O34_N8_S2 <=     O34_N16_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O34_N0_S3;		always @(posedge clk) O34_N0_S3 <=     O34_N0_S2  +  O34_N2_S2 ;
 logic signed [22:0] O34_N2_S3;		always @(posedge clk) O34_N2_S3 <=     O34_N4_S2  +  O34_N6_S2 ;
 logic signed [22:0] O34_N4_S3;		always @(posedge clk) O34_N4_S3 <=     O34_N8_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O34_N0_S4;		always @(posedge clk) O34_N0_S4 <=     O34_N0_S3  +  O34_N2_S3 ;
 logic signed [23:0] O34_N2_S4;		always @(posedge clk) O34_N2_S4 <=     O34_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O34_N0_S5;		always @(posedge clk) O34_N0_S5 <=     O34_N0_S4  +  O34_N2_S4 ;
 assign conv_mac_34 = O34_N0_S5;

logic signed [31:0] conv_mac_35;
logic signed [63:0] chainout_0_O35; 
logic signed [63:0] O35_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O35(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay(-9'sd1),.bx(input_fmap_4[7:0]),.by(-9'sd1),.cx(input_fmap_7[7:0]),.cy(-9'sd1),.dx(input_fmap_8[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O35_N0_S1),.chainout(chainout_0_O35));
logic signed [63:0] chainout_2_O35; 
logic signed [63:0] O35_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O35(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_10[7:0]),.ay(-9'sd1),.bx(input_fmap_11[7:0]),.by( 9'sd1),.cx(input_fmap_13[7:0]),.cy(-9'sd1),.dx(input_fmap_16[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O35_N2_S1),.chainout(chainout_2_O35));
logic signed [63:0] chainout_4_O35; 
logic signed [63:0] O35_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O35(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_18[7:0]),.ay(-9'sd1),.bx(input_fmap_19[7:0]),.by( 9'sd1),.cx(input_fmap_21[7:0]),.cy( 9'sd2),.dx(input_fmap_22[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O35_N4_S1),.chainout(chainout_4_O35));
logic signed [63:0] chainout_6_O35; 
logic signed [63:0] O35_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O35(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_31[7:0]),.ay(-9'sd1),.bx(input_fmap_32[7:0]),.by(-9'sd1),.cx(input_fmap_33[7:0]),.cy(-9'sd1),.dx(input_fmap_35[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O35_N6_S1),.chainout(chainout_6_O35));
logic signed [63:0] chainout_8_O35; 
logic signed [63:0] O35_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O35(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_40[7:0]),.ay( 9'sd1),.bx(input_fmap_42[7:0]),.by( 9'sd2),.cx(input_fmap_48[7:0]),.cy( 9'sd1),.dx(input_fmap_57[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O35_N8_S1),.chainout(chainout_8_O35));
logic signed [63:0] chainout_10_O35; 
logic signed [63:0] O35_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O35(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_58[7:0]),.ay(-9'sd1),.bx(input_fmap_59[7:0]),.by(-9'sd1),.cx(input_fmap_60[7:0]),.cy(-9'sd1),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O35_N10_S1),.chainout(chainout_10_O35));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O35_N0_S2;		always @(posedge clk) O35_N0_S2 <=     O35_N0_S1  +  O35_N2_S1 ;
 logic signed [21:0] O35_N2_S2;		always @(posedge clk) O35_N2_S2 <=     O35_N4_S1  +  O35_N6_S1 ;
 logic signed [21:0] O35_N4_S2;		always @(posedge clk) O35_N4_S2 <=     O35_N8_S1  +  O35_N10_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O35_N0_S3;		always @(posedge clk) O35_N0_S3 <=     O35_N0_S2  +  O35_N2_S2 ;
 logic signed [22:0] O35_N2_S3;		always @(posedge clk) O35_N2_S3 <=     O35_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O35_N0_S4;		always @(posedge clk) O35_N0_S4 <=     O35_N0_S3  +  O35_N2_S3 ;
 assign conv_mac_35 = O35_N0_S4;

logic signed [31:0] conv_mac_36;
logic signed [63:0] chainout_0_O36; 
logic signed [63:0] O36_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O36(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd3),.bx(input_fmap_7[7:0]),.by(-9'sd1),.cx(input_fmap_8[7:0]),.cy( 9'sd1),.dx(input_fmap_10[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O36_N0_S1),.chainout(chainout_0_O36));
logic signed [63:0] chainout_2_O36; 
logic signed [63:0] O36_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O36(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_12[7:0]),.ay(-9'sd1),.bx(input_fmap_13[7:0]),.by(-9'sd1),.cx(input_fmap_16[7:0]),.cy( 9'sd1),.dx(input_fmap_18[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O36_N2_S1),.chainout(chainout_2_O36));
logic signed [63:0] chainout_4_O36; 
logic signed [63:0] O36_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O36(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_19[7:0]),.ay( 9'sd2),.bx(input_fmap_20[7:0]),.by( 9'sd1),.cx(input_fmap_21[7:0]),.cy( 9'sd1),.dx(input_fmap_22[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O36_N4_S1),.chainout(chainout_4_O36));
logic signed [63:0] chainout_6_O36; 
logic signed [63:0] O36_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O36(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_24[7:0]),.ay( 9'sd1),.bx(input_fmap_25[7:0]),.by(-9'sd2),.cx(input_fmap_32[7:0]),.cy( 9'sd1),.dx(input_fmap_33[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O36_N6_S1),.chainout(chainout_6_O36));
logic signed [63:0] chainout_8_O36; 
logic signed [63:0] O36_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O36(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_34[7:0]),.ay( 9'sd1),.bx(input_fmap_35[7:0]),.by(-9'sd1),.cx(input_fmap_37[7:0]),.cy(-9'sd1),.dx(input_fmap_43[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O36_N8_S1),.chainout(chainout_8_O36));
logic signed [63:0] chainout_10_O36; 
logic signed [63:0] O36_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O36(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_44[7:0]),.ay( 9'sd1),.bx(input_fmap_46[7:0]),.by(-9'sd1),.cx(input_fmap_47[7:0]),.cy(-9'sd1),.dx(input_fmap_48[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O36_N10_S1),.chainout(chainout_10_O36));
logic signed [63:0] chainout_12_O36; 
logic signed [63:0] O36_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O36(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_49[7:0]),.ay(-9'sd1),.bx(input_fmap_51[7:0]),.by(-9'sd2),.cx(input_fmap_53[7:0]),.cy( 9'sd1),.dx(input_fmap_55[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O36_N12_S1),.chainout(chainout_12_O36));
logic signed [63:0] chainout_14_O36; 
logic signed [63:0] O36_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O36(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_56[7:0]),.ay( 9'sd1),.bx(input_fmap_57[7:0]),.by(-9'sd1),.cx(input_fmap_58[7:0]),.cy( 9'sd1),.dx(input_fmap_61[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O36_N14_S1),.chainout(chainout_14_O36));
logic signed [63:0] chainout_16_O36; 
logic signed [63:0] O36_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O36(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_62[7:0]),.ay( 9'sd1),.bx(input_fmap_63[7:0]),.by(-9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O36_N16_S1),.chainout(chainout_16_O36));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O36_N0_S2;		always @(posedge clk) O36_N0_S2 <=     O36_N0_S1  +  O36_N2_S1 ;
 logic signed [21:0] O36_N2_S2;		always @(posedge clk) O36_N2_S2 <=     O36_N4_S1  +  O36_N6_S1 ;
 logic signed [21:0] O36_N4_S2;		always @(posedge clk) O36_N4_S2 <=     O36_N8_S1  +  O36_N10_S1 ;
 logic signed [21:0] O36_N6_S2;		always @(posedge clk) O36_N6_S2 <=     O36_N12_S1  +  O36_N14_S1 ;
 logic signed [21:0] O36_N8_S2;		always @(posedge clk) O36_N8_S2 <=     O36_N16_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O36_N0_S3;		always @(posedge clk) O36_N0_S3 <=     O36_N0_S2  +  O36_N2_S2 ;
 logic signed [22:0] O36_N2_S3;		always @(posedge clk) O36_N2_S3 <=     O36_N4_S2  +  O36_N6_S2 ;
 logic signed [22:0] O36_N4_S3;		always @(posedge clk) O36_N4_S3 <=     O36_N8_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O36_N0_S4;		always @(posedge clk) O36_N0_S4 <=     O36_N0_S3  +  O36_N2_S3 ;
 logic signed [23:0] O36_N2_S4;		always @(posedge clk) O36_N2_S4 <=     O36_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O36_N0_S5;		always @(posedge clk) O36_N0_S5 <=     O36_N0_S4  +  O36_N2_S4 ;
 assign conv_mac_36 = O36_N0_S5;

logic signed [31:0] conv_mac_37;
logic signed [63:0] chainout_0_O37; 
logic signed [63:0] O37_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O37(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay(-9'sd1),.bx(input_fmap_2[7:0]),.by(-9'sd1),.cx(input_fmap_5[7:0]),.cy( 9'sd1),.dx(input_fmap_6[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O37_N0_S1),.chainout(chainout_0_O37));
logic signed [63:0] chainout_2_O37; 
logic signed [63:0] O37_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O37(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_11[7:0]),.ay( 9'sd2),.bx(input_fmap_15[7:0]),.by( 9'sd1),.cx(input_fmap_16[7:0]),.cy( 9'sd2),.dx(input_fmap_19[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O37_N2_S1),.chainout(chainout_2_O37));
logic signed [63:0] chainout_4_O37; 
logic signed [63:0] O37_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O37(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_24[7:0]),.ay(-9'sd1),.bx(input_fmap_28[7:0]),.by(-9'sd1),.cx(input_fmap_29[7:0]),.cy( 9'sd1),.dx(input_fmap_30[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O37_N4_S1),.chainout(chainout_4_O37));
logic signed [63:0] chainout_6_O37; 
logic signed [63:0] O37_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O37(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_32[7:0]),.ay( 9'sd1),.bx(input_fmap_33[7:0]),.by( 9'sd1),.cx(input_fmap_34[7:0]),.cy( 9'sd1),.dx(input_fmap_35[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O37_N6_S1),.chainout(chainout_6_O37));
logic signed [63:0] chainout_8_O37; 
logic signed [63:0] O37_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O37(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_38[7:0]),.ay(-9'sd1),.bx(input_fmap_39[7:0]),.by(-9'sd1),.cx(input_fmap_42[7:0]),.cy(-9'sd1),.dx(input_fmap_50[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O37_N8_S1),.chainout(chainout_8_O37));
logic signed [63:0] chainout_10_O37; 
logic signed [63:0] O37_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O37(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_52[7:0]),.ay( 9'sd1),.bx(input_fmap_53[7:0]),.by( 9'sd1),.cx(input_fmap_57[7:0]),.cy( 9'sd2),.dx(input_fmap_59[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O37_N10_S1),.chainout(chainout_10_O37));
logic signed [63:0] chainout_12_O37; 
logic signed [63:0] O37_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O37(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_61[7:0]),.ay(-9'sd2),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O37_N12_S1),.chainout(chainout_12_O37));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O37_N0_S2;		always @(posedge clk) O37_N0_S2 <=     O37_N0_S1  +  O37_N2_S1 ;
 logic signed [21:0] O37_N2_S2;		always @(posedge clk) O37_N2_S2 <=     O37_N4_S1  +  O37_N6_S1 ;
 logic signed [21:0] O37_N4_S2;		always @(posedge clk) O37_N4_S2 <=     O37_N8_S1  +  O37_N10_S1 ;
 logic signed [21:0] O37_N6_S2;		always @(posedge clk) O37_N6_S2 <=     O37_N12_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O37_N0_S3;		always @(posedge clk) O37_N0_S3 <=     O37_N0_S2  +  O37_N2_S2 ;
 logic signed [22:0] O37_N2_S3;		always @(posedge clk) O37_N2_S3 <=     O37_N4_S2  +  O37_N6_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O37_N0_S4;		always @(posedge clk) O37_N0_S4 <=     O37_N0_S3  +  O37_N2_S3 ;
 assign conv_mac_37 = O37_N0_S4;

logic signed [31:0] conv_mac_38;
logic signed [63:0] chainout_0_O38; 
logic signed [63:0] O38_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O38(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay( 9'sd1),.bx(input_fmap_5[7:0]),.by(-9'sd1),.cx(input_fmap_13[7:0]),.cy( 9'sd1),.dx(input_fmap_14[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O38_N0_S1),.chainout(chainout_0_O38));
logic signed [63:0] chainout_2_O38; 
logic signed [63:0] O38_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O38(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_17[7:0]),.ay(-9'sd1),.bx(input_fmap_19[7:0]),.by( 9'sd1),.cx(input_fmap_20[7:0]),.cy( 9'sd1),.dx(input_fmap_21[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O38_N2_S1),.chainout(chainout_2_O38));
logic signed [63:0] chainout_4_O38; 
logic signed [63:0] O38_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O38(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_24[7:0]),.ay( 9'sd1),.bx(input_fmap_27[7:0]),.by(-9'sd1),.cx(input_fmap_28[7:0]),.cy(-9'sd1),.dx(input_fmap_29[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O38_N4_S1),.chainout(chainout_4_O38));
logic signed [63:0] chainout_6_O38; 
logic signed [63:0] O38_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O38(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_31[7:0]),.ay(-9'sd1),.bx(input_fmap_32[7:0]),.by( 9'sd2),.cx(input_fmap_33[7:0]),.cy(-9'sd1),.dx(input_fmap_34[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O38_N6_S1),.chainout(chainout_6_O38));
logic signed [63:0] chainout_8_O38; 
logic signed [63:0] O38_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O38(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_35[7:0]),.ay( 9'sd1),.bx(input_fmap_36[7:0]),.by( 9'sd1),.cx(input_fmap_38[7:0]),.cy(-9'sd1),.dx(input_fmap_40[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O38_N8_S1),.chainout(chainout_8_O38));
logic signed [63:0] chainout_10_O38; 
logic signed [63:0] O38_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O38(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_43[7:0]),.ay( 9'sd1),.bx(input_fmap_45[7:0]),.by(-9'sd1),.cx(input_fmap_47[7:0]),.cy(-9'sd1),.dx(input_fmap_49[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O38_N10_S1),.chainout(chainout_10_O38));
logic signed [63:0] chainout_12_O38; 
logic signed [63:0] O38_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O38(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_50[7:0]),.ay(-9'sd1),.bx(input_fmap_52[7:0]),.by(-9'sd1),.cx(input_fmap_53[7:0]),.cy( 9'sd1),.dx(input_fmap_55[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O38_N12_S1),.chainout(chainout_12_O38));
logic signed [63:0] chainout_14_O38; 
logic signed [63:0] O38_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O38(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_57[7:0]),.ay( 9'sd1),.bx(input_fmap_61[7:0]),.by(-9'sd1),.cx(input_fmap_63[7:0]),.cy(-9'sd1),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O38_N14_S1),.chainout(chainout_14_O38));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O38_N0_S2;		always @(posedge clk) O38_N0_S2 <=     O38_N0_S1  +  O38_N2_S1 ;
 logic signed [21:0] O38_N2_S2;		always @(posedge clk) O38_N2_S2 <=     O38_N4_S1  +  O38_N6_S1 ;
 logic signed [21:0] O38_N4_S2;		always @(posedge clk) O38_N4_S2 <=     O38_N8_S1  +  O38_N10_S1 ;
 logic signed [21:0] O38_N6_S2;		always @(posedge clk) O38_N6_S2 <=     O38_N12_S1  +  O38_N14_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O38_N0_S3;		always @(posedge clk) O38_N0_S3 <=     O38_N0_S2  +  O38_N2_S2 ;
 logic signed [22:0] O38_N2_S3;		always @(posedge clk) O38_N2_S3 <=     O38_N4_S2  +  O38_N6_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O38_N0_S4;		always @(posedge clk) O38_N0_S4 <=     O38_N0_S3  +  O38_N2_S3 ;
 assign conv_mac_38 = O38_N0_S4;

logic signed [31:0] conv_mac_39;
logic signed [63:0] chainout_0_O39; 
logic signed [63:0] O39_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O39(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_2[7:0]),.ay(-9'sd1),.bx(input_fmap_3[7:0]),.by( 9'sd1),.cx(input_fmap_4[7:0]),.cy( 9'sd1),.dx(input_fmap_5[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O39_N0_S1),.chainout(chainout_0_O39));
logic signed [63:0] chainout_2_O39; 
logic signed [63:0] O39_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O39(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_6[7:0]),.ay( 9'sd1),.bx(input_fmap_12[7:0]),.by( 9'sd1),.cx(input_fmap_13[7:0]),.cy( 9'sd1),.dx(input_fmap_15[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O39_N2_S1),.chainout(chainout_2_O39));
logic signed [63:0] chainout_4_O39; 
logic signed [63:0] O39_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O39(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_18[7:0]),.ay( 9'sd1),.bx(input_fmap_19[7:0]),.by( 9'sd1),.cx(input_fmap_22[7:0]),.cy( 9'sd1),.dx(input_fmap_26[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O39_N4_S1),.chainout(chainout_4_O39));
logic signed [63:0] chainout_6_O39; 
logic signed [63:0] O39_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O39(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_29[7:0]),.ay( 9'sd1),.bx(input_fmap_47[7:0]),.by(-9'sd1),.cx(input_fmap_48[7:0]),.cy( 9'sd1),.dx(input_fmap_51[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O39_N6_S1),.chainout(chainout_6_O39));
logic signed [63:0] chainout_8_O39; 
logic signed [63:0] O39_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O39(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_55[7:0]),.ay( 9'sd1),.bx(input_fmap_59[7:0]),.by( 9'sd2),.cx(input_fmap_60[7:0]),.cy(-9'sd1),.dx(input_fmap_62[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O39_N8_S1),.chainout(chainout_8_O39));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O39_N0_S2;		always @(posedge clk) O39_N0_S2 <=     O39_N0_S1  +  O39_N2_S1 ;
 logic signed [21:0] O39_N2_S2;		always @(posedge clk) O39_N2_S2 <=     O39_N4_S1  +  O39_N6_S1 ;
 logic signed [21:0] O39_N4_S2;		always @(posedge clk) O39_N4_S2 <=     O39_N8_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O39_N0_S3;		always @(posedge clk) O39_N0_S3 <=     O39_N0_S2  +  O39_N2_S2 ;
 logic signed [22:0] O39_N2_S3;		always @(posedge clk) O39_N2_S3 <=     O39_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O39_N0_S4;		always @(posedge clk) O39_N0_S4 <=     O39_N0_S3  +  O39_N2_S3 ;
 assign conv_mac_39 = O39_N0_S4;

logic signed [31:0] conv_mac_40;
logic signed [63:0] chainout_0_O40; 
logic signed [63:0] O40_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O40(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay(-9'sd1),.bx(input_fmap_2[7:0]),.by( 9'sd1),.cx(input_fmap_3[7:0]),.cy(-9'sd2),.dx(input_fmap_6[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O40_N0_S1),.chainout(chainout_0_O40));
logic signed [63:0] chainout_2_O40; 
logic signed [63:0] O40_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O40(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_7[7:0]),.ay(-9'sd1),.bx(input_fmap_9[7:0]),.by( 9'sd1),.cx(input_fmap_10[7:0]),.cy(-9'sd1),.dx(input_fmap_11[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O40_N2_S1),.chainout(chainout_2_O40));
logic signed [63:0] chainout_4_O40; 
logic signed [63:0] O40_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O40(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_12[7:0]),.ay( 9'sd2),.bx(input_fmap_15[7:0]),.by( 9'sd3),.cx(input_fmap_16[7:0]),.cy( 9'sd2),.dx(input_fmap_17[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O40_N4_S1),.chainout(chainout_4_O40));
logic signed [63:0] chainout_6_O40; 
logic signed [63:0] O40_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O40(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_19[7:0]),.ay( 9'sd1),.bx(input_fmap_21[7:0]),.by( 9'sd2),.cx(input_fmap_22[7:0]),.cy(-9'sd1),.dx(input_fmap_23[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O40_N6_S1),.chainout(chainout_6_O40));
logic signed [63:0] chainout_8_O40; 
logic signed [63:0] O40_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O40(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_25[7:0]),.ay( 9'sd1),.bx(input_fmap_26[7:0]),.by(-9'sd1),.cx(input_fmap_27[7:0]),.cy( 9'sd1),.dx(input_fmap_28[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O40_N8_S1),.chainout(chainout_8_O40));
logic signed [63:0] chainout_10_O40; 
logic signed [63:0] O40_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O40(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_29[7:0]),.ay(-9'sd2),.bx(input_fmap_30[7:0]),.by(-9'sd1),.cx(input_fmap_31[7:0]),.cy(-9'sd2),.dx(input_fmap_34[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O40_N10_S1),.chainout(chainout_10_O40));
logic signed [63:0] chainout_12_O40; 
logic signed [63:0] O40_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O40(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_35[7:0]),.ay( 9'sd1),.bx(input_fmap_36[7:0]),.by(-9'sd1),.cx(input_fmap_37[7:0]),.cy( 9'sd1),.dx(input_fmap_41[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O40_N12_S1),.chainout(chainout_12_O40));
logic signed [63:0] chainout_14_O40; 
logic signed [63:0] O40_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O40(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_43[7:0]),.ay(-9'sd2),.bx(input_fmap_44[7:0]),.by(-9'sd1),.cx(input_fmap_45[7:0]),.cy(-9'sd1),.dx(input_fmap_47[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O40_N14_S1),.chainout(chainout_14_O40));
logic signed [63:0] chainout_16_O40; 
logic signed [63:0] O40_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O40(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_48[7:0]),.ay(-9'sd1),.bx(input_fmap_50[7:0]),.by(-9'sd1),.cx(input_fmap_51[7:0]),.cy( 9'sd1),.dx(input_fmap_52[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O40_N16_S1),.chainout(chainout_16_O40));
logic signed [63:0] chainout_18_O40; 
logic signed [63:0] O40_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O40(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_54[7:0]),.ay(-9'sd1),.bx(input_fmap_55[7:0]),.by( 9'sd1),.cx(input_fmap_56[7:0]),.cy( 9'sd1),.dx(input_fmap_58[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O40_N18_S1),.chainout(chainout_18_O40));
logic signed [63:0] chainout_20_O40; 
logic signed [63:0] O40_N20_S1; 
 int_sop_4_wrapper int_sop_4_inst_20_O40(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_59[7:0]),.ay( 9'sd1),.bx(input_fmap_60[7:0]),.by(-9'sd1),.cx(input_fmap_61[7:0]),.cy( 9'sd1),.dx(input_fmap_62[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O40_N20_S1),.chainout(chainout_20_O40));
logic signed [63:0] chainout_22_O40; 
logic signed [63:0] O40_N22_S1; 
 int_sop_4_wrapper int_sop_4_inst_22_O40(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_63[7:0]),.ay( 9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O40_N22_S1),.chainout(chainout_22_O40));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O40_N0_S2;		always @(posedge clk) O40_N0_S2 <=     O40_N0_S1  +  O40_N2_S1 ;
 logic signed [21:0] O40_N2_S2;		always @(posedge clk) O40_N2_S2 <=     O40_N4_S1  +  O40_N6_S1 ;
 logic signed [21:0] O40_N4_S2;		always @(posedge clk) O40_N4_S2 <=     O40_N8_S1  +  O40_N10_S1 ;
 logic signed [21:0] O40_N6_S2;		always @(posedge clk) O40_N6_S2 <=     O40_N12_S1  +  O40_N14_S1 ;
 logic signed [21:0] O40_N8_S2;		always @(posedge clk) O40_N8_S2 <=     O40_N16_S1  +  O40_N18_S1 ;
 logic signed [21:0] O40_N10_S2;		always @(posedge clk) O40_N10_S2 <=     O40_N20_S1  +  O40_N22_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O40_N0_S3;		always @(posedge clk) O40_N0_S3 <=     O40_N0_S2  +  O40_N2_S2 ;
 logic signed [22:0] O40_N2_S3;		always @(posedge clk) O40_N2_S3 <=     O40_N4_S2  +  O40_N6_S2 ;
 logic signed [22:0] O40_N4_S3;		always @(posedge clk) O40_N4_S3 <=     O40_N8_S2  +  O40_N10_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O40_N0_S4;		always @(posedge clk) O40_N0_S4 <=     O40_N0_S3  +  O40_N2_S3 ;
 logic signed [23:0] O40_N2_S4;		always @(posedge clk) O40_N2_S4 <=     O40_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O40_N0_S5;		always @(posedge clk) O40_N0_S5 <=     O40_N0_S4  +  O40_N2_S4 ;
 assign conv_mac_40 = O40_N0_S5;

logic signed [31:0] conv_mac_41;
logic signed [63:0] chainout_0_O41; 
logic signed [63:0] O41_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O41(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay(-9'sd1),.bx(input_fmap_9[7:0]),.by(-9'sd2),.cx(input_fmap_12[7:0]),.cy( 9'sd1),.dx(input_fmap_15[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O41_N0_S1),.chainout(chainout_0_O41));
logic signed [63:0] chainout_2_O41; 
logic signed [63:0] O41_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O41(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_19[7:0]),.ay(-9'sd1),.bx(input_fmap_20[7:0]),.by( 9'sd1),.cx(input_fmap_21[7:0]),.cy( 9'sd1),.dx(input_fmap_24[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O41_N2_S1),.chainout(chainout_2_O41));
logic signed [63:0] chainout_4_O41; 
logic signed [63:0] O41_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O41(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_27[7:0]),.ay(-9'sd1),.bx(input_fmap_30[7:0]),.by(-9'sd1),.cx(input_fmap_32[7:0]),.cy( 9'sd2),.dx(input_fmap_34[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O41_N4_S1),.chainout(chainout_4_O41));
logic signed [63:0] chainout_6_O41; 
logic signed [63:0] O41_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O41(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_36[7:0]),.ay( 9'sd2),.bx(input_fmap_37[7:0]),.by( 9'sd1),.cx(input_fmap_38[7:0]),.cy( 9'sd2),.dx(input_fmap_40[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O41_N6_S1),.chainout(chainout_6_O41));
logic signed [63:0] chainout_8_O41; 
logic signed [63:0] O41_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O41(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_44[7:0]),.ay(-9'sd1),.bx(input_fmap_45[7:0]),.by( 9'sd1),.cx(input_fmap_46[7:0]),.cy( 9'sd1),.dx(input_fmap_48[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O41_N8_S1),.chainout(chainout_8_O41));
logic signed [63:0] chainout_10_O41; 
logic signed [63:0] O41_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O41(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_49[7:0]),.ay(-9'sd1),.bx(input_fmap_52[7:0]),.by(-9'sd1),.cx(input_fmap_54[7:0]),.cy( 9'sd1),.dx(input_fmap_55[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O41_N10_S1),.chainout(chainout_10_O41));
logic signed [63:0] chainout_12_O41; 
logic signed [63:0] O41_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O41(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_56[7:0]),.ay( 9'sd1),.bx(input_fmap_57[7:0]),.by(-9'sd1),.cx(input_fmap_58[7:0]),.cy(-9'sd1),.dx(input_fmap_59[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O41_N12_S1),.chainout(chainout_12_O41));
logic signed [63:0] chainout_14_O41; 
logic signed [63:0] O41_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O41(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_60[7:0]),.ay( 9'sd1),.bx(input_fmap_61[7:0]),.by( 9'sd1),.cx(input_fmap_63[7:0]),.cy( 9'sd1),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O41_N14_S1),.chainout(chainout_14_O41));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O41_N0_S2;		always @(posedge clk) O41_N0_S2 <=     O41_N0_S1  +  O41_N2_S1 ;
 logic signed [21:0] O41_N2_S2;		always @(posedge clk) O41_N2_S2 <=     O41_N4_S1  +  O41_N6_S1 ;
 logic signed [21:0] O41_N4_S2;		always @(posedge clk) O41_N4_S2 <=     O41_N8_S1  +  O41_N10_S1 ;
 logic signed [21:0] O41_N6_S2;		always @(posedge clk) O41_N6_S2 <=     O41_N12_S1  +  O41_N14_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O41_N0_S3;		always @(posedge clk) O41_N0_S3 <=     O41_N0_S2  +  O41_N2_S2 ;
 logic signed [22:0] O41_N2_S3;		always @(posedge clk) O41_N2_S3 <=     O41_N4_S2  +  O41_N6_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O41_N0_S4;		always @(posedge clk) O41_N0_S4 <=     O41_N0_S3  +  O41_N2_S3 ;
 assign conv_mac_41 = O41_N0_S4;

logic signed [31:0] conv_mac_42;
logic signed [63:0] chainout_0_O42; 
logic signed [63:0] O42_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O42(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay( 9'sd2),.bx(input_fmap_4[7:0]),.by(-9'sd1),.cx(input_fmap_5[7:0]),.cy(-9'sd1),.dx(input_fmap_6[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O42_N0_S1),.chainout(chainout_0_O42));
logic signed [63:0] chainout_2_O42; 
logic signed [63:0] O42_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O42(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_7[7:0]),.ay(-9'sd1),.bx(input_fmap_8[7:0]),.by(-9'sd1),.cx(input_fmap_9[7:0]),.cy( 9'sd1),.dx(input_fmap_11[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O42_N2_S1),.chainout(chainout_2_O42));
logic signed [63:0] chainout_4_O42; 
logic signed [63:0] O42_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O42(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_12[7:0]),.ay( 9'sd1),.bx(input_fmap_13[7:0]),.by(-9'sd1),.cx(input_fmap_14[7:0]),.cy( 9'sd2),.dx(input_fmap_15[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O42_N4_S1),.chainout(chainout_4_O42));
logic signed [63:0] chainout_6_O42; 
logic signed [63:0] O42_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O42(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_16[7:0]),.ay(-9'sd2),.bx(input_fmap_18[7:0]),.by(-9'sd2),.cx(input_fmap_19[7:0]),.cy( 9'sd1),.dx(input_fmap_22[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O42_N6_S1),.chainout(chainout_6_O42));
logic signed [63:0] chainout_8_O42; 
logic signed [63:0] O42_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O42(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_23[7:0]),.ay( 9'sd1),.bx(input_fmap_25[7:0]),.by(-9'sd1),.cx(input_fmap_28[7:0]),.cy(-9'sd1),.dx(input_fmap_30[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O42_N8_S1),.chainout(chainout_8_O42));
logic signed [63:0] chainout_10_O42; 
logic signed [63:0] O42_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O42(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_31[7:0]),.ay(-9'sd1),.bx(input_fmap_33[7:0]),.by(-9'sd1),.cx(input_fmap_36[7:0]),.cy( 9'sd2),.dx(input_fmap_37[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O42_N10_S1),.chainout(chainout_10_O42));
logic signed [63:0] chainout_12_O42; 
logic signed [63:0] O42_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O42(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_38[7:0]),.ay( 9'sd2),.bx(input_fmap_42[7:0]),.by( 9'sd1),.cx(input_fmap_43[7:0]),.cy(-9'sd1),.dx(input_fmap_44[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O42_N12_S1),.chainout(chainout_12_O42));
logic signed [63:0] chainout_14_O42; 
logic signed [63:0] O42_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O42(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_46[7:0]),.ay( 9'sd1),.bx(input_fmap_48[7:0]),.by(-9'sd1),.cx(input_fmap_52[7:0]),.cy(-9'sd1),.dx(input_fmap_54[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O42_N14_S1),.chainout(chainout_14_O42));
logic signed [63:0] chainout_16_O42; 
logic signed [63:0] O42_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O42(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_55[7:0]),.ay( 9'sd1),.bx(input_fmap_56[7:0]),.by( 9'sd1),.cx(input_fmap_57[7:0]),.cy( 9'sd1),.dx(input_fmap_58[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O42_N16_S1),.chainout(chainout_16_O42));
logic signed [63:0] chainout_18_O42; 
logic signed [63:0] O42_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O42(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_59[7:0]),.ay(-9'sd1),.bx(input_fmap_61[7:0]),.by( 9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O42_N18_S1),.chainout(chainout_18_O42));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O42_N0_S2;		always @(posedge clk) O42_N0_S2 <=     O42_N0_S1  +  O42_N2_S1 ;
 logic signed [21:0] O42_N2_S2;		always @(posedge clk) O42_N2_S2 <=     O42_N4_S1  +  O42_N6_S1 ;
 logic signed [21:0] O42_N4_S2;		always @(posedge clk) O42_N4_S2 <=     O42_N8_S1  +  O42_N10_S1 ;
 logic signed [21:0] O42_N6_S2;		always @(posedge clk) O42_N6_S2 <=     O42_N12_S1  +  O42_N14_S1 ;
 logic signed [21:0] O42_N8_S2;		always @(posedge clk) O42_N8_S2 <=     O42_N16_S1  +  O42_N18_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O42_N0_S3;		always @(posedge clk) O42_N0_S3 <=     O42_N0_S2  +  O42_N2_S2 ;
 logic signed [22:0] O42_N2_S3;		always @(posedge clk) O42_N2_S3 <=     O42_N4_S2  +  O42_N6_S2 ;
 logic signed [22:0] O42_N4_S3;		always @(posedge clk) O42_N4_S3 <=     O42_N8_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O42_N0_S4;		always @(posedge clk) O42_N0_S4 <=     O42_N0_S3  +  O42_N2_S3 ;
 logic signed [23:0] O42_N2_S4;		always @(posedge clk) O42_N2_S4 <=     O42_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O42_N0_S5;		always @(posedge clk) O42_N0_S5 <=     O42_N0_S4  +  O42_N2_S4 ;
 assign conv_mac_42 = O42_N0_S5;

logic signed [31:0] conv_mac_43;
logic signed [63:0] chainout_0_O43; 
logic signed [63:0] O43_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O43(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd3),.bx(input_fmap_3[7:0]),.by( 9'sd1),.cx(input_fmap_6[7:0]),.cy( 9'sd4),.dx(input_fmap_8[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O43_N0_S1),.chainout(chainout_0_O43));
logic signed [63:0] chainout_2_O43; 
logic signed [63:0] O43_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O43(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_9[7:0]),.ay(-9'sd1),.bx(input_fmap_10[7:0]),.by(-9'sd2),.cx(input_fmap_11[7:0]),.cy( 9'sd1),.dx(input_fmap_12[7:0]),.dy(-9'sd3),.chainin(63'd0),.result(O43_N2_S1),.chainout(chainout_2_O43));
logic signed [63:0] chainout_4_O43; 
logic signed [63:0] O43_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O43(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_13[7:0]),.ay(-9'sd1),.bx(input_fmap_14[7:0]),.by(-9'sd2),.cx(input_fmap_16[7:0]),.cy( 9'sd1),.dx(input_fmap_17[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O43_N4_S1),.chainout(chainout_4_O43));
logic signed [63:0] chainout_6_O43; 
logic signed [63:0] O43_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O43(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_18[7:0]),.ay(-9'sd3),.bx(input_fmap_19[7:0]),.by( 9'sd2),.cx(input_fmap_20[7:0]),.cy( 9'sd1),.dx(input_fmap_21[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O43_N6_S1),.chainout(chainout_6_O43));
logic signed [63:0] chainout_8_O43; 
logic signed [63:0] O43_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O43(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_22[7:0]),.ay(-9'sd4),.bx(input_fmap_23[7:0]),.by( 9'sd3),.cx(input_fmap_24[7:0]),.cy(-9'sd3),.dx(input_fmap_25[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O43_N8_S1),.chainout(chainout_8_O43));
logic signed [63:0] chainout_10_O43; 
logic signed [63:0] O43_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O43(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_27[7:0]),.ay(-9'sd1),.bx(input_fmap_28[7:0]),.by( 9'sd4),.cx(input_fmap_29[7:0]),.cy( 9'sd1),.dx(input_fmap_30[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O43_N10_S1),.chainout(chainout_10_O43));
logic signed [63:0] chainout_12_O43; 
logic signed [63:0] O43_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O43(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_31[7:0]),.ay(-9'sd1),.bx(input_fmap_33[7:0]),.by(-9'sd3),.cx(input_fmap_34[7:0]),.cy(-9'sd3),.dx(input_fmap_35[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O43_N12_S1),.chainout(chainout_12_O43));
logic signed [63:0] chainout_14_O43; 
logic signed [63:0] O43_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O43(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_36[7:0]),.ay( 9'sd1),.bx(input_fmap_38[7:0]),.by(-9'sd1),.cx(input_fmap_39[7:0]),.cy( 9'sd1),.dx(input_fmap_40[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O43_N14_S1),.chainout(chainout_14_O43));
logic signed [63:0] chainout_16_O43; 
logic signed [63:0] O43_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O43(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_41[7:0]),.ay( 9'sd2),.bx(input_fmap_42[7:0]),.by( 9'sd4),.cx(input_fmap_43[7:0]),.cy( 9'sd2),.dx(input_fmap_44[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O43_N16_S1),.chainout(chainout_16_O43));
logic signed [63:0] chainout_18_O43; 
logic signed [63:0] O43_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O43(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_46[7:0]),.ay(-9'sd1),.bx(input_fmap_47[7:0]),.by(-9'sd2),.cx(input_fmap_48[7:0]),.cy( 9'sd1),.dx(input_fmap_49[7:0]),.dy( 9'sd3),.chainin(63'd0),.result(O43_N18_S1),.chainout(chainout_18_O43));
logic signed [63:0] chainout_20_O43; 
logic signed [63:0] O43_N20_S1; 
 int_sop_4_wrapper int_sop_4_inst_20_O43(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_50[7:0]),.ay(-9'sd4),.bx(input_fmap_51[7:0]),.by( 9'sd1),.cx(input_fmap_52[7:0]),.cy( 9'sd1),.dx(input_fmap_53[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O43_N20_S1),.chainout(chainout_20_O43));
logic signed [63:0] chainout_22_O43; 
logic signed [63:0] O43_N22_S1; 
 int_sop_4_wrapper int_sop_4_inst_22_O43(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_54[7:0]),.ay(-9'sd2),.bx(input_fmap_55[7:0]),.by( 9'sd3),.cx(input_fmap_56[7:0]),.cy( 9'sd3),.dx(input_fmap_57[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O43_N22_S1),.chainout(chainout_22_O43));
logic signed [63:0] chainout_24_O43; 
logic signed [63:0] O43_N24_S1; 
 int_sop_4_wrapper int_sop_4_inst_24_O43(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_58[7:0]),.ay(-9'sd2),.bx(input_fmap_60[7:0]),.by(-9'sd2),.cx(input_fmap_62[7:0]),.cy(-9'sd1),.dx(input_fmap_63[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O43_N24_S1),.chainout(chainout_24_O43));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O43_N0_S2;		always @(posedge clk) O43_N0_S2 <=     O43_N0_S1  +  O43_N2_S1 ;
 logic signed [21:0] O43_N2_S2;		always @(posedge clk) O43_N2_S2 <=     O43_N4_S1  +  O43_N6_S1 ;
 logic signed [21:0] O43_N4_S2;		always @(posedge clk) O43_N4_S2 <=     O43_N8_S1  +  O43_N10_S1 ;
 logic signed [21:0] O43_N6_S2;		always @(posedge clk) O43_N6_S2 <=     O43_N12_S1  +  O43_N14_S1 ;
 logic signed [21:0] O43_N8_S2;		always @(posedge clk) O43_N8_S2 <=     O43_N16_S1  +  O43_N18_S1 ;
 logic signed [21:0] O43_N10_S2;		always @(posedge clk) O43_N10_S2 <=     O43_N20_S1  +  O43_N22_S1 ;
 logic signed [21:0] O43_N12_S2;		always @(posedge clk) O43_N12_S2 <=     O43_N24_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O43_N0_S3;		always @(posedge clk) O43_N0_S3 <=     O43_N0_S2  +  O43_N2_S2 ;
 logic signed [22:0] O43_N2_S3;		always @(posedge clk) O43_N2_S3 <=     O43_N4_S2  +  O43_N6_S2 ;
 logic signed [22:0] O43_N4_S3;		always @(posedge clk) O43_N4_S3 <=     O43_N8_S2  +  O43_N10_S2 ;
 logic signed [22:0] O43_N6_S3;		always @(posedge clk) O43_N6_S3 <=     O43_N12_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O43_N0_S4;		always @(posedge clk) O43_N0_S4 <=     O43_N0_S3  +  O43_N2_S3 ;
 logic signed [23:0] O43_N2_S4;		always @(posedge clk) O43_N2_S4 <=     O43_N4_S3  +  O43_N6_S3 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O43_N0_S5;		always @(posedge clk) O43_N0_S5 <=     O43_N0_S4  +  O43_N2_S4 ;
 assign conv_mac_43 = O43_N0_S5;

logic signed [31:0] conv_mac_44;
logic signed [63:0] chainout_0_O44; 
logic signed [63:0] O44_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O44(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_2[7:0]),.ay(-9'sd1),.bx(input_fmap_5[7:0]),.by( 9'sd1),.cx(input_fmap_15[7:0]),.cy(-9'sd1),.dx(input_fmap_26[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O44_N0_S1),.chainout(chainout_0_O44));
logic signed [63:0] chainout_2_O44; 
logic signed [63:0] O44_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O44(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_29[7:0]),.ay( 9'sd1),.bx(input_fmap_31[7:0]),.by( 9'sd1),.cx(input_fmap_35[7:0]),.cy(-9'sd1),.dx(input_fmap_47[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O44_N2_S1),.chainout(chainout_2_O44));
logic signed [63:0] chainout_4_O44; 
logic signed [63:0] O44_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O44(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_49[7:0]),.ay( 9'sd1),.bx(input_fmap_51[7:0]),.by( 9'sd1),.cx(input_fmap_54[7:0]),.cy(-9'sd1),.dx(input_fmap_57[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O44_N4_S1),.chainout(chainout_4_O44));
logic signed [63:0] chainout_6_O44; 
logic signed [63:0] O44_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O44(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_59[7:0]),.ay( 9'sd1),.bx(input_fmap_61[7:0]),.by(-9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O44_N6_S1),.chainout(chainout_6_O44));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O44_N0_S2;		always @(posedge clk) O44_N0_S2 <=     O44_N0_S1  +  O44_N2_S1 ;
 logic signed [21:0] O44_N2_S2;		always @(posedge clk) O44_N2_S2 <=     O44_N4_S1  +  O44_N6_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O44_N0_S3;		always @(posedge clk) O44_N0_S3 <=     O44_N0_S2  +  O44_N2_S2 ;
 assign conv_mac_44 = O44_N0_S3;

logic signed [31:0] conv_mac_45;
logic signed [63:0] chainout_0_O45; 
logic signed [63:0] O45_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O45(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd1),.bx(input_fmap_3[7:0]),.by(-9'sd1),.cx(input_fmap_4[7:0]),.cy( 9'sd1),.dx(input_fmap_5[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O45_N0_S1),.chainout(chainout_0_O45));
logic signed [63:0] chainout_2_O45; 
logic signed [63:0] O45_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O45(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_6[7:0]),.ay(-9'sd1),.bx(input_fmap_8[7:0]),.by(-9'sd1),.cx(input_fmap_9[7:0]),.cy(-9'sd1),.dx(input_fmap_10[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O45_N2_S1),.chainout(chainout_2_O45));
logic signed [63:0] chainout_4_O45; 
logic signed [63:0] O45_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O45(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_11[7:0]),.ay( 9'sd3),.bx(input_fmap_12[7:0]),.by(-9'sd1),.cx(input_fmap_13[7:0]),.cy(-9'sd3),.dx(input_fmap_16[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O45_N4_S1),.chainout(chainout_4_O45));
logic signed [63:0] chainout_6_O45; 
logic signed [63:0] O45_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O45(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_18[7:0]),.ay(-9'sd1),.bx(input_fmap_20[7:0]),.by( 9'sd1),.cx(input_fmap_22[7:0]),.cy( 9'sd1),.dx(input_fmap_23[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O45_N6_S1),.chainout(chainout_6_O45));
logic signed [63:0] chainout_8_O45; 
logic signed [63:0] O45_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O45(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_24[7:0]),.ay(-9'sd1),.bx(input_fmap_25[7:0]),.by(-9'sd1),.cx(input_fmap_27[7:0]),.cy(-9'sd1),.dx(input_fmap_28[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O45_N8_S1),.chainout(chainout_8_O45));
logic signed [63:0] chainout_10_O45; 
logic signed [63:0] O45_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O45(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_31[7:0]),.ay(-9'sd1),.bx(input_fmap_32[7:0]),.by(-9'sd1),.cx(input_fmap_33[7:0]),.cy(-9'sd2),.dx(input_fmap_35[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O45_N10_S1),.chainout(chainout_10_O45));
logic signed [63:0] chainout_12_O45; 
logic signed [63:0] O45_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O45(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_36[7:0]),.ay( 9'sd1),.bx(input_fmap_37[7:0]),.by( 9'sd3),.cx(input_fmap_39[7:0]),.cy(-9'sd1),.dx(input_fmap_40[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O45_N12_S1),.chainout(chainout_12_O45));
logic signed [63:0] chainout_14_O45; 
logic signed [63:0] O45_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O45(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_42[7:0]),.ay( 9'sd1),.bx(input_fmap_43[7:0]),.by( 9'sd1),.cx(input_fmap_46[7:0]),.cy(-9'sd1),.dx(input_fmap_47[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O45_N14_S1),.chainout(chainout_14_O45));
logic signed [63:0] chainout_16_O45; 
logic signed [63:0] O45_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O45(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_48[7:0]),.ay(-9'sd2),.bx(input_fmap_49[7:0]),.by(-9'sd1),.cx(input_fmap_50[7:0]),.cy(-9'sd1),.dx(input_fmap_51[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O45_N16_S1),.chainout(chainout_16_O45));
logic signed [63:0] chainout_18_O45; 
logic signed [63:0] O45_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O45(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_52[7:0]),.ay( 9'sd1),.bx(input_fmap_54[7:0]),.by(-9'sd1),.cx(input_fmap_55[7:0]),.cy( 9'sd1),.dx(input_fmap_56[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O45_N18_S1),.chainout(chainout_18_O45));
logic signed [63:0] chainout_20_O45; 
logic signed [63:0] O45_N20_S1; 
 int_sop_4_wrapper int_sop_4_inst_20_O45(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_57[7:0]),.ay( 9'sd1),.bx(input_fmap_58[7:0]),.by(-9'sd1),.cx(input_fmap_59[7:0]),.cy( 9'sd1),.dx(input_fmap_63[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O45_N20_S1),.chainout(chainout_20_O45));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O45_N0_S2;		always @(posedge clk) O45_N0_S2 <=     O45_N0_S1  +  O45_N2_S1 ;
 logic signed [21:0] O45_N2_S2;		always @(posedge clk) O45_N2_S2 <=     O45_N4_S1  +  O45_N6_S1 ;
 logic signed [21:0] O45_N4_S2;		always @(posedge clk) O45_N4_S2 <=     O45_N8_S1  +  O45_N10_S1 ;
 logic signed [21:0] O45_N6_S2;		always @(posedge clk) O45_N6_S2 <=     O45_N12_S1  +  O45_N14_S1 ;
 logic signed [21:0] O45_N8_S2;		always @(posedge clk) O45_N8_S2 <=     O45_N16_S1  +  O45_N18_S1 ;
 logic signed [21:0] O45_N10_S2;		always @(posedge clk) O45_N10_S2 <=     O45_N20_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O45_N0_S3;		always @(posedge clk) O45_N0_S3 <=     O45_N0_S2  +  O45_N2_S2 ;
 logic signed [22:0] O45_N2_S3;		always @(posedge clk) O45_N2_S3 <=     O45_N4_S2  +  O45_N6_S2 ;
 logic signed [22:0] O45_N4_S3;		always @(posedge clk) O45_N4_S3 <=     O45_N8_S2  +  O45_N10_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O45_N0_S4;		always @(posedge clk) O45_N0_S4 <=     O45_N0_S3  +  O45_N2_S3 ;
 logic signed [23:0] O45_N2_S4;		always @(posedge clk) O45_N2_S4 <=     O45_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O45_N0_S5;		always @(posedge clk) O45_N0_S5 <=     O45_N0_S4  +  O45_N2_S4 ;
 assign conv_mac_45 = O45_N0_S5;

logic signed [31:0] conv_mac_46;
logic signed [63:0] chainout_0_O46; 
logic signed [63:0] O46_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O46(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd1),.bx(input_fmap_1[7:0]),.by( 9'sd1),.cx(input_fmap_7[7:0]),.cy(-9'sd1),.dx(input_fmap_9[7:0]),.dy( 9'sd4),.chainin(63'd0),.result(O46_N0_S1),.chainout(chainout_0_O46));
logic signed [63:0] chainout_2_O46; 
logic signed [63:0] O46_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O46(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_14[7:0]),.ay( 9'sd1),.bx(input_fmap_16[7:0]),.by(-9'sd1),.cx(input_fmap_18[7:0]),.cy(-9'sd1),.dx(input_fmap_20[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O46_N2_S1),.chainout(chainout_2_O46));
logic signed [63:0] chainout_4_O46; 
logic signed [63:0] O46_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O46(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_22[7:0]),.ay( 9'sd1),.bx(input_fmap_23[7:0]),.by(-9'sd1),.cx(input_fmap_27[7:0]),.cy( 9'sd1),.dx(input_fmap_30[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O46_N4_S1),.chainout(chainout_4_O46));
logic signed [63:0] chainout_6_O46; 
logic signed [63:0] O46_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O46(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_32[7:0]),.ay(-9'sd1),.bx(input_fmap_33[7:0]),.by(-9'sd1),.cx(input_fmap_35[7:0]),.cy(-9'sd1),.dx(input_fmap_36[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O46_N6_S1),.chainout(chainout_6_O46));
logic signed [63:0] chainout_8_O46; 
logic signed [63:0] O46_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O46(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_38[7:0]),.ay(-9'sd1),.bx(input_fmap_39[7:0]),.by( 9'sd1),.cx(input_fmap_43[7:0]),.cy( 9'sd1),.dx(input_fmap_45[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O46_N8_S1),.chainout(chainout_8_O46));
logic signed [63:0] chainout_10_O46; 
logic signed [63:0] O46_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O46(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_46[7:0]),.ay(-9'sd2),.bx(input_fmap_53[7:0]),.by( 9'sd1),.cx(input_fmap_58[7:0]),.cy( 9'sd1),.dx(input_fmap_60[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O46_N10_S1),.chainout(chainout_10_O46));
logic signed [63:0] chainout_12_O46; 
logic signed [63:0] O46_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O46(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_63[7:0]),.ay( 9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O46_N12_S1),.chainout(chainout_12_O46));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O46_N0_S2;		always @(posedge clk) O46_N0_S2 <=     O46_N0_S1  +  O46_N2_S1 ;
 logic signed [21:0] O46_N2_S2;		always @(posedge clk) O46_N2_S2 <=     O46_N4_S1  +  O46_N6_S1 ;
 logic signed [21:0] O46_N4_S2;		always @(posedge clk) O46_N4_S2 <=     O46_N8_S1  +  O46_N10_S1 ;
 logic signed [21:0] O46_N6_S2;		always @(posedge clk) O46_N6_S2 <=     O46_N12_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O46_N0_S3;		always @(posedge clk) O46_N0_S3 <=     O46_N0_S2  +  O46_N2_S2 ;
 logic signed [22:0] O46_N2_S3;		always @(posedge clk) O46_N2_S3 <=     O46_N4_S2  +  O46_N6_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O46_N0_S4;		always @(posedge clk) O46_N0_S4 <=     O46_N0_S3  +  O46_N2_S3 ;
 assign conv_mac_46 = O46_N0_S4;

logic signed [31:0] conv_mac_47;
logic signed [63:0] chainout_0_O47; 
logic signed [63:0] O47_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O47(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd1),.bx(input_fmap_2[7:0]),.by(-9'sd1),.cx(input_fmap_18[7:0]),.cy(-9'sd1),.dx(input_fmap_19[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O47_N0_S1),.chainout(chainout_0_O47));
logic signed [63:0] chainout_2_O47; 
logic signed [63:0] O47_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O47(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_25[7:0]),.ay(-9'sd1),.bx(input_fmap_40[7:0]),.by( 9'sd1),.cx(input_fmap_43[7:0]),.cy(-9'sd1),.dx(input_fmap_46[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O47_N2_S1),.chainout(chainout_2_O47));
logic signed [63:0] chainout_4_O47; 
logic signed [63:0] O47_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O47(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_57[7:0]),.ay(-9'sd1),.bx(input_fmap_60[7:0]),.by( 9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O47_N4_S1),.chainout(chainout_4_O47));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O47_N0_S2;		always @(posedge clk) O47_N0_S2 <=     O47_N0_S1  +  O47_N2_S1 ;
 logic signed [21:0] O47_N2_S2;		always @(posedge clk) O47_N2_S2 <=     O47_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O47_N0_S3;		always @(posedge clk) O47_N0_S3 <=     O47_N0_S2  +  O47_N2_S2 ;
 assign conv_mac_47 = O47_N0_S3;

logic signed [31:0] conv_mac_48;
logic signed [63:0] chainout_0_O48; 
logic signed [63:0] O48_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O48(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd1),.bx(input_fmap_1[7:0]),.by( 9'sd2),.cx(input_fmap_3[7:0]),.cy(-9'sd1),.dx(input_fmap_5[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O48_N0_S1),.chainout(chainout_0_O48));
logic signed [63:0] chainout_2_O48; 
logic signed [63:0] O48_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O48(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_6[7:0]),.ay(-9'sd1),.bx(input_fmap_7[7:0]),.by(-9'sd1),.cx(input_fmap_8[7:0]),.cy( 9'sd1),.dx(input_fmap_10[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O48_N2_S1),.chainout(chainout_2_O48));
logic signed [63:0] chainout_4_O48; 
logic signed [63:0] O48_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O48(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_12[7:0]),.ay(-9'sd1),.bx(input_fmap_13[7:0]),.by( 9'sd1),.cx(input_fmap_14[7:0]),.cy(-9'sd1),.dx(input_fmap_17[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O48_N4_S1),.chainout(chainout_4_O48));
logic signed [63:0] chainout_6_O48; 
logic signed [63:0] O48_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O48(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_18[7:0]),.ay(-9'sd1),.bx(input_fmap_19[7:0]),.by(-9'sd1),.cx(input_fmap_21[7:0]),.cy(-9'sd1),.dx(input_fmap_22[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O48_N6_S1),.chainout(chainout_6_O48));
logic signed [63:0] chainout_8_O48; 
logic signed [63:0] O48_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O48(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_25[7:0]),.ay(-9'sd4),.bx(input_fmap_26[7:0]),.by( 9'sd2),.cx(input_fmap_27[7:0]),.cy( 9'sd1),.dx(input_fmap_29[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O48_N8_S1),.chainout(chainout_8_O48));
logic signed [63:0] chainout_10_O48; 
logic signed [63:0] O48_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O48(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_31[7:0]),.ay( 9'sd1),.bx(input_fmap_32[7:0]),.by(-9'sd1),.cx(input_fmap_34[7:0]),.cy(-9'sd1),.dx(input_fmap_35[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O48_N10_S1),.chainout(chainout_10_O48));
logic signed [63:0] chainout_12_O48; 
logic signed [63:0] O48_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O48(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_36[7:0]),.ay(-9'sd1),.bx(input_fmap_39[7:0]),.by(-9'sd1),.cx(input_fmap_40[7:0]),.cy( 9'sd1),.dx(input_fmap_42[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O48_N12_S1),.chainout(chainout_12_O48));
logic signed [63:0] chainout_14_O48; 
logic signed [63:0] O48_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O48(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_44[7:0]),.ay( 9'sd1),.bx(input_fmap_45[7:0]),.by(-9'sd2),.cx(input_fmap_49[7:0]),.cy(-9'sd2),.dx(input_fmap_50[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O48_N14_S1),.chainout(chainout_14_O48));
logic signed [63:0] chainout_16_O48; 
logic signed [63:0] O48_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O48(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_51[7:0]),.ay(-9'sd1),.bx(input_fmap_52[7:0]),.by(-9'sd2),.cx(input_fmap_57[7:0]),.cy( 9'sd1),.dx(input_fmap_59[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O48_N16_S1),.chainout(chainout_16_O48));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O48_N0_S2;		always @(posedge clk) O48_N0_S2 <=     O48_N0_S1  +  O48_N2_S1 ;
 logic signed [21:0] O48_N2_S2;		always @(posedge clk) O48_N2_S2 <=     O48_N4_S1  +  O48_N6_S1 ;
 logic signed [21:0] O48_N4_S2;		always @(posedge clk) O48_N4_S2 <=     O48_N8_S1  +  O48_N10_S1 ;
 logic signed [21:0] O48_N6_S2;		always @(posedge clk) O48_N6_S2 <=     O48_N12_S1  +  O48_N14_S1 ;
 logic signed [21:0] O48_N8_S2;		always @(posedge clk) O48_N8_S2 <=     O48_N16_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O48_N0_S3;		always @(posedge clk) O48_N0_S3 <=     O48_N0_S2  +  O48_N2_S2 ;
 logic signed [22:0] O48_N2_S3;		always @(posedge clk) O48_N2_S3 <=     O48_N4_S2  +  O48_N6_S2 ;
 logic signed [22:0] O48_N4_S3;		always @(posedge clk) O48_N4_S3 <=     O48_N8_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O48_N0_S4;		always @(posedge clk) O48_N0_S4 <=     O48_N0_S3  +  O48_N2_S3 ;
 logic signed [23:0] O48_N2_S4;		always @(posedge clk) O48_N2_S4 <=     O48_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O48_N0_S5;		always @(posedge clk) O48_N0_S5 <=     O48_N0_S4  +  O48_N2_S4 ;
 assign conv_mac_48 = O48_N0_S5;

logic signed [31:0] conv_mac_49;
logic signed [63:0] chainout_0_O49; 
logic signed [63:0] O49_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O49(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd1),.bx(input_fmap_1[7:0]),.by(-9'sd1),.cx(input_fmap_2[7:0]),.cy(-9'sd1),.dx(input_fmap_3[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O49_N0_S1),.chainout(chainout_0_O49));
logic signed [63:0] chainout_2_O49; 
logic signed [63:0] O49_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O49(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_4[7:0]),.ay( 9'sd3),.bx(input_fmap_5[7:0]),.by(-9'sd2),.cx(input_fmap_6[7:0]),.cy( 9'sd1),.dx(input_fmap_8[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O49_N2_S1),.chainout(chainout_2_O49));
logic signed [63:0] chainout_4_O49; 
logic signed [63:0] O49_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O49(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_9[7:0]),.ay( 9'sd1),.bx(input_fmap_10[7:0]),.by(-9'sd1),.cx(input_fmap_11[7:0]),.cy( 9'sd2),.dx(input_fmap_12[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O49_N4_S1),.chainout(chainout_4_O49));
logic signed [63:0] chainout_6_O49; 
logic signed [63:0] O49_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O49(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_14[7:0]),.ay( 9'sd1),.bx(input_fmap_17[7:0]),.by( 9'sd4),.cx(input_fmap_19[7:0]),.cy( 9'sd1),.dx(input_fmap_21[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O49_N6_S1),.chainout(chainout_6_O49));
logic signed [63:0] chainout_8_O49; 
logic signed [63:0] O49_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O49(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_22[7:0]),.ay(-9'sd2),.bx(input_fmap_27[7:0]),.by( 9'sd1),.cx(input_fmap_29[7:0]),.cy(-9'sd2),.dx(input_fmap_30[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O49_N8_S1),.chainout(chainout_8_O49));
logic signed [63:0] chainout_10_O49; 
logic signed [63:0] O49_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O49(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_33[7:0]),.ay(-9'sd1),.bx(input_fmap_34[7:0]),.by(-9'sd2),.cx(input_fmap_37[7:0]),.cy(-9'sd2),.dx(input_fmap_39[7:0]),.dy( 9'sd3),.chainin(63'd0),.result(O49_N10_S1),.chainout(chainout_10_O49));
logic signed [63:0] chainout_12_O49; 
logic signed [63:0] O49_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O49(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_40[7:0]),.ay(-9'sd1),.bx(input_fmap_42[7:0]),.by( 9'sd2),.cx(input_fmap_43[7:0]),.cy( 9'sd1),.dx(input_fmap_44[7:0]),.dy( 9'sd3),.chainin(63'd0),.result(O49_N12_S1),.chainout(chainout_12_O49));
logic signed [63:0] chainout_14_O49; 
logic signed [63:0] O49_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O49(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_46[7:0]),.ay(-9'sd1),.bx(input_fmap_48[7:0]),.by( 9'sd1),.cx(input_fmap_50[7:0]),.cy( 9'sd4),.dx(input_fmap_51[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O49_N14_S1),.chainout(chainout_14_O49));
logic signed [63:0] chainout_16_O49; 
logic signed [63:0] O49_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O49(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_52[7:0]),.ay(-9'sd2),.bx(input_fmap_54[7:0]),.by(-9'sd1),.cx(input_fmap_55[7:0]),.cy(-9'sd1),.dx(input_fmap_61[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O49_N16_S1),.chainout(chainout_16_O49));
logic signed [63:0] chainout_18_O49; 
logic signed [63:0] O49_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O49(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_62[7:0]),.ay(-9'sd2),.bx(input_fmap_63[7:0]),.by(-9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O49_N18_S1),.chainout(chainout_18_O49));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O49_N0_S2;		always @(posedge clk) O49_N0_S2 <=     O49_N0_S1  +  O49_N2_S1 ;
 logic signed [21:0] O49_N2_S2;		always @(posedge clk) O49_N2_S2 <=     O49_N4_S1  +  O49_N6_S1 ;
 logic signed [21:0] O49_N4_S2;		always @(posedge clk) O49_N4_S2 <=     O49_N8_S1  +  O49_N10_S1 ;
 logic signed [21:0] O49_N6_S2;		always @(posedge clk) O49_N6_S2 <=     O49_N12_S1  +  O49_N14_S1 ;
 logic signed [21:0] O49_N8_S2;		always @(posedge clk) O49_N8_S2 <=     O49_N16_S1  +  O49_N18_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O49_N0_S3;		always @(posedge clk) O49_N0_S3 <=     O49_N0_S2  +  O49_N2_S2 ;
 logic signed [22:0] O49_N2_S3;		always @(posedge clk) O49_N2_S3 <=     O49_N4_S2  +  O49_N6_S2 ;
 logic signed [22:0] O49_N4_S3;		always @(posedge clk) O49_N4_S3 <=     O49_N8_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O49_N0_S4;		always @(posedge clk) O49_N0_S4 <=     O49_N0_S3  +  O49_N2_S3 ;
 logic signed [23:0] O49_N2_S4;		always @(posedge clk) O49_N2_S4 <=     O49_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O49_N0_S5;		always @(posedge clk) O49_N0_S5 <=     O49_N0_S4  +  O49_N2_S4 ;
 assign conv_mac_49 = O49_N0_S5;

logic signed [31:0] conv_mac_50;
logic signed [63:0] chainout_0_O50; 
logic signed [63:0] O50_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O50(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay(-9'sd1),.bx(input_fmap_2[7:0]),.by( 9'sd1),.cx(input_fmap_10[7:0]),.cy(-9'sd1),.dx(input_fmap_12[7:0]),.dy( 9'sd5),.chainin(63'd0),.result(O50_N0_S1),.chainout(chainout_0_O50));
logic signed [63:0] chainout_2_O50; 
logic signed [63:0] O50_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O50(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_15[7:0]),.ay( 9'sd1),.bx(input_fmap_16[7:0]),.by(-9'sd1),.cx(input_fmap_17[7:0]),.cy( 9'sd1),.dx(input_fmap_18[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O50_N2_S1),.chainout(chainout_2_O50));
logic signed [63:0] chainout_4_O50; 
logic signed [63:0] O50_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O50(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_21[7:0]),.ay( 9'sd1),.bx(input_fmap_24[7:0]),.by(-9'sd1),.cx(input_fmap_28[7:0]),.cy(-9'sd2),.dx(input_fmap_29[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O50_N4_S1),.chainout(chainout_4_O50));
logic signed [63:0] chainout_6_O50; 
logic signed [63:0] O50_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O50(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_31[7:0]),.ay(-9'sd1),.bx(input_fmap_33[7:0]),.by( 9'sd1),.cx(input_fmap_36[7:0]),.cy(-9'sd1),.dx(input_fmap_41[7:0]),.dy( 9'sd3),.chainin(63'd0),.result(O50_N6_S1),.chainout(chainout_6_O50));
logic signed [63:0] chainout_8_O50; 
logic signed [63:0] O50_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O50(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_47[7:0]),.ay(-9'sd1),.bx(input_fmap_53[7:0]),.by( 9'sd1),.cx(input_fmap_55[7:0]),.cy( 9'sd1),.dx(input_fmap_56[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O50_N8_S1),.chainout(chainout_8_O50));
logic signed [63:0] chainout_10_O50; 
logic signed [63:0] O50_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O50(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_57[7:0]),.ay(-9'sd1),.bx(input_fmap_59[7:0]),.by(-9'sd1),.cx(input_fmap_63[7:0]),.cy(-9'sd1),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O50_N10_S1),.chainout(chainout_10_O50));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O50_N0_S2;		always @(posedge clk) O50_N0_S2 <=     O50_N0_S1  +  O50_N2_S1 ;
 logic signed [21:0] O50_N2_S2;		always @(posedge clk) O50_N2_S2 <=     O50_N4_S1  +  O50_N6_S1 ;
 logic signed [21:0] O50_N4_S2;		always @(posedge clk) O50_N4_S2 <=     O50_N8_S1  +  O50_N10_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O50_N0_S3;		always @(posedge clk) O50_N0_S3 <=     O50_N0_S2  +  O50_N2_S2 ;
 logic signed [22:0] O50_N2_S3;		always @(posedge clk) O50_N2_S3 <=     O50_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O50_N0_S4;		always @(posedge clk) O50_N0_S4 <=     O50_N0_S3  +  O50_N2_S3 ;
 assign conv_mac_50 = O50_N0_S4;

logic signed [31:0] conv_mac_51;
logic signed [63:0] chainout_0_O51; 
logic signed [63:0] O51_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O51(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd1),.bx(input_fmap_4[7:0]),.by( 9'sd1),.cx(input_fmap_6[7:0]),.cy( 9'sd2),.dx(input_fmap_7[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O51_N0_S1),.chainout(chainout_0_O51));
logic signed [63:0] chainout_2_O51; 
logic signed [63:0] O51_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O51(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_8[7:0]),.ay(-9'sd1),.bx(input_fmap_12[7:0]),.by( 9'sd2),.cx(input_fmap_14[7:0]),.cy( 9'sd1),.dx(input_fmap_15[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O51_N2_S1),.chainout(chainout_2_O51));
logic signed [63:0] chainout_4_O51; 
logic signed [63:0] O51_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O51(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_16[7:0]),.ay(-9'sd1),.bx(input_fmap_18[7:0]),.by( 9'sd1),.cx(input_fmap_19[7:0]),.cy(-9'sd1),.dx(input_fmap_21[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O51_N4_S1),.chainout(chainout_4_O51));
logic signed [63:0] chainout_6_O51; 
logic signed [63:0] O51_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O51(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_29[7:0]),.ay( 9'sd1),.bx(input_fmap_34[7:0]),.by(-9'sd1),.cx(input_fmap_35[7:0]),.cy( 9'sd1),.dx(input_fmap_39[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O51_N6_S1),.chainout(chainout_6_O51));
logic signed [63:0] chainout_8_O51; 
logic signed [63:0] O51_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O51(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_40[7:0]),.ay( 9'sd1),.bx(input_fmap_47[7:0]),.by( 9'sd1),.cx(input_fmap_48[7:0]),.cy( 9'sd1),.dx(input_fmap_49[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O51_N8_S1),.chainout(chainout_8_O51));
logic signed [63:0] chainout_10_O51; 
logic signed [63:0] O51_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O51(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_53[7:0]),.ay(-9'sd1),.bx(input_fmap_57[7:0]),.by(-9'sd1),.cx(input_fmap_59[7:0]),.cy(-9'sd1),.dx(input_fmap_60[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O51_N10_S1),.chainout(chainout_10_O51));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O51_N0_S2;		always @(posedge clk) O51_N0_S2 <=     O51_N0_S1  +  O51_N2_S1 ;
 logic signed [21:0] O51_N2_S2;		always @(posedge clk) O51_N2_S2 <=     O51_N4_S1  +  O51_N6_S1 ;
 logic signed [21:0] O51_N4_S2;		always @(posedge clk) O51_N4_S2 <=     O51_N8_S1  +  O51_N10_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O51_N0_S3;		always @(posedge clk) O51_N0_S3 <=     O51_N0_S2  +  O51_N2_S2 ;
 logic signed [22:0] O51_N2_S3;		always @(posedge clk) O51_N2_S3 <=     O51_N4_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O51_N0_S4;		always @(posedge clk) O51_N0_S4 <=     O51_N0_S3  +  O51_N2_S3 ;
 assign conv_mac_51 = O51_N0_S4;

logic signed [31:0] conv_mac_52;
logic signed [63:0] chainout_0_O52; 
logic signed [63:0] O52_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O52(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_2[7:0]),.ay(-9'sd1),.bx(input_fmap_3[7:0]),.by(-9'sd1),.cx(input_fmap_6[7:0]),.cy(-9'sd1),.dx(input_fmap_7[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O52_N0_S1),.chainout(chainout_0_O52));
logic signed [63:0] chainout_2_O52; 
logic signed [63:0] O52_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O52(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_8[7:0]),.ay(-9'sd1),.bx(input_fmap_10[7:0]),.by( 9'sd1),.cx(input_fmap_12[7:0]),.cy( 9'sd3),.dx(input_fmap_15[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O52_N2_S1),.chainout(chainout_2_O52));
logic signed [63:0] chainout_4_O52; 
logic signed [63:0] O52_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O52(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_17[7:0]),.ay( 9'sd1),.bx(input_fmap_19[7:0]),.by( 9'sd2),.cx(input_fmap_20[7:0]),.cy( 9'sd1),.dx(input_fmap_21[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O52_N4_S1),.chainout(chainout_4_O52));
logic signed [63:0] chainout_6_O52; 
logic signed [63:0] O52_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O52(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_22[7:0]),.ay(-9'sd1),.bx(input_fmap_26[7:0]),.by( 9'sd1),.cx(input_fmap_31[7:0]),.cy( 9'sd1),.dx(input_fmap_34[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O52_N6_S1),.chainout(chainout_6_O52));
logic signed [63:0] chainout_8_O52; 
logic signed [63:0] O52_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O52(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_35[7:0]),.ay(-9'sd1),.bx(input_fmap_36[7:0]),.by(-9'sd1),.cx(input_fmap_37[7:0]),.cy( 9'sd2),.dx(input_fmap_38[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O52_N8_S1),.chainout(chainout_8_O52));
logic signed [63:0] chainout_10_O52; 
logic signed [63:0] O52_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O52(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_41[7:0]),.ay( 9'sd2),.bx(input_fmap_42[7:0]),.by(-9'sd1),.cx(input_fmap_44[7:0]),.cy( 9'sd1),.dx(input_fmap_47[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O52_N10_S1),.chainout(chainout_10_O52));
logic signed [63:0] chainout_12_O52; 
logic signed [63:0] O52_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O52(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_50[7:0]),.ay(-9'sd1),.bx(input_fmap_53[7:0]),.by( 9'sd1),.cx(input_fmap_54[7:0]),.cy(-9'sd1),.dx(input_fmap_58[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O52_N12_S1),.chainout(chainout_12_O52));
logic signed [63:0] chainout_14_O52; 
logic signed [63:0] O52_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O52(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_60[7:0]),.ay( 9'sd1),.bx(input_fmap_61[7:0]),.by(-9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O52_N14_S1),.chainout(chainout_14_O52));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O52_N0_S2;		always @(posedge clk) O52_N0_S2 <=     O52_N0_S1  +  O52_N2_S1 ;
 logic signed [21:0] O52_N2_S2;		always @(posedge clk) O52_N2_S2 <=     O52_N4_S1  +  O52_N6_S1 ;
 logic signed [21:0] O52_N4_S2;		always @(posedge clk) O52_N4_S2 <=     O52_N8_S1  +  O52_N10_S1 ;
 logic signed [21:0] O52_N6_S2;		always @(posedge clk) O52_N6_S2 <=     O52_N12_S1  +  O52_N14_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O52_N0_S3;		always @(posedge clk) O52_N0_S3 <=     O52_N0_S2  +  O52_N2_S2 ;
 logic signed [22:0] O52_N2_S3;		always @(posedge clk) O52_N2_S3 <=     O52_N4_S2  +  O52_N6_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O52_N0_S4;		always @(posedge clk) O52_N0_S4 <=     O52_N0_S3  +  O52_N2_S3 ;
 assign conv_mac_52 = O52_N0_S4;

logic signed [31:0] conv_mac_53;
logic signed [63:0] chainout_0_O53; 
logic signed [63:0] O53_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O53(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd2),.bx(input_fmap_2[7:0]),.by(-9'sd1),.cx(input_fmap_3[7:0]),.cy(-9'sd1),.dx(input_fmap_4[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O53_N0_S1),.chainout(chainout_0_O53));
logic signed [63:0] chainout_2_O53; 
logic signed [63:0] O53_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O53(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_7[7:0]),.ay( 9'sd1),.bx(input_fmap_10[7:0]),.by( 9'sd2),.cx(input_fmap_12[7:0]),.cy(-9'sd1),.dx(input_fmap_14[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O53_N2_S1),.chainout(chainout_2_O53));
logic signed [63:0] chainout_4_O53; 
logic signed [63:0] O53_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O53(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_16[7:0]),.ay( 9'sd3),.bx(input_fmap_18[7:0]),.by( 9'sd1),.cx(input_fmap_19[7:0]),.cy(-9'sd2),.dx(input_fmap_20[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O53_N4_S1),.chainout(chainout_4_O53));
logic signed [63:0] chainout_6_O53; 
logic signed [63:0] O53_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O53(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_21[7:0]),.ay(-9'sd2),.bx(input_fmap_22[7:0]),.by(-9'sd1),.cx(input_fmap_23[7:0]),.cy( 9'sd2),.dx(input_fmap_27[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O53_N6_S1),.chainout(chainout_6_O53));
logic signed [63:0] chainout_8_O53; 
logic signed [63:0] O53_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O53(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_28[7:0]),.ay(-9'sd1),.bx(input_fmap_29[7:0]),.by( 9'sd1),.cx(input_fmap_31[7:0]),.cy(-9'sd1),.dx(input_fmap_33[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O53_N8_S1),.chainout(chainout_8_O53));
logic signed [63:0] chainout_10_O53; 
logic signed [63:0] O53_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O53(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_34[7:0]),.ay(-9'sd1),.bx(input_fmap_35[7:0]),.by(-9'sd3),.cx(input_fmap_36[7:0]),.cy( 9'sd1),.dx(input_fmap_38[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O53_N10_S1),.chainout(chainout_10_O53));
logic signed [63:0] chainout_12_O53; 
logic signed [63:0] O53_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O53(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_39[7:0]),.ay( 9'sd1),.bx(input_fmap_40[7:0]),.by(-9'sd1),.cx(input_fmap_41[7:0]),.cy(-9'sd2),.dx(input_fmap_42[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O53_N12_S1),.chainout(chainout_12_O53));
logic signed [63:0] chainout_14_O53; 
logic signed [63:0] O53_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O53(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_45[7:0]),.ay( 9'sd1),.bx(input_fmap_46[7:0]),.by( 9'sd1),.cx(input_fmap_47[7:0]),.cy(-9'sd1),.dx(input_fmap_51[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O53_N14_S1),.chainout(chainout_14_O53));
logic signed [63:0] chainout_16_O53; 
logic signed [63:0] O53_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O53(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_54[7:0]),.ay(-9'sd1),.bx(input_fmap_55[7:0]),.by(-9'sd1),.cx(input_fmap_56[7:0]),.cy( 9'sd1),.dx(input_fmap_57[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O53_N16_S1),.chainout(chainout_16_O53));
logic signed [63:0] chainout_18_O53; 
logic signed [63:0] O53_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O53(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_59[7:0]),.ay( 9'sd1),.bx(input_fmap_60[7:0]),.by( 9'sd2),.cx(input_fmap_61[7:0]),.cy( 9'sd1),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O53_N18_S1),.chainout(chainout_18_O53));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O53_N0_S2;		always @(posedge clk) O53_N0_S2 <=     O53_N0_S1  +  O53_N2_S1 ;
 logic signed [21:0] O53_N2_S2;		always @(posedge clk) O53_N2_S2 <=     O53_N4_S1  +  O53_N6_S1 ;
 logic signed [21:0] O53_N4_S2;		always @(posedge clk) O53_N4_S2 <=     O53_N8_S1  +  O53_N10_S1 ;
 logic signed [21:0] O53_N6_S2;		always @(posedge clk) O53_N6_S2 <=     O53_N12_S1  +  O53_N14_S1 ;
 logic signed [21:0] O53_N8_S2;		always @(posedge clk) O53_N8_S2 <=     O53_N16_S1  +  O53_N18_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O53_N0_S3;		always @(posedge clk) O53_N0_S3 <=     O53_N0_S2  +  O53_N2_S2 ;
 logic signed [22:0] O53_N2_S3;		always @(posedge clk) O53_N2_S3 <=     O53_N4_S2  +  O53_N6_S2 ;
 logic signed [22:0] O53_N4_S3;		always @(posedge clk) O53_N4_S3 <=     O53_N8_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O53_N0_S4;		always @(posedge clk) O53_N0_S4 <=     O53_N0_S3  +  O53_N2_S3 ;
 logic signed [23:0] O53_N2_S4;		always @(posedge clk) O53_N2_S4 <=     O53_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O53_N0_S5;		always @(posedge clk) O53_N0_S5 <=     O53_N0_S4  +  O53_N2_S4 ;
 assign conv_mac_53 = O53_N0_S5;

logic signed [31:0] conv_mac_54;
logic signed [63:0] chainout_0_O54; 
logic signed [63:0] O54_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O54(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd2),.bx(input_fmap_5[7:0]),.by( 9'sd1),.cx(input_fmap_7[7:0]),.cy(-9'sd1),.dx(input_fmap_8[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O54_N0_S1),.chainout(chainout_0_O54));
logic signed [63:0] chainout_2_O54; 
logic signed [63:0] O54_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O54(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_10[7:0]),.ay( 9'sd1),.bx(input_fmap_11[7:0]),.by( 9'sd1),.cx(input_fmap_12[7:0]),.cy(-9'sd1),.dx(input_fmap_13[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O54_N2_S1),.chainout(chainout_2_O54));
logic signed [63:0] chainout_4_O54; 
logic signed [63:0] O54_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O54(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_15[7:0]),.ay( 9'sd2),.bx(input_fmap_16[7:0]),.by(-9'sd1),.cx(input_fmap_19[7:0]),.cy( 9'sd1),.dx(input_fmap_20[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O54_N4_S1),.chainout(chainout_4_O54));
logic signed [63:0] chainout_6_O54; 
logic signed [63:0] O54_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O54(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_21[7:0]),.ay(-9'sd1),.bx(input_fmap_22[7:0]),.by(-9'sd1),.cx(input_fmap_24[7:0]),.cy( 9'sd1),.dx(input_fmap_25[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O54_N6_S1),.chainout(chainout_6_O54));
logic signed [63:0] chainout_8_O54; 
logic signed [63:0] O54_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O54(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_27[7:0]),.ay(-9'sd1),.bx(input_fmap_28[7:0]),.by( 9'sd1),.cx(input_fmap_29[7:0]),.cy( 9'sd2),.dx(input_fmap_30[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O54_N8_S1),.chainout(chainout_8_O54));
logic signed [63:0] chainout_10_O54; 
logic signed [63:0] O54_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O54(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_35[7:0]),.ay( 9'sd1),.bx(input_fmap_36[7:0]),.by( 9'sd1),.cx(input_fmap_38[7:0]),.cy(-9'sd1),.dx(input_fmap_39[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O54_N10_S1),.chainout(chainout_10_O54));
logic signed [63:0] chainout_12_O54; 
logic signed [63:0] O54_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O54(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_41[7:0]),.ay(-9'sd2),.bx(input_fmap_42[7:0]),.by( 9'sd1),.cx(input_fmap_43[7:0]),.cy(-9'sd1),.dx(input_fmap_45[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O54_N12_S1),.chainout(chainout_12_O54));
logic signed [63:0] chainout_14_O54; 
logic signed [63:0] O54_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O54(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_46[7:0]),.ay( 9'sd1),.bx(input_fmap_47[7:0]),.by( 9'sd1),.cx(input_fmap_50[7:0]),.cy(-9'sd1),.dx(input_fmap_51[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O54_N14_S1),.chainout(chainout_14_O54));
logic signed [63:0] chainout_16_O54; 
logic signed [63:0] O54_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O54(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_53[7:0]),.ay( 9'sd1),.bx(input_fmap_57[7:0]),.by(-9'sd1),.cx(input_fmap_59[7:0]),.cy(-9'sd1),.dx(input_fmap_61[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O54_N16_S1),.chainout(chainout_16_O54));
logic signed [63:0] chainout_18_O54; 
logic signed [63:0] O54_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O54(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_63[7:0]),.ay( 9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O54_N18_S1),.chainout(chainout_18_O54));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O54_N0_S2;		always @(posedge clk) O54_N0_S2 <=     O54_N0_S1  +  O54_N2_S1 ;
 logic signed [21:0] O54_N2_S2;		always @(posedge clk) O54_N2_S2 <=     O54_N4_S1  +  O54_N6_S1 ;
 logic signed [21:0] O54_N4_S2;		always @(posedge clk) O54_N4_S2 <=     O54_N8_S1  +  O54_N10_S1 ;
 logic signed [21:0] O54_N6_S2;		always @(posedge clk) O54_N6_S2 <=     O54_N12_S1  +  O54_N14_S1 ;
 logic signed [21:0] O54_N8_S2;		always @(posedge clk) O54_N8_S2 <=     O54_N16_S1  +  O54_N18_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O54_N0_S3;		always @(posedge clk) O54_N0_S3 <=     O54_N0_S2  +  O54_N2_S2 ;
 logic signed [22:0] O54_N2_S3;		always @(posedge clk) O54_N2_S3 <=     O54_N4_S2  +  O54_N6_S2 ;
 logic signed [22:0] O54_N4_S3;		always @(posedge clk) O54_N4_S3 <=     O54_N8_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O54_N0_S4;		always @(posedge clk) O54_N0_S4 <=     O54_N0_S3  +  O54_N2_S3 ;
 logic signed [23:0] O54_N2_S4;		always @(posedge clk) O54_N2_S4 <=     O54_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O54_N0_S5;		always @(posedge clk) O54_N0_S5 <=     O54_N0_S4  +  O54_N2_S4 ;
 assign conv_mac_54 = O54_N0_S5;

logic signed [31:0] conv_mac_55;
logic signed [63:0] chainout_0_O55; 
logic signed [63:0] O55_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O55(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd1),.bx(input_fmap_1[7:0]),.by( 9'sd1),.cx(input_fmap_4[7:0]),.cy( 9'sd1),.dx(input_fmap_7[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O55_N0_S1),.chainout(chainout_0_O55));
logic signed [63:0] chainout_2_O55; 
logic signed [63:0] O55_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O55(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_10[7:0]),.ay(-9'sd1),.bx(input_fmap_14[7:0]),.by( 9'sd1),.cx(input_fmap_17[7:0]),.cy( 9'sd1),.dx(input_fmap_20[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O55_N2_S1),.chainout(chainout_2_O55));
logic signed [63:0] chainout_4_O55; 
logic signed [63:0] O55_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O55(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_25[7:0]),.ay( 9'sd1),.bx(input_fmap_26[7:0]),.by(-9'sd1),.cx(input_fmap_27[7:0]),.cy(-9'sd1),.dx(input_fmap_30[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O55_N4_S1),.chainout(chainout_4_O55));
logic signed [63:0] chainout_6_O55; 
logic signed [63:0] O55_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O55(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_32[7:0]),.ay( 9'sd6),.bx(input_fmap_33[7:0]),.by( 9'sd1),.cx(input_fmap_35[7:0]),.cy(-9'sd1),.dx(input_fmap_36[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O55_N6_S1),.chainout(chainout_6_O55));
logic signed [63:0] chainout_8_O55; 
logic signed [63:0] O55_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O55(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_37[7:0]),.ay(-9'sd1),.bx(input_fmap_38[7:0]),.by(-9'sd1),.cx(input_fmap_42[7:0]),.cy(-9'sd1),.dx(input_fmap_43[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O55_N8_S1),.chainout(chainout_8_O55));
logic signed [63:0] chainout_10_O55; 
logic signed [63:0] O55_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O55(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_46[7:0]),.ay( 9'sd1),.bx(input_fmap_54[7:0]),.by(-9'sd1),.cx(input_fmap_57[7:0]),.cy( 9'sd1),.dx(input_fmap_58[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O55_N10_S1),.chainout(chainout_10_O55));
logic signed [63:0] chainout_12_O55; 
logic signed [63:0] O55_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O55(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_61[7:0]),.ay(-9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O55_N12_S1),.chainout(chainout_12_O55));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O55_N0_S2;		always @(posedge clk) O55_N0_S2 <=     O55_N0_S1  +  O55_N2_S1 ;
 logic signed [21:0] O55_N2_S2;		always @(posedge clk) O55_N2_S2 <=     O55_N4_S1  +  O55_N6_S1 ;
 logic signed [21:0] O55_N4_S2;		always @(posedge clk) O55_N4_S2 <=     O55_N8_S1  +  O55_N10_S1 ;
 logic signed [21:0] O55_N6_S2;		always @(posedge clk) O55_N6_S2 <=     O55_N12_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O55_N0_S3;		always @(posedge clk) O55_N0_S3 <=     O55_N0_S2  +  O55_N2_S2 ;
 logic signed [22:0] O55_N2_S3;		always @(posedge clk) O55_N2_S3 <=     O55_N4_S2  +  O55_N6_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O55_N0_S4;		always @(posedge clk) O55_N0_S4 <=     O55_N0_S3  +  O55_N2_S3 ;
 assign conv_mac_55 = O55_N0_S4;

logic signed [31:0] conv_mac_56;
logic signed [63:0] chainout_0_O56; 
logic signed [63:0] O56_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O56(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_5[7:0]),.ay(-9'sd1),.bx(input_fmap_6[7:0]),.by( 9'sd1),.cx(input_fmap_10[7:0]),.cy( 9'sd1),.dx(input_fmap_12[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O56_N0_S1),.chainout(chainout_0_O56));
logic signed [63:0] chainout_2_O56; 
logic signed [63:0] O56_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O56(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_13[7:0]),.ay( 9'sd1),.bx(input_fmap_14[7:0]),.by( 9'sd1),.cx(input_fmap_15[7:0]),.cy( 9'sd1),.dx(input_fmap_16[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O56_N2_S1),.chainout(chainout_2_O56));
logic signed [63:0] chainout_4_O56; 
logic signed [63:0] O56_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O56(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_17[7:0]),.ay(-9'sd1),.bx(input_fmap_18[7:0]),.by( 9'sd1),.cx(input_fmap_21[7:0]),.cy( 9'sd4),.dx(input_fmap_26[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O56_N4_S1),.chainout(chainout_4_O56));
logic signed [63:0] chainout_6_O56; 
logic signed [63:0] O56_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O56(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_27[7:0]),.ay( 9'sd1),.bx(input_fmap_29[7:0]),.by( 9'sd1),.cx(input_fmap_34[7:0]),.cy(-9'sd1),.dx(input_fmap_36[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O56_N6_S1),.chainout(chainout_6_O56));
logic signed [63:0] chainout_8_O56; 
logic signed [63:0] O56_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O56(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_37[7:0]),.ay(-9'sd1),.bx(input_fmap_40[7:0]),.by( 9'sd1),.cx(input_fmap_41[7:0]),.cy(-9'sd1),.dx(input_fmap_42[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O56_N8_S1),.chainout(chainout_8_O56));
logic signed [63:0] chainout_10_O56; 
logic signed [63:0] O56_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O56(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_45[7:0]),.ay(-9'sd1),.bx(input_fmap_47[7:0]),.by( 9'sd1),.cx(input_fmap_54[7:0]),.cy(-9'sd1),.dx(input_fmap_60[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O56_N10_S1),.chainout(chainout_10_O56));
logic signed [63:0] chainout_12_O56; 
logic signed [63:0] O56_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O56(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_63[7:0]),.ay( 9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O56_N12_S1),.chainout(chainout_12_O56));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O56_N0_S2;		always @(posedge clk) O56_N0_S2 <=     O56_N0_S1  +  O56_N2_S1 ;
 logic signed [21:0] O56_N2_S2;		always @(posedge clk) O56_N2_S2 <=     O56_N4_S1  +  O56_N6_S1 ;
 logic signed [21:0] O56_N4_S2;		always @(posedge clk) O56_N4_S2 <=     O56_N8_S1  +  O56_N10_S1 ;
 logic signed [21:0] O56_N6_S2;		always @(posedge clk) O56_N6_S2 <=     O56_N12_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O56_N0_S3;		always @(posedge clk) O56_N0_S3 <=     O56_N0_S2  +  O56_N2_S2 ;
 logic signed [22:0] O56_N2_S3;		always @(posedge clk) O56_N2_S3 <=     O56_N4_S2  +  O56_N6_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O56_N0_S4;		always @(posedge clk) O56_N0_S4 <=     O56_N0_S3  +  O56_N2_S3 ;
 assign conv_mac_56 = O56_N0_S4;

logic signed [31:0] conv_mac_57;
logic signed [63:0] chainout_0_O57; 
logic signed [63:0] O57_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O57(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay(-9'sd2),.bx(input_fmap_3[7:0]),.by(-9'sd1),.cx(input_fmap_4[7:0]),.cy(-9'sd1),.dx(input_fmap_5[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O57_N0_S1),.chainout(chainout_0_O57));
logic signed [63:0] chainout_2_O57; 
logic signed [63:0] O57_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O57(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_9[7:0]),.ay( 9'sd2),.bx(input_fmap_10[7:0]),.by(-9'sd1),.cx(input_fmap_17[7:0]),.cy( 9'sd1),.dx(input_fmap_19[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O57_N2_S1),.chainout(chainout_2_O57));
logic signed [63:0] chainout_4_O57; 
logic signed [63:0] O57_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O57(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_21[7:0]),.ay( 9'sd1),.bx(input_fmap_22[7:0]),.by(-9'sd1),.cx(input_fmap_23[7:0]),.cy( 9'sd1),.dx(input_fmap_26[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O57_N4_S1),.chainout(chainout_4_O57));
logic signed [63:0] chainout_6_O57; 
logic signed [63:0] O57_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O57(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_27[7:0]),.ay( 9'sd2),.bx(input_fmap_28[7:0]),.by( 9'sd1),.cx(input_fmap_29[7:0]),.cy( 9'sd1),.dx(input_fmap_31[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O57_N6_S1),.chainout(chainout_6_O57));
logic signed [63:0] chainout_8_O57; 
logic signed [63:0] O57_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O57(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_36[7:0]),.ay(-9'sd1),.bx(input_fmap_38[7:0]),.by( 9'sd1),.cx(input_fmap_40[7:0]),.cy(-9'sd1),.dx(input_fmap_43[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O57_N8_S1),.chainout(chainout_8_O57));
logic signed [63:0] chainout_10_O57; 
logic signed [63:0] O57_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O57(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_44[7:0]),.ay( 9'sd1),.bx(input_fmap_46[7:0]),.by( 9'sd1),.cx(input_fmap_47[7:0]),.cy(-9'sd2),.dx(input_fmap_50[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O57_N10_S1),.chainout(chainout_10_O57));
logic signed [63:0] chainout_12_O57; 
logic signed [63:0] O57_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O57(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_51[7:0]),.ay(-9'sd1),.bx(input_fmap_54[7:0]),.by( 9'sd1),.cx(input_fmap_57[7:0]),.cy( 9'sd1),.dx(input_fmap_58[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O57_N12_S1),.chainout(chainout_12_O57));
logic signed [63:0] chainout_14_O57; 
logic signed [63:0] O57_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O57(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_60[7:0]),.ay( 9'sd1),.bx(input_fmap_62[7:0]),.by( 9'sd1),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O57_N14_S1),.chainout(chainout_14_O57));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O57_N0_S2;		always @(posedge clk) O57_N0_S2 <=     O57_N0_S1  +  O57_N2_S1 ;
 logic signed [21:0] O57_N2_S2;		always @(posedge clk) O57_N2_S2 <=     O57_N4_S1  +  O57_N6_S1 ;
 logic signed [21:0] O57_N4_S2;		always @(posedge clk) O57_N4_S2 <=     O57_N8_S1  +  O57_N10_S1 ;
 logic signed [21:0] O57_N6_S2;		always @(posedge clk) O57_N6_S2 <=     O57_N12_S1  +  O57_N14_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O57_N0_S3;		always @(posedge clk) O57_N0_S3 <=     O57_N0_S2  +  O57_N2_S2 ;
 logic signed [22:0] O57_N2_S3;		always @(posedge clk) O57_N2_S3 <=     O57_N4_S2  +  O57_N6_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O57_N0_S4;		always @(posedge clk) O57_N0_S4 <=     O57_N0_S3  +  O57_N2_S3 ;
 assign conv_mac_57 = O57_N0_S4;

logic signed [31:0] conv_mac_58;
logic signed [63:0] chainout_0_O58; 
logic signed [63:0] O58_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O58(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay(-9'sd1),.bx(input_fmap_3[7:0]),.by( 9'sd2),.cx(input_fmap_4[7:0]),.cy(-9'sd2),.dx(input_fmap_5[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O58_N0_S1),.chainout(chainout_0_O58));
logic signed [63:0] chainout_2_O58; 
logic signed [63:0] O58_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O58(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_7[7:0]),.ay(-9'sd1),.bx(input_fmap_8[7:0]),.by( 9'sd1),.cx(input_fmap_9[7:0]),.cy( 9'sd1),.dx(input_fmap_10[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O58_N2_S1),.chainout(chainout_2_O58));
logic signed [63:0] chainout_4_O58; 
logic signed [63:0] O58_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O58(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_12[7:0]),.ay( 9'sd1),.bx(input_fmap_13[7:0]),.by( 9'sd1),.cx(input_fmap_17[7:0]),.cy(-9'sd1),.dx(input_fmap_18[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O58_N4_S1),.chainout(chainout_4_O58));
logic signed [63:0] chainout_6_O58; 
logic signed [63:0] O58_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O58(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_19[7:0]),.ay(-9'sd4),.bx(input_fmap_20[7:0]),.by( 9'sd2),.cx(input_fmap_23[7:0]),.cy( 9'sd2),.dx(input_fmap_24[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O58_N6_S1),.chainout(chainout_6_O58));
logic signed [63:0] chainout_8_O58; 
logic signed [63:0] O58_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O58(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_25[7:0]),.ay(-9'sd2),.bx(input_fmap_26[7:0]),.by( 9'sd1),.cx(input_fmap_27[7:0]),.cy( 9'sd1),.dx(input_fmap_28[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O58_N8_S1),.chainout(chainout_8_O58));
logic signed [63:0] chainout_10_O58; 
logic signed [63:0] O58_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O58(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_29[7:0]),.ay(-9'sd2),.bx(input_fmap_30[7:0]),.by(-9'sd2),.cx(input_fmap_32[7:0]),.cy( 9'sd1),.dx(input_fmap_33[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O58_N10_S1),.chainout(chainout_10_O58));
logic signed [63:0] chainout_12_O58; 
logic signed [63:0] O58_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O58(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_36[7:0]),.ay(-9'sd1),.bx(input_fmap_37[7:0]),.by(-9'sd3),.cx(input_fmap_38[7:0]),.cy( 9'sd4),.dx(input_fmap_41[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O58_N12_S1),.chainout(chainout_12_O58));
logic signed [63:0] chainout_14_O58; 
logic signed [63:0] O58_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O58(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_42[7:0]),.ay( 9'sd1),.bx(input_fmap_44[7:0]),.by( 9'sd2),.cx(input_fmap_45[7:0]),.cy( 9'sd2),.dx(input_fmap_46[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O58_N14_S1),.chainout(chainout_14_O58));
logic signed [63:0] chainout_16_O58; 
logic signed [63:0] O58_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O58(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_48[7:0]),.ay(-9'sd1),.bx(input_fmap_49[7:0]),.by(-9'sd1),.cx(input_fmap_50[7:0]),.cy(-9'sd1),.dx(input_fmap_52[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O58_N16_S1),.chainout(chainout_16_O58));
logic signed [63:0] chainout_18_O58; 
logic signed [63:0] O58_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O58(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_53[7:0]),.ay( 9'sd1),.bx(input_fmap_55[7:0]),.by( 9'sd1),.cx(input_fmap_56[7:0]),.cy( 9'sd2),.dx(input_fmap_57[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O58_N18_S1),.chainout(chainout_18_O58));
logic signed [63:0] chainout_20_O58; 
logic signed [63:0] O58_N20_S1; 
 int_sop_4_wrapper int_sop_4_inst_20_O58(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_58[7:0]),.ay( 9'sd1),.bx(input_fmap_59[7:0]),.by( 9'sd1),.cx(input_fmap_62[7:0]),.cy( 9'sd1),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O58_N20_S1),.chainout(chainout_20_O58));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O58_N0_S2;		always @(posedge clk) O58_N0_S2 <=     O58_N0_S1  +  O58_N2_S1 ;
 logic signed [21:0] O58_N2_S2;		always @(posedge clk) O58_N2_S2 <=     O58_N4_S1  +  O58_N6_S1 ;
 logic signed [21:0] O58_N4_S2;		always @(posedge clk) O58_N4_S2 <=     O58_N8_S1  +  O58_N10_S1 ;
 logic signed [21:0] O58_N6_S2;		always @(posedge clk) O58_N6_S2 <=     O58_N12_S1  +  O58_N14_S1 ;
 logic signed [21:0] O58_N8_S2;		always @(posedge clk) O58_N8_S2 <=     O58_N16_S1  +  O58_N18_S1 ;
 logic signed [21:0] O58_N10_S2;		always @(posedge clk) O58_N10_S2 <=     O58_N20_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O58_N0_S3;		always @(posedge clk) O58_N0_S3 <=     O58_N0_S2  +  O58_N2_S2 ;
 logic signed [22:0] O58_N2_S3;		always @(posedge clk) O58_N2_S3 <=     O58_N4_S2  +  O58_N6_S2 ;
 logic signed [22:0] O58_N4_S3;		always @(posedge clk) O58_N4_S3 <=     O58_N8_S2  +  O58_N10_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O58_N0_S4;		always @(posedge clk) O58_N0_S4 <=     O58_N0_S3  +  O58_N2_S3 ;
 logic signed [23:0] O58_N2_S4;		always @(posedge clk) O58_N2_S4 <=     O58_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O58_N0_S5;		always @(posedge clk) O58_N0_S5 <=     O58_N0_S4  +  O58_N2_S4 ;
 assign conv_mac_58 = O58_N0_S5;

logic signed [31:0] conv_mac_59;
logic signed [63:0] chainout_0_O59; 
logic signed [63:0] O59_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O59(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_2[7:0]),.ay(-9'sd2),.bx(input_fmap_3[7:0]),.by(-9'sd2),.cx(input_fmap_5[7:0]),.cy( 9'sd2),.dx(input_fmap_7[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O59_N0_S1),.chainout(chainout_0_O59));
logic signed [63:0] chainout_2_O59; 
logic signed [63:0] O59_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O59(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_8[7:0]),.ay(-9'sd1),.bx(input_fmap_9[7:0]),.by(-9'sd1),.cx(input_fmap_10[7:0]),.cy(-9'sd1),.dx(input_fmap_12[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O59_N2_S1),.chainout(chainout_2_O59));
logic signed [63:0] chainout_4_O59; 
logic signed [63:0] O59_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O59(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_16[7:0]),.ay(-9'sd1),.bx(input_fmap_18[7:0]),.by( 9'sd1),.cx(input_fmap_19[7:0]),.cy(-9'sd1),.dx(input_fmap_21[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O59_N4_S1),.chainout(chainout_4_O59));
logic signed [63:0] chainout_6_O59; 
logic signed [63:0] O59_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O59(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_22[7:0]),.ay(-9'sd1),.bx(input_fmap_23[7:0]),.by( 9'sd1),.cx(input_fmap_25[7:0]),.cy( 9'sd1),.dx(input_fmap_27[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O59_N6_S1),.chainout(chainout_6_O59));
logic signed [63:0] chainout_8_O59; 
logic signed [63:0] O59_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O59(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_31[7:0]),.ay(-9'sd1),.bx(input_fmap_32[7:0]),.by(-9'sd1),.cx(input_fmap_35[7:0]),.cy(-9'sd1),.dx(input_fmap_36[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O59_N8_S1),.chainout(chainout_8_O59));
logic signed [63:0] chainout_10_O59; 
logic signed [63:0] O59_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O59(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_42[7:0]),.ay( 9'sd1),.bx(input_fmap_43[7:0]),.by(-9'sd2),.cx(input_fmap_44[7:0]),.cy(-9'sd1),.dx(input_fmap_47[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O59_N10_S1),.chainout(chainout_10_O59));
logic signed [63:0] chainout_12_O59; 
logic signed [63:0] O59_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O59(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_49[7:0]),.ay( 9'sd1),.bx(input_fmap_51[7:0]),.by( 9'sd1),.cx(input_fmap_55[7:0]),.cy(-9'sd1),.dx(input_fmap_56[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O59_N12_S1),.chainout(chainout_12_O59));
logic signed [63:0] chainout_14_O59; 
logic signed [63:0] O59_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O59(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_57[7:0]),.ay(-9'sd1),.bx(input_fmap_60[7:0]),.by( 9'sd1),.cx(input_fmap_61[7:0]),.cy(-9'sd1),.dx(input_fmap_62[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O59_N14_S1),.chainout(chainout_14_O59));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O59_N0_S2;		always @(posedge clk) O59_N0_S2 <=     O59_N0_S1  +  O59_N2_S1 ;
 logic signed [21:0] O59_N2_S2;		always @(posedge clk) O59_N2_S2 <=     O59_N4_S1  +  O59_N6_S1 ;
 logic signed [21:0] O59_N4_S2;		always @(posedge clk) O59_N4_S2 <=     O59_N8_S1  +  O59_N10_S1 ;
 logic signed [21:0] O59_N6_S2;		always @(posedge clk) O59_N6_S2 <=     O59_N12_S1  +  O59_N14_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O59_N0_S3;		always @(posedge clk) O59_N0_S3 <=     O59_N0_S2  +  O59_N2_S2 ;
 logic signed [22:0] O59_N2_S3;		always @(posedge clk) O59_N2_S3 <=     O59_N4_S2  +  O59_N6_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O59_N0_S4;		always @(posedge clk) O59_N0_S4 <=     O59_N0_S3  +  O59_N2_S3 ;
 assign conv_mac_59 = O59_N0_S4;

logic signed [31:0] conv_mac_60;
logic signed [63:0] chainout_0_O60; 
logic signed [63:0] O60_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O60(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay( 9'sd1),.bx(input_fmap_3[7:0]),.by(-9'sd1),.cx(input_fmap_4[7:0]),.cy( 9'sd2),.dx(input_fmap_5[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O60_N0_S1),.chainout(chainout_0_O60));
logic signed [63:0] chainout_2_O60; 
logic signed [63:0] O60_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O60(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_6[7:0]),.ay( 9'sd2),.bx(input_fmap_7[7:0]),.by(-9'sd3),.cx(input_fmap_8[7:0]),.cy( 9'sd1),.dx(input_fmap_9[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O60_N2_S1),.chainout(chainout_2_O60));
logic signed [63:0] chainout_4_O60; 
logic signed [63:0] O60_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O60(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_10[7:0]),.ay(-9'sd1),.bx(input_fmap_11[7:0]),.by( 9'sd2),.cx(input_fmap_12[7:0]),.cy( 9'sd1),.dx(input_fmap_14[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O60_N4_S1),.chainout(chainout_4_O60));
logic signed [63:0] chainout_6_O60; 
logic signed [63:0] O60_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O60(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_15[7:0]),.ay(-9'sd1),.bx(input_fmap_18[7:0]),.by(-9'sd1),.cx(input_fmap_24[7:0]),.cy(-9'sd1),.dx(input_fmap_25[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O60_N6_S1),.chainout(chainout_6_O60));
logic signed [63:0] chainout_8_O60; 
logic signed [63:0] O60_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O60(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_30[7:0]),.ay( 9'sd1),.bx(input_fmap_31[7:0]),.by( 9'sd1),.cx(input_fmap_32[7:0]),.cy( 9'sd1),.dx(input_fmap_34[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O60_N8_S1),.chainout(chainout_8_O60));
logic signed [63:0] chainout_10_O60; 
logic signed [63:0] O60_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O60(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_35[7:0]),.ay(-9'sd2),.bx(input_fmap_36[7:0]),.by(-9'sd1),.cx(input_fmap_37[7:0]),.cy(-9'sd1),.dx(input_fmap_38[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O60_N10_S1),.chainout(chainout_10_O60));
logic signed [63:0] chainout_12_O60; 
logic signed [63:0] O60_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O60(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_39[7:0]),.ay( 9'sd2),.bx(input_fmap_40[7:0]),.by(-9'sd1),.cx(input_fmap_43[7:0]),.cy( 9'sd2),.dx(input_fmap_44[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O60_N12_S1),.chainout(chainout_12_O60));
logic signed [63:0] chainout_14_O60; 
logic signed [63:0] O60_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O60(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_45[7:0]),.ay( 9'sd1),.bx(input_fmap_46[7:0]),.by( 9'sd1),.cx(input_fmap_47[7:0]),.cy(-9'sd1),.dx(input_fmap_48[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O60_N14_S1),.chainout(chainout_14_O60));
logic signed [63:0] chainout_16_O60; 
logic signed [63:0] O60_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O60(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_50[7:0]),.ay( 9'sd1),.bx(input_fmap_51[7:0]),.by(-9'sd2),.cx(input_fmap_52[7:0]),.cy(-9'sd2),.dx(input_fmap_54[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O60_N16_S1),.chainout(chainout_16_O60));
logic signed [63:0] chainout_18_O60; 
logic signed [63:0] O60_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O60(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_55[7:0]),.ay(-9'sd1),.bx(input_fmap_56[7:0]),.by(-9'sd1),.cx(input_fmap_59[7:0]),.cy( 9'sd2),.dx(input_fmap_61[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O60_N18_S1),.chainout(chainout_18_O60));
logic signed [63:0] chainout_20_O60; 
logic signed [63:0] O60_N20_S1; 
 int_sop_4_wrapper int_sop_4_inst_20_O60(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_63[7:0]),.ay(-9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O60_N20_S1),.chainout(chainout_20_O60));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O60_N0_S2;		always @(posedge clk) O60_N0_S2 <=     O60_N0_S1  +  O60_N2_S1 ;
 logic signed [21:0] O60_N2_S2;		always @(posedge clk) O60_N2_S2 <=     O60_N4_S1  +  O60_N6_S1 ;
 logic signed [21:0] O60_N4_S2;		always @(posedge clk) O60_N4_S2 <=     O60_N8_S1  +  O60_N10_S1 ;
 logic signed [21:0] O60_N6_S2;		always @(posedge clk) O60_N6_S2 <=     O60_N12_S1  +  O60_N14_S1 ;
 logic signed [21:0] O60_N8_S2;		always @(posedge clk) O60_N8_S2 <=     O60_N16_S1  +  O60_N18_S1 ;
 logic signed [21:0] O60_N10_S2;		always @(posedge clk) O60_N10_S2 <=     O60_N20_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O60_N0_S3;		always @(posedge clk) O60_N0_S3 <=     O60_N0_S2  +  O60_N2_S2 ;
 logic signed [22:0] O60_N2_S3;		always @(posedge clk) O60_N2_S3 <=     O60_N4_S2  +  O60_N6_S2 ;
 logic signed [22:0] O60_N4_S3;		always @(posedge clk) O60_N4_S3 <=     O60_N8_S2  +  O60_N10_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O60_N0_S4;		always @(posedge clk) O60_N0_S4 <=     O60_N0_S3  +  O60_N2_S3 ;
 logic signed [23:0] O60_N2_S4;		always @(posedge clk) O60_N2_S4 <=     O60_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O60_N0_S5;		always @(posedge clk) O60_N0_S5 <=     O60_N0_S4  +  O60_N2_S4 ;
 assign conv_mac_60 = O60_N0_S5;

logic signed [31:0] conv_mac_61;
logic signed [63:0] chainout_0_O61; 
logic signed [63:0] O61_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O61(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_0[7:0]),.ay( 9'sd2),.bx(input_fmap_2[7:0]),.by(-9'sd2),.cx(input_fmap_3[7:0]),.cy(-9'sd1),.dx(input_fmap_5[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O61_N0_S1),.chainout(chainout_0_O61));
logic signed [63:0] chainout_2_O61; 
logic signed [63:0] O61_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O61(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_6[7:0]),.ay( 9'sd1),.bx(input_fmap_8[7:0]),.by(-9'sd1),.cx(input_fmap_9[7:0]),.cy( 9'sd1),.dx(input_fmap_12[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O61_N2_S1),.chainout(chainout_2_O61));
logic signed [63:0] chainout_4_O61; 
logic signed [63:0] O61_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O61(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_13[7:0]),.ay( 9'sd1),.bx(input_fmap_14[7:0]),.by( 9'sd5),.cx(input_fmap_15[7:0]),.cy( 9'sd3),.dx(input_fmap_16[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O61_N4_S1),.chainout(chainout_4_O61));
logic signed [63:0] chainout_6_O61; 
logic signed [63:0] O61_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O61(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_18[7:0]),.ay( 9'sd1),.bx(input_fmap_19[7:0]),.by(-9'sd1),.cx(input_fmap_20[7:0]),.cy( 9'sd1),.dx(input_fmap_22[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O61_N6_S1),.chainout(chainout_6_O61));
logic signed [63:0] chainout_8_O61; 
logic signed [63:0] O61_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O61(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_23[7:0]),.ay(-9'sd1),.bx(input_fmap_24[7:0]),.by( 9'sd1),.cx(input_fmap_25[7:0]),.cy(-9'sd1),.dx(input_fmap_26[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O61_N8_S1),.chainout(chainout_8_O61));
logic signed [63:0] chainout_10_O61; 
logic signed [63:0] O61_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O61(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_27[7:0]),.ay( 9'sd1),.bx(input_fmap_28[7:0]),.by( 9'sd2),.cx(input_fmap_31[7:0]),.cy( 9'sd2),.dx(input_fmap_34[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O61_N10_S1),.chainout(chainout_10_O61));
logic signed [63:0] chainout_12_O61; 
logic signed [63:0] O61_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O61(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_35[7:0]),.ay(-9'sd1),.bx(input_fmap_36[7:0]),.by(-9'sd2),.cx(input_fmap_38[7:0]),.cy(-9'sd1),.dx(input_fmap_39[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O61_N12_S1),.chainout(chainout_12_O61));
logic signed [63:0] chainout_14_O61; 
logic signed [63:0] O61_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O61(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_40[7:0]),.ay( 9'sd1),.bx(input_fmap_41[7:0]),.by(-9'sd2),.cx(input_fmap_42[7:0]),.cy( 9'sd2),.dx(input_fmap_43[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O61_N14_S1),.chainout(chainout_14_O61));
logic signed [63:0] chainout_16_O61; 
logic signed [63:0] O61_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O61(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_44[7:0]),.ay( 9'sd1),.bx(input_fmap_46[7:0]),.by( 9'sd2),.cx(input_fmap_47[7:0]),.cy( 9'sd1),.dx(input_fmap_48[7:0]),.dy(-9'sd3),.chainin(63'd0),.result(O61_N16_S1),.chainout(chainout_16_O61));
logic signed [63:0] chainout_18_O61; 
logic signed [63:0] O61_N18_S1; 
 int_sop_4_wrapper int_sop_4_inst_18_O61(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_50[7:0]),.ay( 9'sd1),.bx(input_fmap_52[7:0]),.by( 9'sd1),.cx(input_fmap_53[7:0]),.cy(-9'sd4),.dx(input_fmap_54[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O61_N18_S1),.chainout(chainout_18_O61));
logic signed [63:0] chainout_20_O61; 
logic signed [63:0] O61_N20_S1; 
 int_sop_4_wrapper int_sop_4_inst_20_O61(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_55[7:0]),.ay( 9'sd1),.bx(input_fmap_56[7:0]),.by( 9'sd2),.cx(input_fmap_57[7:0]),.cy(-9'sd1),.dx(input_fmap_59[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O61_N20_S1),.chainout(chainout_20_O61));
logic signed [63:0] chainout_22_O61; 
logic signed [63:0] O61_N22_S1; 
 int_sop_4_wrapper int_sop_4_inst_22_O61(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_61[7:0]),.ay(-9'sd1),.bx(input_fmap_62[7:0]),.by(-9'sd1),.cx(input_fmap_63[7:0]),.cy( 9'sd1),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O61_N22_S1),.chainout(chainout_22_O61));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O61_N0_S2;		always @(posedge clk) O61_N0_S2 <=     O61_N0_S1  +  O61_N2_S1 ;
 logic signed [21:0] O61_N2_S2;		always @(posedge clk) O61_N2_S2 <=     O61_N4_S1  +  O61_N6_S1 ;
 logic signed [21:0] O61_N4_S2;		always @(posedge clk) O61_N4_S2 <=     O61_N8_S1  +  O61_N10_S1 ;
 logic signed [21:0] O61_N6_S2;		always @(posedge clk) O61_N6_S2 <=     O61_N12_S1  +  O61_N14_S1 ;
 logic signed [21:0] O61_N8_S2;		always @(posedge clk) O61_N8_S2 <=     O61_N16_S1  +  O61_N18_S1 ;
 logic signed [21:0] O61_N10_S2;		always @(posedge clk) O61_N10_S2 <=     O61_N20_S1  +  O61_N22_S1 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O61_N0_S3;		always @(posedge clk) O61_N0_S3 <=     O61_N0_S2  +  O61_N2_S2 ;
 logic signed [22:0] O61_N2_S3;		always @(posedge clk) O61_N2_S3 <=     O61_N4_S2  +  O61_N6_S2 ;
 logic signed [22:0] O61_N4_S3;		always @(posedge clk) O61_N4_S3 <=     O61_N8_S2  +  O61_N10_S2 ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O61_N0_S4;		always @(posedge clk) O61_N0_S4 <=     O61_N0_S3  +  O61_N2_S3 ;
 logic signed [23:0] O61_N2_S4;		always @(posedge clk) O61_N2_S4 <=     O61_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O61_N0_S5;		always @(posedge clk) O61_N0_S5 <=     O61_N0_S4  +  O61_N2_S4 ;
 assign conv_mac_61 = O61_N0_S5;

logic signed [31:0] conv_mac_62;
logic signed [63:0] chainout_0_O62; 
logic signed [63:0] O62_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O62(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_5[7:0]),.ay( 9'sd1),.bx(input_fmap_6[7:0]),.by(-9'sd1),.cx(input_fmap_15[7:0]),.cy( 9'sd1),.dx(input_fmap_25[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O62_N0_S1),.chainout(chainout_0_O62));
logic signed [63:0] chainout_2_O62; 
logic signed [63:0] O62_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O62(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_31[7:0]),.ay( 9'sd1),.bx(input_fmap_40[7:0]),.by( 9'sd1),.cx(input_fmap_41[7:0]),.cy( 9'sd1),.dx(input_fmap_45[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O62_N2_S1),.chainout(chainout_2_O62));
logic signed [63:0] chainout_4_O62; 
logic signed [63:0] O62_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O62(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_50[7:0]),.ay( 9'sd1),.bx(input_fmap_51[7:0]),.by(-9'sd1),.cx(input_fmap_56[7:0]),.cy( 9'sd1),.dx(input_fmap_61[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O62_N4_S1),.chainout(chainout_4_O62));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O62_N0_S2;		always @(posedge clk) O62_N0_S2 <=     O62_N0_S1  +  O62_N2_S1 ;
 logic signed [21:0] O62_N2_S2;		always @(posedge clk) O62_N2_S2 <=     O62_N4_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O62_N0_S3;		always @(posedge clk) O62_N0_S3 <=     O62_N0_S2  +  O62_N2_S2 ;
 assign conv_mac_62 = O62_N0_S3;

logic signed [31:0] conv_mac_63;
logic signed [63:0] chainout_0_O63; 
logic signed [63:0] O63_N0_S1; 
 int_sop_4_wrapper int_sop_4_inst_0_O63(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_1[7:0]),.ay( 9'sd1),.bx(input_fmap_4[7:0]),.by(-9'sd1),.cx(input_fmap_8[7:0]),.cy(-9'sd1),.dx(input_fmap_12[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O63_N0_S1),.chainout(chainout_0_O63));
logic signed [63:0] chainout_2_O63; 
logic signed [63:0] O63_N2_S1; 
 int_sop_4_wrapper int_sop_4_inst_2_O63(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_15[7:0]),.ay( 9'sd1),.bx(input_fmap_16[7:0]),.by(-9'sd1),.cx(input_fmap_18[7:0]),.cy( 9'sd1),.dx(input_fmap_19[7:0]),.dy(-9'sd2),.chainin(63'd0),.result(O63_N2_S1),.chainout(chainout_2_O63));
logic signed [63:0] chainout_4_O63; 
logic signed [63:0] O63_N4_S1; 
 int_sop_4_wrapper int_sop_4_inst_4_O63(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_23[7:0]),.ay( 9'sd1),.bx(input_fmap_25[7:0]),.by( 9'sd2),.cx(input_fmap_26[7:0]),.cy(-9'sd1),.dx(input_fmap_27[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O63_N4_S1),.chainout(chainout_4_O63));
logic signed [63:0] chainout_6_O63; 
logic signed [63:0] O63_N6_S1; 
 int_sop_4_wrapper int_sop_4_inst_6_O63(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_28[7:0]),.ay( 9'sd1),.bx(input_fmap_29[7:0]),.by(-9'sd1),.cx(input_fmap_33[7:0]),.cy(-9'sd1),.dx(input_fmap_35[7:0]),.dy( 9'sd2),.chainin(63'd0),.result(O63_N6_S1),.chainout(chainout_6_O63));
logic signed [63:0] chainout_8_O63; 
logic signed [63:0] O63_N8_S1; 
 int_sop_4_wrapper int_sop_4_inst_8_O63(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_37[7:0]),.ay(-9'sd1),.bx(input_fmap_41[7:0]),.by(-9'sd1),.cx(input_fmap_42[7:0]),.cy( 9'sd1),.dx(input_fmap_43[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O63_N8_S1),.chainout(chainout_8_O63));
logic signed [63:0] chainout_10_O63; 
logic signed [63:0] O63_N10_S1; 
 int_sop_4_wrapper int_sop_4_inst_10_O63(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_45[7:0]),.ay( 9'sd2),.bx(input_fmap_46[7:0]),.by( 9'sd1),.cx(input_fmap_47[7:0]),.cy( 9'sd1),.dx(input_fmap_48[7:0]),.dy(-9'sd1),.chainin(63'd0),.result(O63_N10_S1),.chainout(chainout_10_O63));
logic signed [63:0] chainout_12_O63; 
logic signed [63:0] O63_N12_S1; 
 int_sop_4_wrapper int_sop_4_inst_12_O63(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_50[7:0]),.ay(-9'sd1),.bx(input_fmap_51[7:0]),.by( 9'sd3),.cx(input_fmap_54[7:0]),.cy( 9'sd1),.dx(input_fmap_55[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O63_N12_S1),.chainout(chainout_12_O63));
logic signed [63:0] chainout_14_O63; 
logic signed [63:0] O63_N14_S1; 
 int_sop_4_wrapper int_sop_4_inst_14_O63(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_56[7:0]),.ay( 9'sd1),.bx(input_fmap_58[7:0]),.by( 9'sd1),.cx(input_fmap_59[7:0]),.cy(-9'sd1),.dx(input_fmap_60[7:0]),.dy( 9'sd1),.chainin(63'd0),.result(O63_N14_S1),.chainout(chainout_14_O63));
logic signed [63:0] chainout_16_O63; 
logic signed [63:0] O63_N16_S1; 
 int_sop_4_wrapper int_sop_4_inst_16_O63(.clk(clk),.reset(rstn),.mode_sigs(12'd0),.ax(input_fmap_61[7:0]),.ay( 9'sd1),.bx(zero_number[8:0]),.by( 9'sd0),.cx(zero_number[8:0]),.cy( 9'sd0),.dx(zero_number[8:0]),.dy( 9'sd0),.chainin(63'd0),.result(O63_N16_S1),.chainout(chainout_16_O63));
//----------------------adder tree stage complete--------------------------------//
//----------------------adder tree stage complete--------------------------------//
logic signed [21:0] O63_N0_S2;		always @(posedge clk) O63_N0_S2 <=     O63_N0_S1  +  O63_N2_S1 ;
 logic signed [21:0] O63_N2_S2;		always @(posedge clk) O63_N2_S2 <=     O63_N4_S1  +  O63_N6_S1 ;
 logic signed [21:0] O63_N4_S2;		always @(posedge clk) O63_N4_S2 <=     O63_N8_S1  +  O63_N10_S1 ;
 logic signed [21:0] O63_N6_S2;		always @(posedge clk) O63_N6_S2 <=     O63_N12_S1  +  O63_N14_S1 ;
 logic signed [21:0] O63_N8_S2;		always @(posedge clk) O63_N8_S2 <=     O63_N16_S1     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [22:0] O63_N0_S3;		always @(posedge clk) O63_N0_S3 <=     O63_N0_S2  +  O63_N2_S2 ;
 logic signed [22:0] O63_N2_S3;		always @(posedge clk) O63_N2_S3 <=     O63_N4_S2  +  O63_N6_S2 ;
 logic signed [22:0] O63_N4_S3;		always @(posedge clk) O63_N4_S3 <=     O63_N8_S2     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [23:0] O63_N0_S4;		always @(posedge clk) O63_N0_S4 <=     O63_N0_S3  +  O63_N2_S3 ;
 logic signed [23:0] O63_N2_S4;		always @(posedge clk) O63_N2_S4 <=     O63_N4_S3     ;
 //----------------------adder tree stage complete--------------------------------//
logic signed [24:0] O63_N0_S5;		always @(posedge clk) O63_N0_S5 <=     O63_N0_S4  +  O63_N2_S4 ;
 assign conv_mac_63 = O63_N0_S5;

logic valid_D1;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D1<= 0 ;
	else valid_D1<=valid;
end
logic valid_D2;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D2<= 0 ;
	else valid_D2<=valid_D1;
end
logic valid_D3;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D3<= 0 ;
	else valid_D3<=valid_D2;
end
logic valid_D4;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D4<= 0 ;
	else valid_D4<=valid_D3;
end
logic valid_D5;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D5<= 0 ;
	else valid_D5<=valid_D4;
end
logic valid_D6;
always_ff @(posedge clk) begin
	if (rstn == 0) valid_D6<= 0 ;
	else valid_D6<=valid_D5;
end
always_ff @(posedge clk) begin
	if (rstn == 0) ready <= 0 ;
	else ready <=valid_D6;
end
logic [31:0] bias_add_0;
assign bias_add_0 = conv_mac_0 + 4'd6;
logic [31:0] bias_add_1;
assign bias_add_1 = conv_mac_1 - 5'd11;
logic [31:0] bias_add_2;
assign bias_add_2 = conv_mac_2 - 3'd3;
logic [31:0] bias_add_3;
assign bias_add_3 = conv_mac_3 + 5'd8;
logic [31:0] bias_add_4;
assign bias_add_4 = conv_mac_4 + 5'd10;
logic [31:0] bias_add_5;
assign bias_add_5 = conv_mac_5 + 2'd1;
logic [31:0] bias_add_6;
assign bias_add_6 = conv_mac_6 - 4'd5;
logic [31:0] bias_add_7;
assign bias_add_7 = conv_mac_7 + 5'd9;
logic [31:0] bias_add_8;
assign bias_add_8 = conv_mac_8 + 4'd5;
logic [31:0] bias_add_9;
assign bias_add_9 = conv_mac_9 + 6'd20;
logic [31:0] bias_add_10;
assign bias_add_10 = conv_mac_10 + 3'd2;
logic [31:0] bias_add_11;
assign bias_add_11 = conv_mac_11 - 4'd7;
logic [31:0] bias_add_12;
assign bias_add_12 = conv_mac_12 + 4'd6;
logic [31:0] bias_add_13;
assign bias_add_13 = conv_mac_13 + 3'd3;
logic [31:0] bias_add_14;
assign bias_add_14 = conv_mac_14 + 6'd22;
logic [31:0] bias_add_15;
assign bias_add_15 = conv_mac_15 + 5'd11;
logic [31:0] bias_add_16;
assign bias_add_16 = conv_mac_16 - 3'd3;
logic [31:0] bias_add_17;
assign bias_add_17 = conv_mac_17 + 5'd11;
logic [31:0] bias_add_18;
assign bias_add_18 = conv_mac_18 + 4'd6;
logic [31:0] bias_add_19;
assign bias_add_19 = conv_mac_19 + 6'd18;
logic [31:0] bias_add_20;
assign bias_add_20 = conv_mac_20 + 3'd2;
logic [31:0] bias_add_21;
assign bias_add_21 = conv_mac_21 + 5'd14;
logic [31:0] bias_add_22;
assign bias_add_22 = conv_mac_22 + 4'd6;
logic [31:0] bias_add_23;
assign bias_add_23 = conv_mac_23 + 5'd13;
logic [31:0] bias_add_24;
assign bias_add_24 = conv_mac_24 + 5'd12;
logic [31:0] bias_add_25;
assign bias_add_25 = conv_mac_25 + 6'd18;
logic [31:0] bias_add_26;
assign bias_add_26 = conv_mac_26 + 6'd16;
logic [31:0] bias_add_27;
assign bias_add_27 = conv_mac_27 + 5'd8;
logic [31:0] bias_add_28;
assign bias_add_28 = conv_mac_28 + 3'd2;
logic [31:0] bias_add_29;
assign bias_add_29 = conv_mac_29 - 5'd10;
logic [31:0] bias_add_30;
assign bias_add_30 = conv_mac_30 + 3'd2;
logic [31:0] bias_add_31;
assign bias_add_31 = conv_mac_31 + 4'd4;
logic [31:0] bias_add_32;
assign bias_add_32 = conv_mac_32 + 5'd10;
logic [31:0] bias_add_33;
assign bias_add_33 = conv_mac_33 + 6'd21;
logic [31:0] bias_add_34;
assign bias_add_34 = conv_mac_34 + 5'd8;
logic [31:0] bias_add_35;
assign bias_add_35 = conv_mac_35 + 6'd16;
logic [31:0] bias_add_36;
assign bias_add_36 = conv_mac_36 + 6'd17;
logic [31:0] bias_add_37;
assign bias_add_37 = conv_mac_37 + 4'd6;
logic [31:0] bias_add_38;
assign bias_add_38 = conv_mac_38 + 5'd15;
logic [31:0] bias_add_39;
assign bias_add_39 = conv_mac_39 + 4'd4;
logic [31:0] bias_add_40;
assign bias_add_40 = conv_mac_40 + 4'd5;
logic [31:0] bias_add_41;
assign bias_add_41 = conv_mac_41 + 3'd2;
logic [31:0] bias_add_42;
assign bias_add_42 = conv_mac_42 + 4'd6;
logic [31:0] bias_add_43;
assign bias_add_43 = conv_mac_43 + 5'd8;
logic [31:0] bias_add_44;
assign bias_add_44 = conv_mac_44 + 5'd9;
logic [31:0] bias_add_45;
assign bias_add_45 = conv_mac_45 + 4'd5;
logic [31:0] bias_add_46;
assign bias_add_46 = conv_mac_46 + 4'd5;
logic [31:0] bias_add_47;
assign bias_add_47 = conv_mac_47 + 6'd18;
logic [31:0] bias_add_48;
assign bias_add_48 = conv_mac_48 + 6'd20;
logic [31:0] bias_add_49;
assign bias_add_49 = conv_mac_49 - 6'd16;
logic [31:0] bias_add_50;
assign bias_add_50 = conv_mac_50 + 4'd6;
logic [31:0] bias_add_51;
assign bias_add_51 = conv_mac_51 + 4'd4;
logic [31:0] bias_add_52;
assign bias_add_52 = conv_mac_52 + 4'd6;
logic [31:0] bias_add_53;
assign bias_add_53 = conv_mac_53 - 6'd17;
logic [31:0] bias_add_54;
assign bias_add_54 = conv_mac_54 + 4'd6;
logic [31:0] bias_add_55;
assign bias_add_55 = conv_mac_55 - 4'd4;
logic [31:0] bias_add_56;
assign bias_add_56 = conv_mac_56 + 4'd7;
logic [31:0] bias_add_57;
assign bias_add_57 = conv_mac_57 + 4'd6;
logic [31:0] bias_add_58;
assign bias_add_58 = conv_mac_58 + 5'd9;
logic [31:0] bias_add_59;
assign bias_add_59 = conv_mac_59 + 6'd16;
logic [31:0] bias_add_60;
assign bias_add_60 = conv_mac_60 - 3'd2;
logic [31:0] bias_add_61;
assign bias_add_61 = conv_mac_61 + 2'd1;
logic [31:0] bias_add_62;
assign bias_add_62 = conv_mac_62 + 6'd17;
logic [31:0] bias_add_63;
assign bias_add_63 = conv_mac_63 - 4'd7;

logic [7:0] relu_0;
assign relu_0[7:0] = (bias_add_0[31]==0) ? ((bias_add_0<3'd6) ? {{bias_add_0[31],bias_add_0[10:4]}} :'d6) : '0;
logic [7:0] relu_1;
assign relu_1[7:0] = (bias_add_1[31]==0) ? ((bias_add_1<3'd6) ? {{bias_add_1[31],bias_add_1[10:4]}} :'d6) : '0;
logic [7:0] relu_2;
assign relu_2[7:0] = (bias_add_2[31]==0) ? ((bias_add_2<3'd6) ? {{bias_add_2[31],bias_add_2[10:4]}} :'d6) : '0;
logic [7:0] relu_3;
assign relu_3[7:0] = (bias_add_3[31]==0) ? ((bias_add_3<3'd6) ? {{bias_add_3[31],bias_add_3[10:4]}} :'d6) : '0;
logic [7:0] relu_4;
assign relu_4[7:0] = (bias_add_4[31]==0) ? ((bias_add_4<3'd6) ? {{bias_add_4[31],bias_add_4[10:4]}} :'d6) : '0;
logic [7:0] relu_5;
assign relu_5[7:0] = (bias_add_5[31]==0) ? ((bias_add_5<3'd6) ? {{bias_add_5[31],bias_add_5[10:4]}} :'d6) : '0;
logic [7:0] relu_6;
assign relu_6[7:0] = (bias_add_6[31]==0) ? ((bias_add_6<3'd6) ? {{bias_add_6[31],bias_add_6[10:4]}} :'d6) : '0;
logic [7:0] relu_7;
assign relu_7[7:0] = (bias_add_7[31]==0) ? ((bias_add_7<3'd6) ? {{bias_add_7[31],bias_add_7[10:4]}} :'d6) : '0;
logic [7:0] relu_8;
assign relu_8[7:0] = (bias_add_8[31]==0) ? ((bias_add_8<3'd6) ? {{bias_add_8[31],bias_add_8[10:4]}} :'d6) : '0;
logic [7:0] relu_9;
assign relu_9[7:0] = (bias_add_9[31]==0) ? ((bias_add_9<3'd6) ? {{bias_add_9[31],bias_add_9[10:4]}} :'d6) : '0;
logic [7:0] relu_10;
assign relu_10[7:0] = (bias_add_10[31]==0) ? ((bias_add_10<3'd6) ? {{bias_add_10[31],bias_add_10[10:4]}} :'d6) : '0;
logic [7:0] relu_11;
assign relu_11[7:0] = (bias_add_11[31]==0) ? ((bias_add_11<3'd6) ? {{bias_add_11[31],bias_add_11[10:4]}} :'d6) : '0;
logic [7:0] relu_12;
assign relu_12[7:0] = (bias_add_12[31]==0) ? ((bias_add_12<3'd6) ? {{bias_add_12[31],bias_add_12[10:4]}} :'d6) : '0;
logic [7:0] relu_13;
assign relu_13[7:0] = (bias_add_13[31]==0) ? ((bias_add_13<3'd6) ? {{bias_add_13[31],bias_add_13[10:4]}} :'d6) : '0;
logic [7:0] relu_14;
assign relu_14[7:0] = (bias_add_14[31]==0) ? ((bias_add_14<3'd6) ? {{bias_add_14[31],bias_add_14[10:4]}} :'d6) : '0;
logic [7:0] relu_15;
assign relu_15[7:0] = (bias_add_15[31]==0) ? ((bias_add_15<3'd6) ? {{bias_add_15[31],bias_add_15[10:4]}} :'d6) : '0;
logic [7:0] relu_16;
assign relu_16[7:0] = (bias_add_16[31]==0) ? ((bias_add_16<3'd6) ? {{bias_add_16[31],bias_add_16[10:4]}} :'d6) : '0;
logic [7:0] relu_17;
assign relu_17[7:0] = (bias_add_17[31]==0) ? ((bias_add_17<3'd6) ? {{bias_add_17[31],bias_add_17[10:4]}} :'d6) : '0;
logic [7:0] relu_18;
assign relu_18[7:0] = (bias_add_18[31]==0) ? ((bias_add_18<3'd6) ? {{bias_add_18[31],bias_add_18[10:4]}} :'d6) : '0;
logic [7:0] relu_19;
assign relu_19[7:0] = (bias_add_19[31]==0) ? ((bias_add_19<3'd6) ? {{bias_add_19[31],bias_add_19[10:4]}} :'d6) : '0;
logic [7:0] relu_20;
assign relu_20[7:0] = (bias_add_20[31]==0) ? ((bias_add_20<3'd6) ? {{bias_add_20[31],bias_add_20[10:4]}} :'d6) : '0;
logic [7:0] relu_21;
assign relu_21[7:0] = (bias_add_21[31]==0) ? ((bias_add_21<3'd6) ? {{bias_add_21[31],bias_add_21[10:4]}} :'d6) : '0;
logic [7:0] relu_22;
assign relu_22[7:0] = (bias_add_22[31]==0) ? ((bias_add_22<3'd6) ? {{bias_add_22[31],bias_add_22[10:4]}} :'d6) : '0;
logic [7:0] relu_23;
assign relu_23[7:0] = (bias_add_23[31]==0) ? ((bias_add_23<3'd6) ? {{bias_add_23[31],bias_add_23[10:4]}} :'d6) : '0;
logic [7:0] relu_24;
assign relu_24[7:0] = (bias_add_24[31]==0) ? ((bias_add_24<3'd6) ? {{bias_add_24[31],bias_add_24[10:4]}} :'d6) : '0;
logic [7:0] relu_25;
assign relu_25[7:0] = (bias_add_25[31]==0) ? ((bias_add_25<3'd6) ? {{bias_add_25[31],bias_add_25[10:4]}} :'d6) : '0;
logic [7:0] relu_26;
assign relu_26[7:0] = (bias_add_26[31]==0) ? ((bias_add_26<3'd6) ? {{bias_add_26[31],bias_add_26[10:4]}} :'d6) : '0;
logic [7:0] relu_27;
assign relu_27[7:0] = (bias_add_27[31]==0) ? ((bias_add_27<3'd6) ? {{bias_add_27[31],bias_add_27[10:4]}} :'d6) : '0;
logic [7:0] relu_28;
assign relu_28[7:0] = (bias_add_28[31]==0) ? ((bias_add_28<3'd6) ? {{bias_add_28[31],bias_add_28[10:4]}} :'d6) : '0;
logic [7:0] relu_29;
assign relu_29[7:0] = (bias_add_29[31]==0) ? ((bias_add_29<3'd6) ? {{bias_add_29[31],bias_add_29[10:4]}} :'d6) : '0;
logic [7:0] relu_30;
assign relu_30[7:0] = (bias_add_30[31]==0) ? ((bias_add_30<3'd6) ? {{bias_add_30[31],bias_add_30[10:4]}} :'d6) : '0;
logic [7:0] relu_31;
assign relu_31[7:0] = (bias_add_31[31]==0) ? ((bias_add_31<3'd6) ? {{bias_add_31[31],bias_add_31[10:4]}} :'d6) : '0;
logic [7:0] relu_32;
assign relu_32[7:0] = (bias_add_32[31]==0) ? ((bias_add_32<3'd6) ? {{bias_add_32[31],bias_add_32[10:4]}} :'d6) : '0;
logic [7:0] relu_33;
assign relu_33[7:0] = (bias_add_33[31]==0) ? ((bias_add_33<3'd6) ? {{bias_add_33[31],bias_add_33[10:4]}} :'d6) : '0;
logic [7:0] relu_34;
assign relu_34[7:0] = (bias_add_34[31]==0) ? ((bias_add_34<3'd6) ? {{bias_add_34[31],bias_add_34[10:4]}} :'d6) : '0;
logic [7:0] relu_35;
assign relu_35[7:0] = (bias_add_35[31]==0) ? ((bias_add_35<3'd6) ? {{bias_add_35[31],bias_add_35[10:4]}} :'d6) : '0;
logic [7:0] relu_36;
assign relu_36[7:0] = (bias_add_36[31]==0) ? ((bias_add_36<3'd6) ? {{bias_add_36[31],bias_add_36[10:4]}} :'d6) : '0;
logic [7:0] relu_37;
assign relu_37[7:0] = (bias_add_37[31]==0) ? ((bias_add_37<3'd6) ? {{bias_add_37[31],bias_add_37[10:4]}} :'d6) : '0;
logic [7:0] relu_38;
assign relu_38[7:0] = (bias_add_38[31]==0) ? ((bias_add_38<3'd6) ? {{bias_add_38[31],bias_add_38[10:4]}} :'d6) : '0;
logic [7:0] relu_39;
assign relu_39[7:0] = (bias_add_39[31]==0) ? ((bias_add_39<3'd6) ? {{bias_add_39[31],bias_add_39[10:4]}} :'d6) : '0;
logic [7:0] relu_40;
assign relu_40[7:0] = (bias_add_40[31]==0) ? ((bias_add_40<3'd6) ? {{bias_add_40[31],bias_add_40[10:4]}} :'d6) : '0;
logic [7:0] relu_41;
assign relu_41[7:0] = (bias_add_41[31]==0) ? ((bias_add_41<3'd6) ? {{bias_add_41[31],bias_add_41[10:4]}} :'d6) : '0;
logic [7:0] relu_42;
assign relu_42[7:0] = (bias_add_42[31]==0) ? ((bias_add_42<3'd6) ? {{bias_add_42[31],bias_add_42[10:4]}} :'d6) : '0;
logic [7:0] relu_43;
assign relu_43[7:0] = (bias_add_43[31]==0) ? ((bias_add_43<3'd6) ? {{bias_add_43[31],bias_add_43[10:4]}} :'d6) : '0;
logic [7:0] relu_44;
assign relu_44[7:0] = (bias_add_44[31]==0) ? ((bias_add_44<3'd6) ? {{bias_add_44[31],bias_add_44[10:4]}} :'d6) : '0;
logic [7:0] relu_45;
assign relu_45[7:0] = (bias_add_45[31]==0) ? ((bias_add_45<3'd6) ? {{bias_add_45[31],bias_add_45[10:4]}} :'d6) : '0;
logic [7:0] relu_46;
assign relu_46[7:0] = (bias_add_46[31]==0) ? ((bias_add_46<3'd6) ? {{bias_add_46[31],bias_add_46[10:4]}} :'d6) : '0;
logic [7:0] relu_47;
assign relu_47[7:0] = (bias_add_47[31]==0) ? ((bias_add_47<3'd6) ? {{bias_add_47[31],bias_add_47[10:4]}} :'d6) : '0;
logic [7:0] relu_48;
assign relu_48[7:0] = (bias_add_48[31]==0) ? ((bias_add_48<3'd6) ? {{bias_add_48[31],bias_add_48[10:4]}} :'d6) : '0;
logic [7:0] relu_49;
assign relu_49[7:0] = (bias_add_49[31]==0) ? ((bias_add_49<3'd6) ? {{bias_add_49[31],bias_add_49[10:4]}} :'d6) : '0;
logic [7:0] relu_50;
assign relu_50[7:0] = (bias_add_50[31]==0) ? ((bias_add_50<3'd6) ? {{bias_add_50[31],bias_add_50[10:4]}} :'d6) : '0;
logic [7:0] relu_51;
assign relu_51[7:0] = (bias_add_51[31]==0) ? ((bias_add_51<3'd6) ? {{bias_add_51[31],bias_add_51[10:4]}} :'d6) : '0;
logic [7:0] relu_52;
assign relu_52[7:0] = (bias_add_52[31]==0) ? ((bias_add_52<3'd6) ? {{bias_add_52[31],bias_add_52[10:4]}} :'d6) : '0;
logic [7:0] relu_53;
assign relu_53[7:0] = (bias_add_53[31]==0) ? ((bias_add_53<3'd6) ? {{bias_add_53[31],bias_add_53[10:4]}} :'d6) : '0;
logic [7:0] relu_54;
assign relu_54[7:0] = (bias_add_54[31]==0) ? ((bias_add_54<3'd6) ? {{bias_add_54[31],bias_add_54[10:4]}} :'d6) : '0;
logic [7:0] relu_55;
assign relu_55[7:0] = (bias_add_55[31]==0) ? ((bias_add_55<3'd6) ? {{bias_add_55[31],bias_add_55[10:4]}} :'d6) : '0;
logic [7:0] relu_56;
assign relu_56[7:0] = (bias_add_56[31]==0) ? ((bias_add_56<3'd6) ? {{bias_add_56[31],bias_add_56[10:4]}} :'d6) : '0;
logic [7:0] relu_57;
assign relu_57[7:0] = (bias_add_57[31]==0) ? ((bias_add_57<3'd6) ? {{bias_add_57[31],bias_add_57[10:4]}} :'d6) : '0;
logic [7:0] relu_58;
assign relu_58[7:0] = (bias_add_58[31]==0) ? ((bias_add_58<3'd6) ? {{bias_add_58[31],bias_add_58[10:4]}} :'d6) : '0;
logic [7:0] relu_59;
assign relu_59[7:0] = (bias_add_59[31]==0) ? ((bias_add_59<3'd6) ? {{bias_add_59[31],bias_add_59[10:4]}} :'d6) : '0;
logic [7:0] relu_60;
assign relu_60[7:0] = (bias_add_60[31]==0) ? ((bias_add_60<3'd6) ? {{bias_add_60[31],bias_add_60[10:4]}} :'d6) : '0;
logic [7:0] relu_61;
assign relu_61[7:0] = (bias_add_61[31]==0) ? ((bias_add_61<3'd6) ? {{bias_add_61[31],bias_add_61[10:4]}} :'d6) : '0;
logic [7:0] relu_62;
assign relu_62[7:0] = (bias_add_62[31]==0) ? ((bias_add_62<3'd6) ? {{bias_add_62[31],bias_add_62[10:4]}} :'d6) : '0;
logic [7:0] relu_63;
assign relu_63[7:0] = (bias_add_63[31]==0) ? ((bias_add_63<3'd6) ? {{bias_add_63[31],bias_add_63[10:4]}} :'d6) : '0;

assign output_act = {
	relu_63,
	relu_62,
	relu_61,
	relu_60,
	relu_59,
	relu_58,
	relu_57,
	relu_56,
	relu_55,
	relu_54,
	relu_53,
	relu_52,
	relu_51,
	relu_50,
	relu_49,
	relu_48,
	relu_47,
	relu_46,
	relu_45,
	relu_44,
	relu_43,
	relu_42,
	relu_41,
	relu_40,
	relu_39,
	relu_38,
	relu_37,
	relu_36,
	relu_35,
	relu_34,
	relu_33,
	relu_32,
	relu_31,
	relu_30,
	relu_29,
	relu_28,
	relu_27,
	relu_26,
	relu_25,
	relu_24,
	relu_23,
	relu_22,
	relu_21,
	relu_20,
	relu_19,
	relu_18,
	relu_17,
	relu_16,
	relu_15,
	relu_14,
	relu_13,
	relu_12,
	relu_11,
	relu_10,
	relu_9,
	relu_8,
	relu_7,
	relu_6,
	relu_5,
	relu_4,
	relu_3,
	relu_2,
	relu_1,
	relu_0
};

endmodule

module line_buffer_array_k7
#(
    parameter KER_SIZE = 7,
    parameter BITWIDTH = 8,
    parameter AW       = 8,
    parameter PAD      = 1
)
(
    input logic clk,
    input logic rstn,
    input logic [BITWIDTH*KER_SIZE-1:0] pixel_in,
    input logic [3-1:0] col_ptr,
    input logic [3-1:0] init_col_ptr,
    input logic [KER_SIZE-1:0] left_pad_mask,
    input logic [KER_SIZE-1:0] right_pad_mask,
    output logic [BITWIDTH*KER_SIZE*KER_SIZE-1:0] pixel_out   
);

// wires
//logic [KER_SIZE*BITWIDTH-1:0] pixel_col [KER_SIZE-1:0];
logic [KER_SIZE*KER_SIZE*BITWIDTH-1:0] pixel_col;

//logic [KER_SIZE*BITWIDTH-1:0] pixel_row [KER_SIZE-1:0];
logic [KER_SIZE*KER_SIZE*BITWIDTH-1:0] pixel_row;

//logic [KER_SIZE*BITWIDTH-1:0] padded_pixel_row [KER_SIZE-1:0];
logic [KER_SIZE*KER_SIZE*BITWIDTH-1:0] padded_pixel_row;

//logic [KER_SIZE*BITWIDTH-1:0] left_padded_pixel_col [KER_SIZE-1:0];
logic [KER_SIZE*KER_SIZE*BITWIDTH-1:0] left_padded_pixel_col;

//logic [KER_SIZE*BITWIDTH-1:0] right_padded_pixel_col [KER_SIZE-1:0];
logic [KER_SIZE*KER_SIZE*BITWIDTH-1:0] right_padded_pixel_col; 

logic [KER_SIZE*KER_SIZE*BITWIDTH-1:0] pixel_out_wire;
logic [KER_SIZE*KER_SIZE*BITWIDTH-1:0] stored_pixel_out;
logic ready;

logic [8-1:0] global_col_ptr;
logic ready_reg;

// reg array
genvar i,j;
generate

for (i = 0; i < KER_SIZE; i++) begin: genblk_14
    d_flop #(
        .BITWIDTH (BITWIDTH*KER_SIZE)
    ) reg_inst (
        .clk (clk),
        .rstn (rstn),
        .valid (col_ptr == i),
        .D (pixel_in),
        .Q (pixel_col[(i+1)*KER_SIZE*BITWIDTH -1:i*KER_SIZE*BITWIDTH])
    ); // each d_flop stores a column of data
//always@(posedge clk) begin 
assign left_padded_pixel_col[(i+1)*KER_SIZE*BITWIDTH -1:i*KER_SIZE*BITWIDTH] = (left_pad_mask[i]==1)? {(KER_SIZE*BITWIDTH){1'b0}} : pixel_col[(i+1)*KER_SIZE*BITWIDTH -1:i*KER_SIZE*BITWIDTH];//left padding
//end 
end
endgenerate

// reshape
always_comb begin
    case (1'b1)
(col_ptr == 'd4): pixel_out_wire = {pixel_in[7*BITWIDTH-1:6*BITWIDTH],left_padded_pixel_col[4*7*BITWIDTH-1:4*6*BITWIDTH],left_padded_pixel_col[3*7*BITWIDTH-1:3*6*BITWIDTH],left_padded_pixel_col[2*7*BITWIDTH-1:2*6*BITWIDTH],left_padded_pixel_col[7*BITWIDTH-1:6*BITWIDTH],left_padded_pixel_col[7*7*BITWIDTH-1:7*6*BITWIDTH],left_padded_pixel_col[6*7*BITWIDTH-1:6*6*BITWIDTH],
                                    pixel_in[6*BITWIDTH-1:5*BITWIDTH],left_padded_pixel_col[4*6*BITWIDTH-1:4*5*BITWIDTH],left_padded_pixel_col[3*6*BITWIDTH-1:3*5*BITWIDTH],left_padded_pixel_col[2*6*BITWIDTH-1:2*5*BITWIDTH],left_padded_pixel_col[6*BITWIDTH-1:5*BITWIDTH],left_padded_pixel_col[7*6*BITWIDTH-1:7*5*BITWIDTH],left_padded_pixel_col[6*6*BITWIDTH-1:6*5*BITWIDTH],
                                    pixel_in[5*BITWIDTH-1:4*BITWIDTH],left_padded_pixel_col[4*5*BITWIDTH-1:4*4*BITWIDTH],left_padded_pixel_col[3*5*BITWIDTH-1:3*4*BITWIDTH],left_padded_pixel_col[2*5*BITWIDTH-1:2*4*BITWIDTH],left_padded_pixel_col[5*BITWIDTH-1:4*BITWIDTH],left_padded_pixel_col[7*5*BITWIDTH-1:7*4*BITWIDTH],left_padded_pixel_col[6*5*BITWIDTH-1:6*4*BITWIDTH],
                                    pixel_in[4*BITWIDTH-1:3*BITWIDTH],left_padded_pixel_col[4*4*BITWIDTH-1:4*3*BITWIDTH],left_padded_pixel_col[3*4*BITWIDTH-1:3*3*BITWIDTH],left_padded_pixel_col[2*4*BITWIDTH-1:2*3*BITWIDTH],left_padded_pixel_col[4*BITWIDTH-1:3*BITWIDTH],left_padded_pixel_col[7*4*BITWIDTH-1:7*3*BITWIDTH],left_padded_pixel_col[6*4*BITWIDTH-1:6*3*BITWIDTH],
                                    pixel_in[3*BITWIDTH-1:2*BITWIDTH],left_padded_pixel_col[4*3*BITWIDTH-1:4*2*BITWIDTH],left_padded_pixel_col[3*3*BITWIDTH-1:3*2*BITWIDTH],left_padded_pixel_col[2*3*BITWIDTH-1:2*2*BITWIDTH],left_padded_pixel_col[3*BITWIDTH-1:2*BITWIDTH],left_padded_pixel_col[7*3*BITWIDTH-1:7*2*BITWIDTH],left_padded_pixel_col[6*3*BITWIDTH-1:6*2*BITWIDTH],
                                    pixel_in[2*BITWIDTH-1:1*BITWIDTH],left_padded_pixel_col[4*2*BITWIDTH-1:4*1*BITWIDTH],left_padded_pixel_col[3*2*BITWIDTH-1:3*1*BITWIDTH],left_padded_pixel_col[2*2*BITWIDTH-1:2*1*BITWIDTH],left_padded_pixel_col[2*BITWIDTH-1:1*BITWIDTH],left_padded_pixel_col[7*2*BITWIDTH-1:7*1*BITWIDTH],left_padded_pixel_col[6*2*BITWIDTH-1:6*1*BITWIDTH],
                                    pixel_in[1*BITWIDTH-1:0*BITWIDTH],left_padded_pixel_col[4*1*BITWIDTH-1:4*0*BITWIDTH],left_padded_pixel_col[3*1*BITWIDTH-1:3*0*BITWIDTH],left_padded_pixel_col[2*1*BITWIDTH-1:2*0*BITWIDTH],left_padded_pixel_col[1*BITWIDTH-1:0*BITWIDTH],left_padded_pixel_col[7*1*BITWIDTH-1:7*0*BITWIDTH],left_padded_pixel_col[6*1*BITWIDTH-1:6*0*BITWIDTH]};
                                    
(col_ptr == 'd3): pixel_out_wire = {pixel_in[7*BITWIDTH-1:6*BITWIDTH],left_padded_pixel_col[3*7*BITWIDTH-1:3*6*BITWIDTH],left_padded_pixel_col[2*7*BITWIDTH-1:2*6*BITWIDTH],left_padded_pixel_col[7*BITWIDTH-1:6*BITWIDTH],left_padded_pixel_col[7*7*BITWIDTH-1:7*6*BITWIDTH],left_padded_pixel_col[6*7*BITWIDTH-1:6*6*BITWIDTH],left_padded_pixel_col[5*7*BITWIDTH-1:5*6*BITWIDTH],
                                    pixel_in[6*BITWIDTH-1:5*BITWIDTH],left_padded_pixel_col[3*6*BITWIDTH-1:3*5*BITWIDTH],left_padded_pixel_col[2*6*BITWIDTH-1:2*5*BITWIDTH],left_padded_pixel_col[6*BITWIDTH-1:5*BITWIDTH],left_padded_pixel_col[7*6*BITWIDTH-1:7*5*BITWIDTH],left_padded_pixel_col[6*6*BITWIDTH-1:6*5*BITWIDTH],left_padded_pixel_col[5*6*BITWIDTH-1:5*5*BITWIDTH],
                                    pixel_in[5*BITWIDTH-1:4*BITWIDTH],left_padded_pixel_col[3*5*BITWIDTH-1:3*4*BITWIDTH],left_padded_pixel_col[2*5*BITWIDTH-1:2*4*BITWIDTH],left_padded_pixel_col[5*BITWIDTH-1:4*BITWIDTH],left_padded_pixel_col[7*5*BITWIDTH-1:7*4*BITWIDTH],left_padded_pixel_col[6*5*BITWIDTH-1:6*4*BITWIDTH],left_padded_pixel_col[5*5*BITWIDTH-1:5*4*BITWIDTH],
                                    pixel_in[4*BITWIDTH-1:3*BITWIDTH],left_padded_pixel_col[3*4*BITWIDTH-1:3*3*BITWIDTH],left_padded_pixel_col[2*4*BITWIDTH-1:2*3*BITWIDTH],left_padded_pixel_col[4*BITWIDTH-1:3*BITWIDTH],left_padded_pixel_col[7*4*BITWIDTH-1:7*3*BITWIDTH],left_padded_pixel_col[6*4*BITWIDTH-1:6*3*BITWIDTH],left_padded_pixel_col[5*4*BITWIDTH-1:5*3*BITWIDTH],
                                    pixel_in[3*BITWIDTH-1:2*BITWIDTH],left_padded_pixel_col[3*3*BITWIDTH-1:3*2*BITWIDTH],left_padded_pixel_col[2*3*BITWIDTH-1:2*2*BITWIDTH],left_padded_pixel_col[3*BITWIDTH-1:2*BITWIDTH],left_padded_pixel_col[7*3*BITWIDTH-1:7*2*BITWIDTH],left_padded_pixel_col[6*3*BITWIDTH-1:6*2*BITWIDTH],left_padded_pixel_col[5*3*BITWIDTH-1:5*2*BITWIDTH],
                                    pixel_in[2*BITWIDTH-1:1*BITWIDTH],left_padded_pixel_col[3*2*BITWIDTH-1:3*1*BITWIDTH],left_padded_pixel_col[2*2*BITWIDTH-1:2*1*BITWIDTH],left_padded_pixel_col[2*BITWIDTH-1:1*BITWIDTH],left_padded_pixel_col[7*2*BITWIDTH-1:7*1*BITWIDTH],left_padded_pixel_col[6*2*BITWIDTH-1:6*1*BITWIDTH],left_padded_pixel_col[5*2*BITWIDTH-1:5*1*BITWIDTH],
                                    pixel_in[1*BITWIDTH-1:0*BITWIDTH],left_padded_pixel_col[3*1*BITWIDTH-1:3*0*BITWIDTH],left_padded_pixel_col[2*1*BITWIDTH-1:2*0*BITWIDTH],left_padded_pixel_col[1*BITWIDTH-1:0*BITWIDTH],left_padded_pixel_col[7*1*BITWIDTH-1:7*0*BITWIDTH],left_padded_pixel_col[6*1*BITWIDTH-1:6*0*BITWIDTH],left_padded_pixel_col[5*1*BITWIDTH-1:5*0*BITWIDTH]};
                                    
(col_ptr == 'd2): pixel_out_wire = {pixel_in[7*BITWIDTH-1:6*BITWIDTH],left_padded_pixel_col[2*7*BITWIDTH-1:2*6*BITWIDTH],left_padded_pixel_col[7*BITWIDTH-1:6*BITWIDTH],left_padded_pixel_col[7*7*BITWIDTH-1:7*6*BITWIDTH],left_padded_pixel_col[6*7*BITWIDTH-1:6*6*BITWIDTH],left_padded_pixel_col[5*7*BITWIDTH-1:5*6*BITWIDTH],left_padded_pixel_col[4*7*BITWIDTH-1:4*6*BITWIDTH],
                                    pixel_in[6*BITWIDTH-1:5*BITWIDTH],left_padded_pixel_col[2*6*BITWIDTH-1:2*5*BITWIDTH],left_padded_pixel_col[6*BITWIDTH-1:5*BITWIDTH],left_padded_pixel_col[7*6*BITWIDTH-1:7*5*BITWIDTH],left_padded_pixel_col[6*6*BITWIDTH-1:6*5*BITWIDTH],left_padded_pixel_col[5*6*BITWIDTH-1:5*5*BITWIDTH],left_padded_pixel_col[4*6*BITWIDTH-1:4*5*BITWIDTH],
                                    pixel_in[5*BITWIDTH-1:4*BITWIDTH],left_padded_pixel_col[2*5*BITWIDTH-1:2*4*BITWIDTH],left_padded_pixel_col[5*BITWIDTH-1:4*BITWIDTH],left_padded_pixel_col[7*5*BITWIDTH-1:7*4*BITWIDTH],left_padded_pixel_col[6*5*BITWIDTH-1:6*4*BITWIDTH],left_padded_pixel_col[5*5*BITWIDTH-1:5*4*BITWIDTH],left_padded_pixel_col[4*5*BITWIDTH-1:4*4*BITWIDTH],
                                    pixel_in[4*BITWIDTH-1:3*BITWIDTH],left_padded_pixel_col[2*4*BITWIDTH-1:2*3*BITWIDTH],left_padded_pixel_col[4*BITWIDTH-1:3*BITWIDTH],left_padded_pixel_col[7*4*BITWIDTH-1:7*3*BITWIDTH],left_padded_pixel_col[6*4*BITWIDTH-1:6*3*BITWIDTH],left_padded_pixel_col[5*4*BITWIDTH-1:5*3*BITWIDTH],left_padded_pixel_col[4*4*BITWIDTH-1:4*3*BITWIDTH],
                                    pixel_in[3*BITWIDTH-1:2*BITWIDTH],left_padded_pixel_col[2*3*BITWIDTH-1:2*2*BITWIDTH],left_padded_pixel_col[3*BITWIDTH-1:2*BITWIDTH],left_padded_pixel_col[7*3*BITWIDTH-1:7*2*BITWIDTH],left_padded_pixel_col[6*3*BITWIDTH-1:6*2*BITWIDTH],left_padded_pixel_col[5*3*BITWIDTH-1:5*2*BITWIDTH],left_padded_pixel_col[4*3*BITWIDTH-1:4*2*BITWIDTH],
                                    pixel_in[2*BITWIDTH-1:1*BITWIDTH],left_padded_pixel_col[2*2*BITWIDTH-1:2*1*BITWIDTH],left_padded_pixel_col[2*BITWIDTH-1:1*BITWIDTH],left_padded_pixel_col[7*2*BITWIDTH-1:7*1*BITWIDTH],left_padded_pixel_col[6*2*BITWIDTH-1:6*1*BITWIDTH],left_padded_pixel_col[5*2*BITWIDTH-1:5*1*BITWIDTH],left_padded_pixel_col[4*2*BITWIDTH-1:4*1*BITWIDTH],
                                    pixel_in[1*BITWIDTH-1:0*BITWIDTH],left_padded_pixel_col[2*1*BITWIDTH-1:2*0*BITWIDTH],left_padded_pixel_col[1*BITWIDTH-1:0*BITWIDTH],left_padded_pixel_col[7*1*BITWIDTH-1:7*0*BITWIDTH],left_padded_pixel_col[6*1*BITWIDTH-1:6*0*BITWIDTH],left_padded_pixel_col[5*1*BITWIDTH-1:5*0*BITWIDTH],left_padded_pixel_col[4*1*BITWIDTH-1:4*0*BITWIDTH]};   
                                    
(col_ptr == 'd1): pixel_out_wire = {pixel_in[7*BITWIDTH-1:6*BITWIDTH],left_padded_pixel_col[7*BITWIDTH-1:6*BITWIDTH],left_padded_pixel_col[7*7*BITWIDTH-1:7*6*BITWIDTH],left_padded_pixel_col[6*7*BITWIDTH-1:6*6*BITWIDTH],left_padded_pixel_col[5*7*BITWIDTH-1:5*6*BITWIDTH],left_padded_pixel_col[4*7*BITWIDTH-1:4*6*BITWIDTH],left_padded_pixel_col[3*7*BITWIDTH-1:3*6*BITWIDTH],
                                    pixel_in[6*BITWIDTH-1:5*BITWIDTH],left_padded_pixel_col[6*BITWIDTH-1:5*BITWIDTH],left_padded_pixel_col[7*6*BITWIDTH-1:7*5*BITWIDTH],left_padded_pixel_col[6*6*BITWIDTH-1:6*5*BITWIDTH],left_padded_pixel_col[5*6*BITWIDTH-1:5*5*BITWIDTH],left_padded_pixel_col[4*6*BITWIDTH-1:4*5*BITWIDTH],left_padded_pixel_col[3*6*BITWIDTH-1:3*5*BITWIDTH],
                                    pixel_in[5*BITWIDTH-1:4*BITWIDTH],left_padded_pixel_col[5*BITWIDTH-1:4*BITWIDTH],left_padded_pixel_col[7*5*BITWIDTH-1:7*4*BITWIDTH],left_padded_pixel_col[6*5*BITWIDTH-1:6*4*BITWIDTH],left_padded_pixel_col[5*5*BITWIDTH-1:5*4*BITWIDTH],left_padded_pixel_col[4*5*BITWIDTH-1:4*4*BITWIDTH],left_padded_pixel_col[3*5*BITWIDTH-1:3*4*BITWIDTH],
                                    pixel_in[4*BITWIDTH-1:3*BITWIDTH],left_padded_pixel_col[4*BITWIDTH-1:3*BITWIDTH],left_padded_pixel_col[7*4*BITWIDTH-1:7*3*BITWIDTH],left_padded_pixel_col[6*4*BITWIDTH-1:6*3*BITWIDTH],left_padded_pixel_col[5*4*BITWIDTH-1:5*3*BITWIDTH],left_padded_pixel_col[4*4*BITWIDTH-1:4*3*BITWIDTH],left_padded_pixel_col[3*4*BITWIDTH-1:3*3*BITWIDTH],
                                    pixel_in[3*BITWIDTH-1:2*BITWIDTH],left_padded_pixel_col[3*BITWIDTH-1:2*BITWIDTH],left_padded_pixel_col[7*3*BITWIDTH-1:7*2*BITWIDTH],left_padded_pixel_col[6*3*BITWIDTH-1:6*2*BITWIDTH],left_padded_pixel_col[5*3*BITWIDTH-1:5*2*BITWIDTH],left_padded_pixel_col[4*3*BITWIDTH-1:4*2*BITWIDTH],left_padded_pixel_col[3*3*BITWIDTH-1:3*2*BITWIDTH],
                                    pixel_in[2*BITWIDTH-1:1*BITWIDTH],left_padded_pixel_col[2*BITWIDTH-1:1*BITWIDTH],left_padded_pixel_col[7*2*BITWIDTH-1:7*1*BITWIDTH],left_padded_pixel_col[6*2*BITWIDTH-1:6*1*BITWIDTH],left_padded_pixel_col[5*2*BITWIDTH-1:5*1*BITWIDTH],left_padded_pixel_col[4*2*BITWIDTH-1:4*1*BITWIDTH],left_padded_pixel_col[3*2*BITWIDTH-1:3*1*BITWIDTH],
                                    pixel_in[1*BITWIDTH-1:0*BITWIDTH],left_padded_pixel_col[1*BITWIDTH-1:0*BITWIDTH],left_padded_pixel_col[7*1*BITWIDTH-1:7*0*BITWIDTH],left_padded_pixel_col[6*1*BITWIDTH-1:6*0*BITWIDTH],left_padded_pixel_col[5*1*BITWIDTH-1:5*0*BITWIDTH],left_padded_pixel_col[4*1*BITWIDTH-1:4*0*BITWIDTH],left_padded_pixel_col[3*1*BITWIDTH-1:3*0*BITWIDTH]}; 
                                    
(col_ptr == 'd0): pixel_out_wire = {pixel_in[7*BITWIDTH-1:6*BITWIDTH],left_padded_pixel_col[7*7*BITWIDTH-1:7*6*BITWIDTH],left_padded_pixel_col[6*7*BITWIDTH-1:6*6*BITWIDTH],left_padded_pixel_col[5*7*BITWIDTH-1:5*6*BITWIDTH],left_padded_pixel_col[4*7*BITWIDTH-1:4*6*BITWIDTH],left_padded_pixel_col[3*7*BITWIDTH-1:3*6*BITWIDTH],left_padded_pixel_col[2*7*BITWIDTH-1:2*6*BITWIDTH],
                                    pixel_in[6*BITWIDTH-1:5*BITWIDTH],left_padded_pixel_col[7*6*BITWIDTH-1:7*5*BITWIDTH],left_padded_pixel_col[6*6*BITWIDTH-1:6*5*BITWIDTH],left_padded_pixel_col[5*6*BITWIDTH-1:5*5*BITWIDTH],left_padded_pixel_col[4*6*BITWIDTH-1:4*5*BITWIDTH],left_padded_pixel_col[3*6*BITWIDTH-1:3*5*BITWIDTH],left_padded_pixel_col[2*6*BITWIDTH-1:2*5*BITWIDTH],
                                    pixel_in[5*BITWIDTH-1:4*BITWIDTH],left_padded_pixel_col[7*5*BITWIDTH-1:7*4*BITWIDTH],left_padded_pixel_col[6*5*BITWIDTH-1:6*4*BITWIDTH],left_padded_pixel_col[5*5*BITWIDTH-1:5*4*BITWIDTH],left_padded_pixel_col[4*5*BITWIDTH-1:4*4*BITWIDTH],left_padded_pixel_col[3*5*BITWIDTH-1:3*4*BITWIDTH],left_padded_pixel_col[2*5*BITWIDTH-1:2*4*BITWIDTH],
                                    pixel_in[4*BITWIDTH-1:3*BITWIDTH],left_padded_pixel_col[7*4*BITWIDTH-1:7*3*BITWIDTH],left_padded_pixel_col[6*4*BITWIDTH-1:6*3*BITWIDTH],left_padded_pixel_col[5*4*BITWIDTH-1:5*3*BITWIDTH],left_padded_pixel_col[4*4*BITWIDTH-1:4*3*BITWIDTH],left_padded_pixel_col[3*4*BITWIDTH-1:3*3*BITWIDTH],left_padded_pixel_col[2*4*BITWIDTH-1:2*3*BITWIDTH],
                                    pixel_in[3*BITWIDTH-1:2*BITWIDTH],left_padded_pixel_col[7*3*BITWIDTH-1:7*2*BITWIDTH],left_padded_pixel_col[6*3*BITWIDTH-1:6*2*BITWIDTH],left_padded_pixel_col[5*3*BITWIDTH-1:5*2*BITWIDTH],left_padded_pixel_col[4*3*BITWIDTH-1:4*2*BITWIDTH],left_padded_pixel_col[3*3*BITWIDTH-1:3*2*BITWIDTH],left_padded_pixel_col[2*3*BITWIDTH-1:2*2*BITWIDTH],
                                    pixel_in[2*BITWIDTH-1:1*BITWIDTH],left_padded_pixel_col[7*2*BITWIDTH-1:7*1*BITWIDTH],left_padded_pixel_col[6*2*BITWIDTH-1:6*1*BITWIDTH],left_padded_pixel_col[5*2*BITWIDTH-1:5*1*BITWIDTH],left_padded_pixel_col[4*2*BITWIDTH-1:4*1*BITWIDTH],left_padded_pixel_col[3*2*BITWIDTH-1:3*1*BITWIDTH],left_padded_pixel_col[2*2*BITWIDTH-1:2*1*BITWIDTH],
                                    pixel_in[1*BITWIDTH-1:0*BITWIDTH],left_padded_pixel_col[7*1*BITWIDTH-1:7*0*BITWIDTH],left_padded_pixel_col[6*1*BITWIDTH-1:6*0*BITWIDTH],left_padded_pixel_col[5*1*BITWIDTH-1:5*0*BITWIDTH],left_padded_pixel_col[4*1*BITWIDTH-1:4*0*BITWIDTH],left_padded_pixel_col[3*1*BITWIDTH-1:3*0*BITWIDTH],left_padded_pixel_col[2*1*BITWIDTH-1:2*0*BITWIDTH]};

(col_ptr == 'd5): pixel_out_wire = {pixel_in[7*BITWIDTH-1:6*BITWIDTH],left_padded_pixel_col[5*7*BITWIDTH-1:5*6*BITWIDTH],left_padded_pixel_col[4*7*BITWIDTH-1:4*6*BITWIDTH],left_padded_pixel_col[3*7*BITWIDTH-1:3*6*BITWIDTH],left_padded_pixel_col[2*7*BITWIDTH-1:2*6*BITWIDTH],left_padded_pixel_col[7*BITWIDTH-1:6*BITWIDTH],left_padded_pixel_col[7*7*BITWIDTH-1:7*6*BITWIDTH],
                                    pixel_in[6*BITWIDTH-1:5*BITWIDTH],left_padded_pixel_col[5*6*BITWIDTH-1:5*5*BITWIDTH],left_padded_pixel_col[4*6*BITWIDTH-1:4*5*BITWIDTH],left_padded_pixel_col[3*6*BITWIDTH-1:3*5*BITWIDTH],left_padded_pixel_col[2*6*BITWIDTH-1:2*5*BITWIDTH],left_padded_pixel_col[6*BITWIDTH-1:5*BITWIDTH],left_padded_pixel_col[7*6*BITWIDTH-1:7*5*BITWIDTH],
                                    pixel_in[5*BITWIDTH-1:4*BITWIDTH],left_padded_pixel_col[5*5*BITWIDTH-1:5*4*BITWIDTH],left_padded_pixel_col[4*5*BITWIDTH-1:4*4*BITWIDTH],left_padded_pixel_col[3*5*BITWIDTH-1:3*4*BITWIDTH],left_padded_pixel_col[2*5*BITWIDTH-1:2*4*BITWIDTH],left_padded_pixel_col[5*BITWIDTH-1:4*BITWIDTH],left_padded_pixel_col[7*5*BITWIDTH-1:7*4*BITWIDTH],
                                    pixel_in[4*BITWIDTH-1:3*BITWIDTH],left_padded_pixel_col[5*4*BITWIDTH-1:5*3*BITWIDTH],left_padded_pixel_col[4*4*BITWIDTH-1:4*3*BITWIDTH],left_padded_pixel_col[3*4*BITWIDTH-1:3*3*BITWIDTH],left_padded_pixel_col[2*4*BITWIDTH-1:2*3*BITWIDTH],left_padded_pixel_col[4*BITWIDTH-1:3*BITWIDTH],left_padded_pixel_col[7*4*BITWIDTH-1:7*3*BITWIDTH],
                                    pixel_in[3*BITWIDTH-1:2*BITWIDTH],left_padded_pixel_col[5*3*BITWIDTH-1:5*2*BITWIDTH],left_padded_pixel_col[4*3*BITWIDTH-1:4*2*BITWIDTH],left_padded_pixel_col[3*3*BITWIDTH-1:3*2*BITWIDTH],left_padded_pixel_col[2*3*BITWIDTH-1:2*2*BITWIDTH],left_padded_pixel_col[3*BITWIDTH-1:2*BITWIDTH],left_padded_pixel_col[7*3*BITWIDTH-1:7*2*BITWIDTH],
                                    pixel_in[2*BITWIDTH-1:1*BITWIDTH],left_padded_pixel_col[5*2*BITWIDTH-1:5*1*BITWIDTH],left_padded_pixel_col[4*2*BITWIDTH-1:4*1*BITWIDTH],left_padded_pixel_col[3*2*BITWIDTH-1:3*1*BITWIDTH],left_padded_pixel_col[2*2*BITWIDTH-1:2*1*BITWIDTH],left_padded_pixel_col[2*BITWIDTH-1:1*BITWIDTH],left_padded_pixel_col[7*2*BITWIDTH-1:7*1*BITWIDTH],
                                    pixel_in[1*BITWIDTH-1:0*BITWIDTH],left_padded_pixel_col[5*1*BITWIDTH-1:5*0*BITWIDTH],left_padded_pixel_col[4*1*BITWIDTH-1:4*0*BITWIDTH],left_padded_pixel_col[3*1*BITWIDTH-1:3*0*BITWIDTH],left_padded_pixel_col[2*1*BITWIDTH-1:2*0*BITWIDTH],left_padded_pixel_col[1*BITWIDTH-1:0*BITWIDTH],left_padded_pixel_col[7*1*BITWIDTH-1:7*0*BITWIDTH]};

(col_ptr == 'd6): pixel_out_wire = {pixel_in[7*BITWIDTH-1:6*BITWIDTH],left_padded_pixel_col[6*7*BITWIDTH-1:6*6*BITWIDTH],left_padded_pixel_col[5*7*BITWIDTH-1:5*6*BITWIDTH],left_padded_pixel_col[4*7*BITWIDTH-1:4*6*BITWIDTH],left_padded_pixel_col[3*7*BITWIDTH-1:3*6*BITWIDTH],left_padded_pixel_col[2*7*BITWIDTH-1:2*6*BITWIDTH],left_padded_pixel_col[7*BITWIDTH-1:6*BITWIDTH],
                                    pixel_in[6*BITWIDTH-1:5*BITWIDTH],left_padded_pixel_col[6*6*BITWIDTH-1:6*5*BITWIDTH],left_padded_pixel_col[5*6*BITWIDTH-1:5*5*BITWIDTH],left_padded_pixel_col[4*6*BITWIDTH-1:4*5*BITWIDTH],left_padded_pixel_col[3*6*BITWIDTH-1:3*5*BITWIDTH],left_padded_pixel_col[2*6*BITWIDTH-1:2*5*BITWIDTH],left_padded_pixel_col[6*BITWIDTH-1:5*BITWIDTH],
                                    pixel_in[5*BITWIDTH-1:4*BITWIDTH],left_padded_pixel_col[6*5*BITWIDTH-1:6*4*BITWIDTH],left_padded_pixel_col[5*5*BITWIDTH-1:5*4*BITWIDTH],left_padded_pixel_col[4*5*BITWIDTH-1:4*4*BITWIDTH],left_padded_pixel_col[3*5*BITWIDTH-1:3*4*BITWIDTH],left_padded_pixel_col[2*5*BITWIDTH-1:2*4*BITWIDTH],left_padded_pixel_col[5*BITWIDTH-1:4*BITWIDTH],
                                    pixel_in[4*BITWIDTH-1:3*BITWIDTH],left_padded_pixel_col[6*4*BITWIDTH-1:6*3*BITWIDTH],left_padded_pixel_col[5*4*BITWIDTH-1:5*3*BITWIDTH],left_padded_pixel_col[4*4*BITWIDTH-1:4*3*BITWIDTH],left_padded_pixel_col[3*4*BITWIDTH-1:3*3*BITWIDTH],left_padded_pixel_col[2*4*BITWIDTH-1:2*3*BITWIDTH],left_padded_pixel_col[4*BITWIDTH-1:3*BITWIDTH],
                                    pixel_in[3*BITWIDTH-1:2*BITWIDTH],left_padded_pixel_col[6*3*BITWIDTH-1:6*2*BITWIDTH],left_padded_pixel_col[5*3*BITWIDTH-1:5*2*BITWIDTH],left_padded_pixel_col[4*3*BITWIDTH-1:4*2*BITWIDTH],left_padded_pixel_col[3*3*BITWIDTH-1:3*2*BITWIDTH],left_padded_pixel_col[2*3*BITWIDTH-1:2*2*BITWIDTH],left_padded_pixel_col[3*BITWIDTH-1:2*BITWIDTH],
                                    pixel_in[2*BITWIDTH-1:1*BITWIDTH],left_padded_pixel_col[6*2*BITWIDTH-1:6*1*BITWIDTH],left_padded_pixel_col[5*2*BITWIDTH-1:5*1*BITWIDTH],left_padded_pixel_col[4*2*BITWIDTH-1:4*1*BITWIDTH],left_padded_pixel_col[3*2*BITWIDTH-1:3*1*BITWIDTH],left_padded_pixel_col[2*2*BITWIDTH-1:2*1*BITWIDTH],left_padded_pixel_col[2*BITWIDTH-1:1*BITWIDTH],
                                    pixel_in[1*BITWIDTH-1:0*BITWIDTH],left_padded_pixel_col[6*1*BITWIDTH-1:6*0*BITWIDTH],left_padded_pixel_col[5*1*BITWIDTH-1:5*0*BITWIDTH],left_padded_pixel_col[4*1*BITWIDTH-1:4*0*BITWIDTH],left_padded_pixel_col[3*1*BITWIDTH-1:3*0*BITWIDTH],left_padded_pixel_col[2*1*BITWIDTH-1:2*0*BITWIDTH],left_padded_pixel_col[1*BITWIDTH-1:0*BITWIDTH]};
        default:          pixel_out_wire = '0;
    endcase
end



// output flop
always_ff @(posedge clk) begin
    if (!rstn) begin
        stored_pixel_out <= '0;
    end
    else if (ready) begin
        stored_pixel_out <= pixel_out_wire;
    end
    else begin
        stored_pixel_out <= stored_pixel_out;
    end
end

generate
	for (i = 0; i < KER_SIZE ; i++) begin: genblk_20
		assign pixel_row[(i+1)*KER_SIZE*BITWIDTH-1:i*KER_SIZE*BITWIDTH] = stored_pixel_out[KER_SIZE*BITWIDTH*i+:KER_SIZE*BITWIDTH];
		assign pixel_out[KER_SIZE*BITWIDTH*i+:KER_SIZE*BITWIDTH] = padded_pixel_row[(i+1)*KER_SIZE*BITWIDTH-1:i*KER_SIZE*BITWIDTH];
	end
endgenerate

generate
	for (i = 0; i < KER_SIZE ; i++) begin: genblk_15
	for (j = 0; j < KER_SIZE ; j++) begin: genblk_16
		assign padded_pixel_row[(i*KER_SIZE*BITWIDTH + BITWIDTH*j)+:BITWIDTH] = right_pad_mask[j] ?{BITWIDTH{1'b0}}:pixel_row[(i*KER_SIZE*BITWIDTH + BITWIDTH*j)+:BITWIDTH];
	end
	end

endgenerate


assign ready =  init_col_ptr == KER_SIZE-1;

endmodule

module line_buffer_array_k5
#(
    parameter KER_SIZE = 5,
    parameter BITWIDTH = 8,
    parameter AW       = 8,
    parameter PAD      = 1
)
(
    input logic clk,
    input logic rstn,
    input logic [BITWIDTH*KER_SIZE-1:0] pixel_in,
    input logic [3-1:0] col_ptr,
    input logic [3-1:0] init_col_ptr,
    input logic [KER_SIZE-1:0] left_pad_mask,
    input logic [KER_SIZE-1:0] right_pad_mask,
    output logic [BITWIDTH*KER_SIZE*KER_SIZE-1:0] pixel_out   
);

// wires
//logic [KER_SIZE*BITWIDTH-1:0] pixel_col [KER_SIZE-1:0];
logic [KER_SIZE*KER_SIZE*BITWIDTH-1:0] pixel_col;

//logic [KER_SIZE*BITWIDTH-1:0] pixel_row [KER_SIZE-1:0];
logic [KER_SIZE*KER_SIZE*BITWIDTH-1:0] pixel_row;

//logic [KER_SIZE*BITWIDTH-1:0] padded_pixel_row [KER_SIZE-1:0];
logic [KER_SIZE*KER_SIZE*BITWIDTH-1:0] padded_pixel_row;

//logic [KER_SIZE*BITWIDTH-1:0] left_padded_pixel_col [KER_SIZE-1:0];
logic [KER_SIZE*KER_SIZE*BITWIDTH-1:0] left_padded_pixel_col;

//logic [KER_SIZE*BITWIDTH-1:0] right_padded_pixel_col [KER_SIZE-1:0];
logic [KER_SIZE*KER_SIZE*BITWIDTH-1:0] right_padded_pixel_col; 

logic [KER_SIZE*KER_SIZE*BITWIDTH-1:0] pixel_out_wire;
logic [KER_SIZE*KER_SIZE*BITWIDTH-1:0] stored_pixel_out;
logic ready;

logic [8-1:0] global_col_ptr;
logic ready_reg;

// reg array
genvar i,j;
generate
for (i = 0; i < KER_SIZE; i++) begin: genblk_21
    d_flop #(
        .BITWIDTH (BITWIDTH*KER_SIZE)
    ) reg_inst (
        .clk (clk),
        .rstn (rstn),
        .valid (col_ptr == i),
        .D (pixel_in),
        .Q (pixel_col[(i+1)*KER_SIZE*BITWIDTH -1:i*KER_SIZE*BITWIDTH])
    ); // each d_flop stores a column of data
//always@(posedge clk) begin 
assign left_padded_pixel_col[(i+1)*KER_SIZE*BITWIDTH -1:i*KER_SIZE*BITWIDTH] = (left_pad_mask[i]==1)? {(KER_SIZE*BITWIDTH){1'b0}} : pixel_col[(i+1)*KER_SIZE*BITWIDTH -1:i*KER_SIZE*BITWIDTH];//left padding
//end
end
endgenerate

// reshape
always_comb begin
    case (1'b1)
        (col_ptr == 'd0): pixel_out_wire = {pixel_in[5*BITWIDTH-1:4*BITWIDTH],		left_padded_pixel_col[5*5*BITWIDTH-1:5*4*BITWIDTH],		left_padded_pixel_col[4*5*BITWIDTH-1:4*4*BITWIDTH],		left_padded_pixel_col[3*5*BITWIDTH-1:3*4*BITWIDTH],		left_padded_pixel_col[2*5*BITWIDTH-1:2*4*BITWIDTH],		pixel_in[4*BITWIDTH-1:3*BITWIDTH],		left_padded_pixel_col[5*4*BITWIDTH-1:5*3*BITWIDTH],		left_padded_pixel_col[4*4*BITWIDTH-1:4*3*BITWIDTH],		left_padded_pixel_col[3*4*BITWIDTH-1:3*3*BITWIDTH],		left_padded_pixel_col[2*4*BITWIDTH-1:2*3*BITWIDTH],		pixel_in[3*BITWIDTH-1:2*BITWIDTH],		left_padded_pixel_col[5*3*BITWIDTH-1:5*2*BITWIDTH],		left_padded_pixel_col[4*3*BITWIDTH-1:4*2*BITWIDTH],		left_padded_pixel_col[3*3*BITWIDTH-1:3*2*BITWIDTH],		left_padded_pixel_col[2*3*BITWIDTH-1:2*2*BITWIDTH],		pixel_in[2*BITWIDTH-1:BITWIDTH],		left_padded_pixel_col[5*2*BITWIDTH-1:5*BITWIDTH],		left_padded_pixel_col[4*2*BITWIDTH-1:4*BITWIDTH],		left_padded_pixel_col[3*2*BITWIDTH-1:3*BITWIDTH],		left_padded_pixel_col[2*2*BITWIDTH-1:2*BITWIDTH],		pixel_in[BITWIDTH-1:0],		left_padded_pixel_col[5*BITWIDTH-1:0],		left_padded_pixel_col[4*BITWIDTH-1:0],		left_padded_pixel_col[3*BITWIDTH-1:0],		left_padded_pixel_col[2*BITWIDTH-1:0]};
        (col_ptr == 'd1): pixel_out_wire = {pixel_in[5*BITWIDTH-1:4*BITWIDTH],		left_padded_pixel_col[5*BITWIDTH-1:4*BITWIDTH],		left_padded_pixel_col[5*5*BITWIDTH-1:5*4*BITWIDTH],		left_padded_pixel_col[4*5*BITWIDTH-1:4*4*BITWIDTH],		left_padded_pixel_col[3*5*BITWIDTH-1:3*4*BITWIDTH],		pixel_in[4*BITWIDTH-1:3*BITWIDTH],		left_padded_pixel_col[4*BITWIDTH-1:3*BITWIDTH],		left_padded_pixel_col[5*4*BITWIDTH-1:5*3*BITWIDTH],		left_padded_pixel_col[4*4*BITWIDTH-1:4*3*BITWIDTH],		left_padded_pixel_col[3*4*BITWIDTH-1:3*3*BITWIDTH],		pixel_in[3*BITWIDTH-1:2*BITWIDTH],		left_padded_pixel_col[3*BITWIDTH-1:2*BITWIDTH],		left_padded_pixel_col[5*3*BITWIDTH-1:5*2*BITWIDTH],		left_padded_pixel_col[4*3*BITWIDTH-1:4*2*BITWIDTH],		left_padded_pixel_col[3*3*BITWIDTH-1:3*2*BITWIDTH],		pixel_in[2*BITWIDTH-1:BITWIDTH],		left_padded_pixel_col[2*BITWIDTH-1:BITWIDTH],		left_padded_pixel_col[5*2*BITWIDTH-1:5*BITWIDTH],		left_padded_pixel_col[4*2*BITWIDTH-1:4*BITWIDTH],		left_padded_pixel_col[3*2*BITWIDTH-1:3*BITWIDTH],		pixel_in[BITWIDTH-1:0],		left_padded_pixel_col[BITWIDTH-1:0],		left_padded_pixel_col[5*BITWIDTH-1:0],		left_padded_pixel_col[4*BITWIDTH-1:0],		left_padded_pixel_col[3*BITWIDTH-1:0]};
        (col_ptr == 'd2): pixel_out_wire = {pixel_in[5*BITWIDTH-1:4*BITWIDTH],		left_padded_pixel_col[2*5*BITWIDTH-1:2*4*BITWIDTH],		left_padded_pixel_col[5*BITWIDTH-1:4*BITWIDTH],		left_padded_pixel_col[5*5*BITWIDTH-1:5*4*BITWIDTH],		left_padded_pixel_col[4*5*BITWIDTH-1:4*4*BITWIDTH],		pixel_in[4*BITWIDTH-1:3*BITWIDTH],		left_padded_pixel_col[2*4*BITWIDTH-1:2*3*BITWIDTH],		left_padded_pixel_col[4*BITWIDTH-1:3*BITWIDTH],		left_padded_pixel_col[5*4*BITWIDTH-1:5*3*BITWIDTH],		left_padded_pixel_col[4*4*BITWIDTH-1:4*3*BITWIDTH],		pixel_in[3*BITWIDTH-1:2*BITWIDTH],		left_padded_pixel_col[2*3*BITWIDTH-1:2*2*BITWIDTH],		left_padded_pixel_col[3*BITWIDTH-1:2*BITWIDTH],		left_padded_pixel_col[5*3*BITWIDTH-1:5*2*BITWIDTH],		left_padded_pixel_col[4*3*BITWIDTH-1:4*2*BITWIDTH],		pixel_in[2*BITWIDTH-1:BITWIDTH],		left_padded_pixel_col[2*2*BITWIDTH-1:2*BITWIDTH],		left_padded_pixel_col[2*BITWIDTH-1:BITWIDTH],		left_padded_pixel_col[5*2*BITWIDTH-1:5*BITWIDTH],		left_padded_pixel_col[4*2*BITWIDTH-1:4*BITWIDTH],		pixel_in[BITWIDTH-1:0],		left_padded_pixel_col[2*BITWIDTH-1:0],		left_padded_pixel_col[BITWIDTH-1:0],		left_padded_pixel_col[5*BITWIDTH-1:0],		left_padded_pixel_col[4*BITWIDTH-1:0]};
        (col_ptr == 'd3): pixel_out_wire = {pixel_in[5*BITWIDTH-1:4*BITWIDTH],		left_padded_pixel_col[3*5*BITWIDTH-1:3*4*BITWIDTH],		left_padded_pixel_col[2*5*BITWIDTH-1:2*4*BITWIDTH],		left_padded_pixel_col[5*BITWIDTH-1:4*BITWIDTH],		left_padded_pixel_col[5*5*BITWIDTH-1:5*4*BITWIDTH],		pixel_in[4*BITWIDTH-1:3*BITWIDTH],		left_padded_pixel_col[3*4*BITWIDTH-1:3*3*BITWIDTH],		left_padded_pixel_col[2*4*BITWIDTH-1:2*3*BITWIDTH],		left_padded_pixel_col[4*BITWIDTH-1:3*BITWIDTH],		left_padded_pixel_col[5*4*BITWIDTH-1:5*3*BITWIDTH],		pixel_in[3*BITWIDTH-1:2*BITWIDTH],		left_padded_pixel_col[3*3*BITWIDTH-1:3*2*BITWIDTH],		left_padded_pixel_col[2*3*BITWIDTH-1:2*2*BITWIDTH],		left_padded_pixel_col[3*BITWIDTH-1:2*BITWIDTH],		left_padded_pixel_col[5*3*BITWIDTH-1:5*2*BITWIDTH],		pixel_in[2*BITWIDTH-1:BITWIDTH],		left_padded_pixel_col[3*2*BITWIDTH-1:3*BITWIDTH],		left_padded_pixel_col[2*2*BITWIDTH-1:2*BITWIDTH],		left_padded_pixel_col[2*BITWIDTH-1:BITWIDTH],		left_padded_pixel_col[5*2*BITWIDTH-1:5*BITWIDTH],		pixel_in[BITWIDTH-1:0],		left_padded_pixel_col[3*BITWIDTH-1:0],		left_padded_pixel_col[2*BITWIDTH-1:0],		left_padded_pixel_col[BITWIDTH-1:0],		left_padded_pixel_col[5*BITWIDTH-1:0]};
        (col_ptr == 'd4): pixel_out_wire = {pixel_in[5*BITWIDTH-1:4*BITWIDTH],		left_padded_pixel_col[4*5*BITWIDTH-1:4*4*BITWIDTH],		left_padded_pixel_col[3*5*BITWIDTH-1:3*4*BITWIDTH],		left_padded_pixel_col[2*5*BITWIDTH-1:2*4*BITWIDTH],		left_padded_pixel_col[5*BITWIDTH-1:4*BITWIDTH],		pixel_in[4*BITWIDTH-1:3*BITWIDTH],		left_padded_pixel_col[4*4*BITWIDTH-1:4*3*BITWIDTH],		left_padded_pixel_col[3*4*BITWIDTH-1:3*3*BITWIDTH],		left_padded_pixel_col[2*4*BITWIDTH-1:2*3*BITWIDTH],		left_padded_pixel_col[4*BITWIDTH-1:3*BITWIDTH],		pixel_in[3*BITWIDTH-1:2*BITWIDTH],		left_padded_pixel_col[4*3*BITWIDTH-1:4*2*BITWIDTH],		left_padded_pixel_col[3*3*BITWIDTH-1:3*2*BITWIDTH],		left_padded_pixel_col[2*3*BITWIDTH-1:2*2*BITWIDTH],		left_padded_pixel_col[3*BITWIDTH-1:2*BITWIDTH],		pixel_in[2*BITWIDTH-1:BITWIDTH],		left_padded_pixel_col[4*2*BITWIDTH-1:4*BITWIDTH],		left_padded_pixel_col[3*2*BITWIDTH-1:3*BITWIDTH],		left_padded_pixel_col[2*2*BITWIDTH-1:2*BITWIDTH],		left_padded_pixel_col[2*BITWIDTH-1:BITWIDTH],		pixel_in[BITWIDTH-1:0],		left_padded_pixel_col[4*BITWIDTH-1:0],		left_padded_pixel_col[3*BITWIDTH-1:0],		left_padded_pixel_col[2*BITWIDTH-1:0],		left_padded_pixel_col[BITWIDTH-1:0]};
        default:          pixel_out_wire = '0;
    endcase
end



// output flop
always_ff @(posedge clk) begin
    if (!rstn) begin
        stored_pixel_out <= '0;
    end
    else if (ready) begin
        stored_pixel_out <= pixel_out_wire;
    end
    else begin
        stored_pixel_out <= stored_pixel_out;
    end
end

generate
	for (i = 0; i < KER_SIZE ; i++) begin: genblk_17
		assign pixel_row[(i+1)*KER_SIZE*BITWIDTH-1:i*KER_SIZE*BITWIDTH] = stored_pixel_out[KER_SIZE*BITWIDTH*i+:KER_SIZE*BITWIDTH];
		assign pixel_out[KER_SIZE*BITWIDTH*i+:KER_SIZE*BITWIDTH] = padded_pixel_row[(i+1)*KER_SIZE*BITWIDTH-1:i*KER_SIZE*BITWIDTH];
	end
endgenerate

generate
	for (i = 0; i < KER_SIZE ; i++) begin: genblk_18
	for (j = 0; j < KER_SIZE ; j++) begin: genblk_19
		assign padded_pixel_row[(i*KER_SIZE*BITWIDTH + BITWIDTH*j)+:BITWIDTH] = right_pad_mask[j] ?{BITWIDTH{1'b0}}:pixel_row[(i*KER_SIZE*BITWIDTH + BITWIDTH*j)+:BITWIDTH];
	end
	end
endgenerate

assign ready =  init_col_ptr == KER_SIZE-1;

endmodule

module line_buffer_array_k3
#(
    parameter   KER_SIZE    = 3,
    parameter BITWIDTH  = 8,
    parameter AW                = 8,
		parameter PAD = 1								 
)
(
    input logic clk,
    input logic rstn,
    input logic [BITWIDTH*KER_SIZE-1:0] pixel_in,
    input logic [3-1:0] col_ptr,
    input logic [3-1:0] init_col_ptr,
		input logic [KER_SIZE-1:0] left_pad_mask,																				 
		input logic [KER_SIZE-1:0] right_pad_mask,																					
    output logic [BITWIDTH*KER_SIZE*KER_SIZE-1:0] pixel_out   
);

// wires
//logic [KER_SIZE*BITWIDTH-1:0] pixel_col [KER_SIZE-1:0];
logic [KER_SIZE*KER_SIZE*BITWIDTH-1:0] pixel_col;

//logic [KER_SIZE*BITWIDTH-1:0] pixel_row [KER_SIZE-1:0];
logic [KER_SIZE*KER_SIZE*BITWIDTH-1:0] pixel_row;

//logic [KER_SIZE*BITWIDTH-1:0] padded_pixel_row [KER_SIZE-1:0];
logic [KER_SIZE*KER_SIZE*BITWIDTH-1:0] padded_pixel_row;

//logic [KER_SIZE*BITWIDTH-1:0] left_padded_pixel_col [KER_SIZE-1:0];
logic [KER_SIZE*KER_SIZE*BITWIDTH-1:0] left_padded_pixel_col;

//logic [KER_SIZE*BITWIDTH-1:0] right_padded_pixel_col [KER_SIZE-1:0];
logic [KER_SIZE*KER_SIZE*BITWIDTH-1:0] right_padded_pixel_col; 

logic [KER_SIZE*KER_SIZE*BITWIDTH-1:0] pixel_out_wire;
logic [KER_SIZE*KER_SIZE*BITWIDTH-1:0] stored_pixel_out;
logic ready;

logic [8-1:0] global_col_ptr;
logic ready_reg;													 
// reg array
genvar i,j;
generate
for (i = 0; i < KER_SIZE; i++) begin: genblk_22
    d_flop #(
        .BITWIDTH (BITWIDTH*KER_SIZE)
    ) reg_inst (
        .clk (clk),
        .rstn (rstn),
        .valid (col_ptr == i),
        .D (pixel_in),
        .Q (pixel_col[(i+1)*KER_SIZE*BITWIDTH -1:i*KER_SIZE*BITWIDTH])
    ); // each d_flop stores a column of data
//always@(posedge clk) begin 
assign left_padded_pixel_col[(i+1)*KER_SIZE*BITWIDTH -1:i*KER_SIZE*BITWIDTH] = (left_pad_mask[i]==1)? {(KER_SIZE*BITWIDTH){1'b0}} : pixel_col[(i+1)*KER_SIZE*BITWIDTH -1:i*KER_SIZE*BITWIDTH];//left padding
//end
end
endgenerate

// reshape
always_comb begin
    case (1'b1)
			(col_ptr == 'd0): pixel_out_wire = {pixel_in[3*BITWIDTH-1:2*BITWIDTH],left_padded_pixel_col[3*3*BITWIDTH-1:3*2*BITWIDTH],left_padded_pixel_col[2*3*BITWIDTH-1:2*2*BITWIDTH],pixel_in[2*BITWIDTH-1:BITWIDTH],left_padded_pixel_col[3*2*BITWIDTH-1:3*BITWIDTH],left_padded_pixel_col[2*2*BITWIDTH-1:2*BITWIDTH],pixel_in[BITWIDTH-1:0],left_padded_pixel_col[3*BITWIDTH-1:0],left_padded_pixel_col[2*BITWIDTH-1:0]};
			(col_ptr == 'd1): pixel_out_wire = {pixel_in[3*BITWIDTH-1:2*BITWIDTH],left_padded_pixel_col[3*BITWIDTH-1:2*BITWIDTH],left_padded_pixel_col[3*3*BITWIDTH-1:3*2*BITWIDTH],pixel_in[2*BITWIDTH-1:BITWIDTH],left_padded_pixel_col[2*BITWIDTH-1:BITWIDTH],left_padded_pixel_col[3*2*BITWIDTH-1:3*BITWIDTH],pixel_in[BITWIDTH-1:0],left_padded_pixel_col[BITWIDTH-1:0],left_padded_pixel_col[3*BITWIDTH-1:0]};
			(col_ptr == 'd2): pixel_out_wire = {pixel_in[3*BITWIDTH-1:2*BITWIDTH],left_padded_pixel_col[2*3*BITWIDTH-1:2*2*BITWIDTH],left_padded_pixel_col[3*BITWIDTH-1:2*BITWIDTH],pixel_in[2*BITWIDTH-1:BITWIDTH],left_padded_pixel_col[2*2*BITWIDTH-1:2*BITWIDTH],left_padded_pixel_col[2*BITWIDTH-1:BITWIDTH],pixel_in[BITWIDTH-1:0],left_padded_pixel_col[2*BITWIDTH-1:0],left_padded_pixel_col[BITWIDTH-1:0]};        
			default:          									pixel_out_wire = '0;
    endcase
end

// output flop
always_ff @(posedge clk) begin
    if (!rstn) begin
        stored_pixel_out <= '0;
    end
    else if (ready) begin
        stored_pixel_out <= pixel_out_wire;
    end
    else begin
        stored_pixel_out <= stored_pixel_out;
    end
end

generate
	for (i = 0; i < KER_SIZE ; i++) begin: genblk_23
		assign pixel_row[(i+1)*KER_SIZE*BITWIDTH-1:i*KER_SIZE*BITWIDTH] = stored_pixel_out[KER_SIZE*BITWIDTH*i+:KER_SIZE*BITWIDTH];
		assign pixel_out[KER_SIZE*BITWIDTH*i+:KER_SIZE*BITWIDTH] = padded_pixel_row[(i+1)*KER_SIZE*BITWIDTH-1:i*KER_SIZE*BITWIDTH];
	end
endgenerate

generate
	for (i = 0; i < KER_SIZE ; i++) begin: genblk_24
	for (j = 0; j < KER_SIZE ; j++) begin: genblk_25
		assign padded_pixel_row[(i*KER_SIZE*BITWIDTH + BITWIDTH*j)+:BITWIDTH] = right_pad_mask[j] ?{BITWIDTH{1'b0}}:pixel_row[(i*KER_SIZE*BITWIDTH + BITWIDTH*j)+:BITWIDTH];
	end
	end
endgenerate

assign ready =  init_col_ptr == KER_SIZE-1;

endmodule

module line_buffer_array_k2
#(
    parameter KER_SIZE = 3,
    parameter BITWIDTH = 8,
    parameter AW = 8
)
(
    input logic clk,
    input logic rstn,
    input logic [BITWIDTH*KER_SIZE-1:0] pixel_in,
    input logic [3-1:0] col_ptr,
    input logic [3-1:0] init_col_ptr,
    output logic [BITWIDTH*KER_SIZE*KER_SIZE-1:0] pixel_out
);

// wires
//logic [KER_SIZE*BITWIDTH-1:0] pixel_col [KER_SIZE-1:0];
logic [KER_SIZE*KER_SIZE*BITWIDTH-1:0] pixel_col;

logic [KER_SIZE*KER_SIZE*BITWIDTH-1:0] pixel_out_wire;
logic ready;

// reg array
genvar i;
generate
for (i=0;i<KER_SIZE;i++) begin: genblk_30
    d_flop #(
        .BITWIDTH (BITWIDTH*KER_SIZE)
    ) reg_inst (
        .clk (clk),
        .rstn (rstn),
        .valid (col_ptr == i),
        .D (pixel_in),
        .Q (pixel_col[(i+1)*KER_SIZE*BITWIDTH -1:i*KER_SIZE*BITWIDTH])
    ); // each d_flop stores a column of data
end
endgenerate

// reshape
always_comb begin
    case (1'b1)
        (col_ptr == 'd0): pixel_out_wire = {pixel_in[2*BITWIDTH-1:BITWIDTH],pixel_col[2*2*BITWIDTH-1:2*BITWIDTH],pixel_in[BITWIDTH-1:0],pixel_col[2*BITWIDTH-1:0]};
        (col_ptr == 'd1): pixel_out_wire = {pixel_in[2*BITWIDTH-1:BITWIDTH],pixel_col[2*BITWIDTH-1:BITWIDTH],pixel_in[BITWIDTH-1:0],pixel_col[BITWIDTH-1:0]};
        default:          pixel_out_wire = '0;
    endcase
end

// output flop
always_ff @(posedge clk) begin
    if (!rstn) begin
        pixel_out <= '0;
    end
    else if (ready) begin
        pixel_out <= pixel_out_wire;
    end
    else begin
        pixel_out <= pixel_out;
    end
end

assign ready = (init_col_ptr == KER_SIZE-1);

endmodule

// d_flop
module d_flop
#(
    parameter BITWIDTH = 8
)
(
    input logic clk,
    input logic rstn,
    input logic valid,
    input logic [BITWIDTH-1:0] D,
    output logic [BITWIDTH-1:0] Q
);

always_ff @(posedge clk) begin
    if (rstn == 0) begin
        Q <= '0;
    end
    else if (valid == 1) begin
        Q <= D;
    end
    else begin
        Q <= Q;
    end     
end

endmodule





module line_buffer_controller
#(
    parameter KER_SIZE    = 3,
    parameter INPUT_X_DIM = 3,
    parameter PAD         = 1
)
(
    input logic clk,
    input logic rstn,
    input logic valid,
    input logic row_complete,
    output logic right_pad_valid,
    output logic [3-1:0] col_ptr,
    output logic [KER_SIZE-1:0] left_pad_mask,	 
    output logic [KER_SIZE-1:0] right_pad_mask,	 
    output logic [3-1:0] init_col_ptr
);

logic [3-1:0] init_col_ptr_nxt;
logic [3-1:0] col_ptr_nxt;

logic [7:0] global_col_ptr;
logic [7:0] global_col_ptr_nxt;

//-------------------------------------
logic padrow_complete;
logic row_complete_D1;
logic row_complete_D2;
always_ff @(posedge clk) 
begin
	if (!rstn) 
	begin
			row_complete_D1 	 <='0;
			row_complete_D2 	 <='0;
	end
	else if (padrow_complete)
	begin	
			row_complete_D1 		<= '0;
			row_complete_D2 		<= '0;
	end
	else
	begin
			row_complete_D1 		<= row_complete;
			row_complete_D2 		<= row_complete_D1;
	end
end
assign padrow_complete = row_complete_D1;
//-------------------------------------


// initialize counters
always_ff @(posedge clk) begin
    if (!rstn) begin
        col_ptr 			      <= PAD;//Left padding
        init_col_ptr 		    <= PAD;//Left padding
        global_col_ptr 		  <='0;
    end
    else if (padrow_complete) begin
        col_ptr 				    <= PAD; //Left padding
        init_col_ptr 			  <= PAD;//Left padding
        global_col_ptr 			<= '0;
    end
    else begin
        col_ptr 				    <= col_ptr_nxt;
        init_col_ptr 			  <= init_col_ptr_nxt;
        global_col_ptr 			<= global_col_ptr_nxt;
    end
end


// Increment counters based on conditions
assign col_ptr_nxt 		  	= valid ? (col_ptr==KER_SIZE-1 ? '0 : col_ptr + 1'd1) : col_ptr;
assign global_col_ptr_nxt = padrow_complete ? 'd0 : valid ?  global_col_ptr + 1'd1: global_col_ptr;
assign init_col_ptr_nxt   = valid && init_col_ptr<KER_SIZE-1 ? init_col_ptr + 1'd1 :padrow_complete==1'b1 ? PAD : init_col_ptr;

// Left pad logic
logic [KER_SIZE-1:0]left_pad_shift;

generate
	if(PAD>0) 
	begin
		logic [PAD-1:0] shifted_left_pad_mask;
		always_ff @(posedge clk) 
		begin
			if (!rstn) 
				shifted_left_pad_mask <= {PAD{1'b1}}; 
			else if (padrow_complete) 
				shifted_left_pad_mask <= {PAD{1'b1}}; 
			else if (valid)
				shifted_left_pad_mask <= shifted_left_pad_mask << left_pad_shift; 
			else
				shifted_left_pad_mask <= shifted_left_pad_mask; 
		end
	assign left_pad_mask =  {{KER_SIZE-PAD{1'b0}},shifted_left_pad_mask};
	end
	
	else
	begin
		assign left_pad_mask =  {KER_SIZE{1'b0}};
	end
endgenerate
	
assign left_pad_shift  = global_col_ptr >= KER_SIZE-PAD-1 && global_col_ptr < KER_SIZE-1 ? 1'b1 : 1'b0;

// Right pad logic
logic right_pad_en;
logic [2:0] right_pad_counter;
logic [KER_SIZE-1:0]right_pad_shift;

always_ff @(posedge clk) begin
    if (!rstn) begin
        right_pad_en <= '0;
    end
    else if (global_col_ptr==INPUT_X_DIM-PAD-1) begin
        right_pad_en <= '1;
    end
    else if(right_pad_counter==KER_SIZE-1)begin //PAD + (KER_SIZE-PAD-1)
        right_pad_en <= 0;
    end
end

always_ff @(posedge clk) begin
    if (!rstn) begin
        right_pad_counter <= '0;
    end
    else if (right_pad_counter==KER_SIZE-1) begin
        right_pad_counter <= 0;
    end
    else if (right_pad_en) begin
        right_pad_counter <= right_pad_counter + 1'd1;
    end
    else 
        right_pad_counter <= 0;
end

assign right_pad_shift =  right_pad_en && !(right_pad_counter<PAD+1);
assign right_pad_valid = right_pad_shift;

generate
	if(PAD>0) 
	begin
		logic [KER_SIZE-1:0] right_pad_mask_wire;
		always_ff @(posedge clk) 
		begin
			if (!rstn) 
				right_pad_mask_wire <=  {1'b1,{KER_SIZE-1{1'b0}}};
			else if (global_col_ptr==INPUT_X_DIM-PAD-1) 
				right_pad_mask_wire <=  {1'b1,{KER_SIZE-1{1'b0}}};
			else if (right_pad_shift)
				right_pad_mask_wire <= (right_pad_mask_wire >> 1) | {1'b1,{KER_SIZE-1{1'b0}}};
			else
				right_pad_mask_wire <= {1'b1,{KER_SIZE-1{1'b0}}};
		end
		assign right_pad_mask = right_pad_shift ? right_pad_mask_wire: 0;
	end
	
	else
	begin
		assign right_pad_mask =  {KER_SIZE{1'b0}};
	end
endgenerate
endmodule




module sram_array_k3
#(
    parameter KER_SIZE = 3,
    parameter DW       = 32, // Data width (nbits)
    parameter NW       = 32, // Number of words
    parameter AW       = $clog2(NW)
)
(
    input logic clk,
    input logic rstn,
    input logic [AW-1:0] a, // same for read and write    
    input logic [KER_SIZE-1:0] wen, // active high
    input logic [KER_SIZE-1:0] ren, // active high
    input logic [DW-1:0] d,
    output logic [(KER_SIZE-1)*DW-1:0] q
);

//logic [DW-1:0] q_wire [KER_SIZE-1:0];
logic [KER_SIZE*DW-1:0] q_wire; 

logic [KER_SIZE-1:0] write_en_D1;

always_ff @(posedge clk) begin
    if(!rstn) begin
        write_en_D1 <= '0;
    end
    else begin
        write_en_D1 <= wen;
    end
end

genvar i;
generate
    for (i = 0; i < (KER_SIZE); i++) begin: genblk_26
        array #(
            .DW (DW),
            .NW (NW),
            .AW (AW)
        ) sram_inst (
            .clk (clk),
            .cen (!(wen[i] || ren[i])),
            .gwen (!(wen[i])),
            .a (a),
            .d (d),
            .q (q_wire[(i+1)*DW-1:i*DW])
        );
    end
endgenerate

// reorder rows
always_comb begin
    case (1'b1)
        write_en_D1[0] : q = {q_wire[3*DW-1:2*DW],q_wire[2*DW-1:DW]};
        write_en_D1[1] : q = {q_wire[DW-1:0],q_wire[3*DW-1:2*DW]};
        write_en_D1[2] : q = {q_wire[2*DW-1:DW],q_wire[DW-1:0]};
        default :        q = '0;
    endcase
end

endmodule

module sram_array_k5
#(
    parameter KER_SIZE = 5,
    parameter DW = 32, // Data width (nbits)
    parameter NW = 32, // Number of words
    parameter AW = $clog2(NW)
)
(
    input logic clk,
    input logic rstn,
    input logic [AW-1:0] a, // same for read and write    
    input logic [KER_SIZE-1:0] wen, // active high
    input logic [KER_SIZE-1:0] ren, // active high
    input logic [DW-1:0] d,
    output logic [(KER_SIZE-1)*DW-1:0] q
);

//logic [DW-1:0] q_wire [KER_SIZE-1:0];
logic [KER_SIZE*DW-1:0] q_wire; 

logic [KER_SIZE-1:0] write_en_D1; // delayed write enable because of 1 cycle delay of sram

always_ff @(posedge clk) begin
    if(!rstn) begin
        write_en_D1 <= '0;
    end
    else begin
        write_en_D1 <= wen;
    end
end

genvar i;
generate
    for (i = 0; i < (KER_SIZE); i++) begin: genblk_27
        array #(
            .DW (DW),
            .NW (NW),
            .AW (AW)
        ) sram_inst (
            .clk (clk),
            .cen (!(wen[i] || ren[i])),
            .gwen (!(wen[i])),
            .a (a),
            .d (d),
            .q (q_wire[(i+1)*DW-1:i*DW])
        );
    end
endgenerate

// reorder rows
always_comb begin
    case (1'b1)
        write_en_D1[0] : q = {q_wire[5*DW-1:4*DW],q_wire[4*DW-1:3*DW],q_wire[3*DW-1:2*DW],q_wire[2*DW-1:DW]};
        write_en_D1[1] : q = {q_wire[DW-1:0],q_wire[5*DW-1:4*DW],q_wire[4*DW-1:3*DW],q_wire[3*DW-1:2*DW]};
        write_en_D1[2] : q = {q_wire[2*DW-1:DW],q_wire[DW-1:0],q_wire[5*DW-1:4*DW],q_wire[4*DW-1:3*DW]};
        write_en_D1[3] : q = {q_wire[3*DW-1:2*DW],q_wire[2*DW-1:DW],q_wire[DW-1:DW],q_wire[5*DW-1:4*DW]};
        write_en_D1[4] : q = {q_wire[4*DW-1:3*DW],q_wire[3*DW-1:2*DW],q_wire[2*DW-1:DW],q_wire[DW-1:0]};
        default :        q = '0;
    endcase
end

endmodule

module sram_array_k7
#(
    parameter KER_SIZE = 7,
    parameter DW = 32, // Data width (nbits)
    parameter NW = 32, // Number of words
    parameter AW = $clog2(NW)
)
(
    input logic clk,
    input logic rstn,
    input logic [AW-1:0] a, // same for read and write    
    input logic [KER_SIZE-1:0] wen, // active high
    input logic [KER_SIZE-1:0] ren, // active high
    input logic [DW-1:0] d,
    output logic [(KER_SIZE-1)*DW-1:0] q
);

//logic [DW-1:0] q_wire [KER_SIZE-1:0];
logic [KER_SIZE*DW-1:0] q_wire; 

logic [KER_SIZE-1:0] write_en_D1; // delayed write enable because of 1 cycle delay of sram

always_ff @(posedge clk) begin
    if(!rstn) begin
        write_en_D1 <= '0;
    end
    else begin
        write_en_D1 <= wen;
    end
end

genvar i;
generate
    for (i = 0; i < (KER_SIZE); i++) begin: genblk_28
        array #(
            .DW (DW),
            .NW (NW),
            .AW (AW)
        ) sram_inst (
            .clk (clk),
            .cen (!(wen[i] || ren[i])),
            .gwen (!(wen[i])),
            .a (a),
            .d (d),
            .q (q_wire[(i+1)*DW-1:i*DW])
        );
    end
endgenerate

// reorder rows
always_comb begin
    case (1'b1) 
        write_en_D1[0] : q = {q_wire[7*DW-1:6*DW],q_wire[6*DW-1:5*DW],q_wire[5*DW-1:4*DW],q_wire[4*DW-1:3*DW],q_wire[3*DW-1:2*DW],q_wire[2*DW-1:DW]};
        write_en_D1[1] : q = {q_wire[DW-1:0],q_wire[7*DW-1:6*DW],q_wire[6*DW-1:5*DW],q_wire[5*DW-1:4*DW],q_wire[4*DW-1:3*DW],q_wire[3*DW-1:2*DW]};
        write_en_D1[2] : q = {q_wire[2*DW-1:DW],q_wire[DW-1:0],q_wire[7*DW-1:6*DW],q_wire[6*DW-1:5*DW],q_wire[5*DW-1:4*DW],q_wire[4*DW-1:3*DW]};
        write_en_D1[3] : q = {q_wire[3*DW-1:2*DW],q_wire[2*DW-1:DW],q_wire[DW-1:0],q_wire[7*DW-1:6*DW],q_wire[6*DW-1:5*DW],q_wire[5*DW-1:4*DW]};
        write_en_D1[4] : q = {q_wire[4*DW-1:3*DW],q_wire[3*DW-1:2*DW],q_wire[2*DW-1:DW],q_wire[DW-1:0],q_wire[7*DW-1:6*DW],q_wire[6*DW-1:5*DW]};
        write_en_D1[5] : q = {q_wire[5*DW-1:4*DW],q_wire[4*DW-1:3*DW],q_wire[3*DW-1:2*DW],q_wire[2*DW-1:DW],q_wire[DW-1:0],q_wire[7*DW-1:6*DW]};
        write_en_D1[6] : q = {q_wire[6*DW-1:5*DW],q_wire[5*DW-1:4*DW],q_wire[4*DW-1:3*DW],q_wire[3*DW-1:2*DW],q_wire[2*DW-1:DW],q_wire[DW-1:0]};
        default :        q = '0;
    endcase
end

endmodule

module sram_array_k2
#(
    parameter KER_SIZE = 3,
    parameter DW = 32, // Data width (nbits)
    parameter NW = 32, // Number of words
    parameter AW = $clog2(NW)
)
(
    input logic clk,
    input logic rstn,
    input logic [AW-1:0] a, // same for read and write
    input logic [KER_SIZE-1:0] wen, // active high
    input logic [KER_SIZE-1:0] ren, // active high
    input logic [DW-1:0] d,
    output logic [(KER_SIZE-1)*DW-1:0] q
);

//logic [DW-1:0] q_wire [KER_SIZE-1:0];
logic [KER_SIZE*DW-1:0] q_wire; 

logic [KER_SIZE-1:0] write_en_D1;

always_ff @(posedge clk ) begin
    if(!rstn) begin
        write_en_D1 <= '0;
    end
    else begin
        write_en_D1 <= wen;
    end
end

genvar i;
generate
    for (i = 0; i < (KER_SIZE); i++) begin: genblk_29
        array #(
            .DW (DW),
            .NW (NW),
            .AW (AW)
        ) sram_inst (
            .clk (clk),
            .cen (!(wen[i] || ren[i])),
            .gwen (!(wen[i])),
            .a (a),
            .d (d),
            .q (q_wire[(i+1)*DW-1:i*DW])
        );
    end
endgenerate

// reorder rows
always_comb
begin
    case (1'b1)
        write_en_D1[0] : q = {q_wire[1]};
        write_en_D1[1] : q = {q_wire[0]};
        default :        q = '0;
    endcase
end

endmodule

module array
#(
    parameter DW = 32,
    parameter NW = 32,
    parameter AW = $clog2(NW) 
) 
(
    input logic clk,
    input logic cen, // enable active low
    input logic gwen, // global write enable active low
    input logic [AW-1:0] a,
    input logic [DW-1:0] d,
    output logic [DW-1:0] q
);

logic [DW-1:0] data [0:NW-1];

// write
always @(posedge clk) begin
    if (~cen & ~gwen) begin
        data[a] <= d;
    end
    else begin
        data[a] <= data[a];
    end
end

// read
always @(posedge clk) begin
    if (~cen) begin
        q <= data[a];
    end
    else begin
        q <= q;
    end
end

endmodule

module ram_single #(parameter WORDS = 256, 
                    parameter A_WIDTH =8, 
                    parameter D_WIDTH=12,
                    parameter INIT_FILE="dummy.mif") (q, address, d, we, clk);
   output [D_WIDTH-1:0] q;
   input [D_WIDTH-1:0] d;
   input [A_WIDTH:0] address;
   input we, clk;

`ifdef hard_mem

defparam u_single_port_ram.ADDR_WIDTH = A_WIDTH;
defparam u_single_port_ram.DATA_WIDTH = D_WIDTH;

single_port_ram u_single_port_ram(
.addr(address),
.we(we),
.data(d),
.out(q),
.clk(clk)
);

`elsif QUARTUS
    reg [D_WIDTH-1:0] mem [WORDS-1:0];
    reg [D_WIDTH-1:0] q;

    initial begin
        $readmemb(INIT_FILE, mem);
    end

    always @(posedge clk) begin
        q <= mem[address];
    end

`else

    reg [D_WIDTH-1:0] mem [WORDS-1:0];
    reg [D_WIDTH-1:0] q;
    always @(posedge clk) begin
        if (we)
            mem[address] <= d;
        q <= mem[address];
    end

`endif
endmodule

module sram_controller
#(
    parameter KER_SIZE    = 3,
    parameter BITWIDTH    = 8,
    parameter STRIDE      = 8,
    parameter NFMAPS      = 3,
    parameter INPUT_X_DIM = 28,
    parameter PAD         = 1,
    parameter AW          = 5
)
(
  input logic clk,      
  input logic rstn,     
  input logic valid,
  output logic [AW-1:0] addr, // same for read and write    
  output logic [KER_SIZE-1:0] write_en,     
  output logic [KER_SIZE-1:0] read_en,
  output logic ready,
  output logic [KER_SIZE-1:0] top_pad_mask ,
  output logic bottom_pad_mask,
  output logic row_is_complete
);

genvar i;

logic [KER_SIZE:0] row_ptr          ;
logic [KER_SIZE:0] pad_row_ptr      ;
logic [7:0] global_row_ptr          ;
logic [7:0] global_row_ptr_nxt      ;
logic [AW-1:0] col_ptr              ;
logic [3:0] init_row_counter        ;
logic [KER_SIZE:0] row_ptr_nxt      ;
logic [AW-1:0] col_ptr_nxt          ;
logic [3:0] init_row_counter_nxt    ;
logic [3-1:0] row_stride_counter    ;
logic [3-1:0] row_stride_counter_nxt;

//padding
logic [KER_SIZE-1:0]top_pad_shift;
logic [KER_SIZE-1:0] init_top_pad_mask;

always_ff @(posedge clk) begin
    if (!rstn) begin
        row_ptr 			      <= PAD;//top padding
        global_row_ptr 		  <= 'd0;
        col_ptr 			      <= 'd0;
        init_row_counter 	  <= PAD;//top padding
        row_stride_counter 	<= 'd0;
    end
    else begin
        row_ptr 			      <= row_ptr_nxt;
        global_row_ptr 		  <= global_row_ptr_nxt;
        col_ptr 			      <= col_ptr_nxt;
        init_row_counter 	  <= init_row_counter_nxt;
        row_stride_counter 	<= row_stride_counter_nxt;
    end
end

generate
    for (i=0;i<KER_SIZE;i++) begin: genblk_31
        assign write_en[i] = (row_ptr==i); 
    end
endgenerate

logic col_ptr_done;
logic top_pad_en;
assign col_ptr_done           = col_ptr==(INPUT_X_DIM-1);

assign row_is_complete  	    = valid && col_ptr_done;
assign col_ptr_nxt 			      = valid ? (col_ptr_done ? 'd0 : col_ptr + 1'd1) : col_ptr ; 
assign row_ptr_nxt 			      = valid && col_ptr_done ? (row_ptr==KER_SIZE-1 ? 'd0 : row_ptr + 1'd1): row_ptr;
assign global_row_ptr_nxt 	  = valid && col_ptr_done ?  global_row_ptr + 1'd1 : global_row_ptr;
assign init_row_counter_nxt   = valid && col_ptr_done && (init_row_counter<KER_SIZE-1) 	? init_row_counter + 1'd1 : init_row_counter;

assign read_en 	              = {KER_SIZE{init_row_counter == KER_SIZE-1}} & (~write_en); 
assign addr 	                = col_ptr;
assign ready 	                = (init_row_counter == KER_SIZE-1) && (row_stride_counter==0);
assign row_stride_counter_nxt = (col_ptr==(INPUT_X_DIM-1) && valid && init_row_counter == KER_SIZE-1) ? ((row_stride_counter<STRIDE-1'd1)?row_stride_counter+1'd1:'0 ): row_stride_counter;

generate
if(PAD>0)
	begin
		always_ff @(posedge clk) 
			begin
				if (!rstn) 
					top_pad_en   <= 1'd0; 
				else 
					top_pad_en   <= valid && col_ptr_done; 
			end
			
		always_ff @(posedge clk) 
			begin
				if (!rstn) 
					top_pad_mask <= init_top_pad_mask; 
				else if (top_pad_en)
					top_pad_mask <= top_pad_mask >> top_pad_shift; 
				else
					top_pad_mask <= top_pad_mask; 
			end
			
	assign bottom_pad_mask 	= global_row_ptr > INPUT_X_DIM - 1'd1; // tell line buffer that one row is done, pad zeros if needed at the bottom rows
	assign top_pad_shift 		= global_row_ptr > KER_SIZE-PAD && global_row_ptr <KER_SIZE+1 ? 1'b1 : 1'b0;
	
	end
else 
	begin
		assign top_pad_mask 		= 0;
		assign bottom_pad_mask 	= 0;
		assign top_pad_en 			= 0;
		assign top_pad_shift 		= 0;
	end
endgenerate
		
generate
	for (i=0;i<KER_SIZE;i++) 
	begin: genblk_32
		always_ff @(posedge clk) begin
			if (!rstn) 
				init_top_pad_mask[i] <= i<PAD ? 1'b1 : 1'd0; 
			else 
				init_top_pad_mask[i] <= init_top_pad_mask[i];
		end
    end
endgenerate

endmodule

`ifdef complex_dsp
module int_sop_4_wrapper (
  mode_sigs,
	clk,
	reset,
	ax,
	ay,
	bx,
	by,
  cx,
  cy,
  dx,
  dy,
	chainin,
	result,
	chainout);
input [11:0] mode_sigs;
input clk;
input reset; 
input [8:0] ax, bx, cx, dx;
input [8:0] ay, by, cy, dy;
input [63:0] chainin;
output [63:0] result;
output [63:0] chainout;

int_sop_4 int_sop_4_inst(.clk(clk),.reset(rstn),.mode_sigs(mode_sigs),.ax(ax),.ay(ay),.bx(bx),.by(by),.cx(cx),.cy(cy),.dx(dx),.dy(dy),.chainin(chainin),.result(result),.chainout(chainout));
endmodule
`else
module int_sop_4_wrapper (mode_sigs,
	clk,
	reset,
	ax,
	ay,
	bx,
	by,
  cx,
  cy,
  dx,
  dy,
	chainin,
	result,
	chainout);
input [11:0] mode_sigs;
input clk;
input reset; 
input [8:0] ax, bx, cx, dx;
input [8:0] ay, by, cy, dy;
input [63:0] chainin;
output [63:0] result;
output [63:0] chainout;

reg [8:0] ax_reg;
reg [8:0] ay_reg;
reg [8:0] bx_reg;
reg [8:0] by_reg;
reg [8:0] cx_reg;
reg [8:0] cy_reg;
reg [8:0] dx_reg;
reg [8:0] dy_reg;
reg [63:0] resulta;

reg [17:0] result_a;
reg [17:0] result_b;
reg [17:0] result_c;
reg [17:0] result_d;

always @(posedge clk) begin
  if(reset) begin
    resulta <= 0;
    ax_reg <= 0;
    ay_reg <= 0;
    bx_reg <= 0;
    by_reg <= 0;
    cx_reg <= 0;
    cy_reg <= 0;
    dx_reg <= 0;
    dy_reg <= 0;
  end
  else begin
    ax_reg <= ax;
    ay_reg <= ay;
    bx_reg <= bx;
    by_reg <= by;
    cx_reg <= cx;
    cy_reg <= cy;
    dx_reg <= dx;
    dy_reg <= dy;
    result_a <= ax_reg * ay_reg;
    result_b <= bx_reg * by_reg;
    result_c <= cx_reg * cy_reg;
    result_d <= dx_reg * dy_reg;
    resulta <= result_a + result_b + result_c + result_d + chainin;
  end
end
assign result = resulta;
assign chainout = resulta;
endmodule
`endif


