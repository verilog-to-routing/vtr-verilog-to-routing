`define BINARY_OP(out,a,b) bufif1(out, a, b);
`include "../.generic/wire_test.v"