module and_primitive();
	/*  input declaration	*/
	wire   a;
	wire   b;

	/*	output declaration	*/
	wire	out;

    assign out = a&b; 

endmodule