`define BINARY_OP(out,a,b) or(out, a, b);
`include "wire_test.v"