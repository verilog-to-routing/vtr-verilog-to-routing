`define BINARY_OP(out,a,b) xor(out, a, b);
`include "wire_test.v"