module Fadder_(
  in1,
  in2,
  in3,
  sum,
  carry);

  input in1, in2, in3;
  output sum, carry;

  assign sum=in1^in2^in3;
  assign carry=(in1&in2) | (in2&in3) | (in1&in3);

endmodule 

module Hadder_(
  in1,
  in2,
  sum,
  carry);

  input in1, in2;
  output sum, carry;

  assign sum=in1^in2;
  assign carry=in1&in2;

endmodule 

module mult_(
  a,
  b,
  s,
  c);

  input [63:0] a;
  input [63:0] b;
  output [127:0] s;
  output [126:0] c;

  wire [63:0] a_;
  wire sign_ ;
  reg [65:0] P_0 ;
  reg [65:0] P_1 ;
  reg [65:0] P_2 ;
  reg [65:0] P_3 ;
  reg [65:0] P_4 ;
  reg [65:0] P_5 ;
  reg [65:0] P_6 ;
  reg [65:0] P_7 ;
  reg [65:0] P_8 ;
  reg [65:0] P_9 ;
  reg [65:0] P_10 ;
  reg [65:0] P_11 ;
  reg [65:0] P_12 ;
  reg [65:0] P_13 ;
  reg [65:0] P_14 ;
  reg [65:0] P_15 ;
  reg [65:0] P_16 ;
  reg [65:0] P_17 ;
  reg [65:0] P_18 ;
  reg [65:0] P_19 ;
  reg [65:0] P_20 ;
  reg [65:0] P_21 ;
  reg [65:0] P_22 ;
  reg [65:0] P_23 ;
  reg [65:0] P_24 ;
  reg [65:0] P_25 ;
  reg [65:0] P_26 ;
  reg [65:0] P_27 ;
  reg [65:0] P_28 ;
  reg [65:0] P_29 ;
  reg [65:0] P_30 ;
  reg [65:0] P_31 ;
  reg [63:0] inc ;

  assign sign_ = 1'b1 ;
  assign a_ = ~ a ;

  always @( a or b or a_ )
    begin

    case( b[1:0] ) // synopsys full_case parallel_case
      2'b00:
        begin
        inc[0]=1'b0 ;
        inc[1]=1'b0 ;
        P_0={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      2'b01:
        begin
        inc[0]=1'b0 ;
        inc[1]=1'b0 ;
        P_0={(~a[63]),a[63],a} ;
        end
      2'b10:
        begin
        inc[0]=1'b0 ;
        inc[1]=1'b1 ;
        P_0={(~a_[63]),a_,1'b0} ;
        end
      2'b11:
        begin
        inc[0]=1'b1 ;
        inc[1]=1'b0 ;
        P_0={(~a_[63]),a_[63],a_} ;
        end
    endcase

    case({b[3:1]}) // synopsys full_case parallel_case
      3'b000:
        begin
        inc[2]=1'b0 ;
        inc[3]=1'b0 ;
        P_1={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b111:
        begin
        inc[2]=1'b0 ;
        inc[3]=1'b0 ;
        P_1={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b001:
        begin
        inc[2]=1'b0 ;
        inc[3]=1'b0 ;
        P_1={(~a[63]),a[63],a} ;
        end
      3'b010:
        begin
        inc[2]=1'b0 ;
        inc[3]=1'b0 ;
        P_1={(~a[63]),a[63],a} ;
        end
      3'b100:
        begin
        inc[2]=1'b0 ;
        inc[3]=1'b1 ;
        P_1={(~a_[63]),a_,1'b0} ;
        end
      3'b101:
        begin
        inc[2]=1'b1 ;
        inc[3]=1'b0 ;
        P_1={(~a_[63]),a_[63],a_} ;
        end
      3'b110:
        begin
        inc[2]=1'b1 ;
        inc[3]=1'b0 ;
        P_1={(~a_[63]),a_[63],a_} ;
        end
      3'b011:
        begin
        inc[2]=1'b0 ;
        inc[3]=1'b0 ;
        P_1={(~a[63]),a,1'b0} ;
        end
    endcase

    case({b[5:3]}) // synopsys full_case parallel_case
      3'b000:
        begin
        inc[4]=1'b0 ;
        inc[5]=1'b0 ;
        P_2={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b111:
        begin
        inc[4]=1'b0 ;
        inc[5]=1'b0 ;
        P_2={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b001:
        begin
        inc[4]=1'b0 ;
        inc[5]=1'b0 ;
        P_2={(~a[63]),a[63],a} ;
        end
      3'b010:
        begin
        inc[4]=1'b0 ;
        inc[5]=1'b0 ;
        P_2={(~a[63]),a[63],a} ;
        end
      3'b100:
        begin
        inc[4]=1'b0 ;
        inc[5]=1'b1 ;
        P_2={(~a_[63]),a_,1'b0} ;
        end
      3'b101:
        begin
        inc[4]=1'b1 ;
        inc[5]=1'b0 ;
        P_2={(~a_[63]),a_[63],a_} ;
        end
      3'b110:
        begin
        inc[4]=1'b1 ;
        inc[5]=1'b0 ;
        P_2={(~a_[63]),a_[63],a_} ;
        end
      3'b011:
        begin
        inc[4]=1'b0 ;
        inc[5]=1'b0 ;
        P_2={(~a[63]),a,1'b0} ;
        end
    endcase

    case({b[7:5]}) // synopsys full_case parallel_case
      3'b000:
        begin
        inc[6]=1'b0 ;
        inc[7]=1'b0 ;
        P_3={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b111:
        begin
        inc[6]=1'b0 ;
        inc[7]=1'b0 ;
        P_3={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b001:
        begin
        inc[6]=1'b0 ;
        inc[7]=1'b0 ;
        P_3={(~a[63]),a[63],a} ;
        end
      3'b010:
        begin
        inc[6]=1'b0 ;
        inc[7]=1'b0 ;
        P_3={(~a[63]),a[63],a} ;
        end
      3'b100:
        begin
        inc[6]=1'b0 ;
        inc[7]=1'b1 ;
        P_3={(~a_[63]),a_,1'b0} ;
        end
      3'b101:
        begin
        inc[6]=1'b1 ;
        inc[7]=1'b0 ;
        P_3={(~a_[63]),a_[63],a_} ;
        end
      3'b110:
        begin
        inc[6]=1'b1 ;
        inc[7]=1'b0 ;
        P_3={(~a_[63]),a_[63],a_} ;
        end
      3'b011:
        begin
        inc[6]=1'b0 ;
        inc[7]=1'b0 ;
        P_3={(~a[63]),a,1'b0} ;
        end
    endcase

    case({b[9:7]}) // synopsys full_case parallel_case
      3'b000:
        begin
        inc[8]=1'b0 ;
        inc[9]=1'b0 ;
        P_4={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b111:
        begin
        inc[8]=1'b0 ;
        inc[9]=1'b0 ;
        P_4={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b001:
        begin
        inc[8]=1'b0 ;
        inc[9]=1'b0 ;
        P_4={(~a[63]),a[63],a} ;
        end
      3'b010:
        begin
        inc[8]=1'b0 ;
        inc[9]=1'b0 ;
        P_4={(~a[63]),a[63],a} ;
        end
      3'b100:
        begin
        inc[8]=1'b0 ;
        inc[9]=1'b1 ;
        P_4={(~a_[63]),a_,1'b0} ;
        end
      3'b101:
        begin
        inc[8]=1'b1 ;
        inc[9]=1'b0 ;
        P_4={(~a_[63]),a_[63],a_} ;
        end
      3'b110:
        begin
        inc[8]=1'b1 ;
        inc[9]=1'b0 ;
        P_4={(~a_[63]),a_[63],a_} ;
        end
      3'b011:
        begin
        inc[8]=1'b0 ;
        inc[9]=1'b0 ;
        P_4={(~a[63]),a,1'b0} ;
        end
    endcase

    case({b[11:9]}) // synopsys full_case parallel_case
      3'b000:
        begin
        inc[10]=1'b0 ;
        inc[11]=1'b0 ;
        P_5={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b111:
        begin
        inc[10]=1'b0 ;
        inc[11]=1'b0 ;
        P_5={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b001:
        begin
        inc[10]=1'b0 ;
        inc[11]=1'b0 ;
        P_5={(~a[63]),a[63],a} ;
        end
      3'b010:
        begin
        inc[10]=1'b0 ;
        inc[11]=1'b0 ;
        P_5={(~a[63]),a[63],a} ;
        end
      3'b100:
        begin
        inc[10]=1'b0 ;
        inc[11]=1'b1 ;
        P_5={(~a_[63]),a_,1'b0} ;
        end
      3'b101:
        begin
        inc[10]=1'b1 ;
        inc[11]=1'b0 ;
        P_5={(~a_[63]),a_[63],a_} ;
        end
      3'b110:
        begin
        inc[10]=1'b1 ;
        inc[11]=1'b0 ;
        P_5={(~a_[63]),a_[63],a_} ;
        end
      3'b011:
        begin
        inc[10]=1'b0 ;
        inc[11]=1'b0 ;
        P_5={(~a[63]),a,1'b0} ;
        end
    endcase

    case({b[13:11]}) // synopsys full_case parallel_case
      3'b000:
        begin
        inc[12]=1'b0 ;
        inc[13]=1'b0 ;
        P_6={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b111:
        begin
        inc[12]=1'b0 ;
        inc[13]=1'b0 ;
        P_6={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b001:
        begin
        inc[12]=1'b0 ;
        inc[13]=1'b0 ;
        P_6={(~a[63]),a[63],a} ;
        end
      3'b010:
        begin
        inc[12]=1'b0 ;
        inc[13]=1'b0 ;
        P_6={(~a[63]),a[63],a} ;
        end
      3'b100:
        begin
        inc[12]=1'b0 ;
        inc[13]=1'b1 ;
        P_6={(~a_[63]),a_,1'b0} ;
        end
      3'b101:
        begin
        inc[12]=1'b1 ;
        inc[13]=1'b0 ;
        P_6={(~a_[63]),a_[63],a_} ;
        end
      3'b110:
        begin
        inc[12]=1'b1 ;
        inc[13]=1'b0 ;
        P_6={(~a_[63]),a_[63],a_} ;
        end
      3'b011:
        begin
        inc[12]=1'b0 ;
        inc[13]=1'b0 ;
        P_6={(~a[63]),a,1'b0} ;
        end
    endcase

    case({b[15:13]}) // synopsys full_case parallel_case
      3'b000:
        begin
        inc[14]=1'b0 ;
        inc[15]=1'b0 ;
        P_7={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b111:
        begin
        inc[14]=1'b0 ;
        inc[15]=1'b0 ;
        P_7={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b001:
        begin
        inc[14]=1'b0 ;
        inc[15]=1'b0 ;
        P_7={(~a[63]),a[63],a} ;
        end
      3'b010:
        begin
        inc[14]=1'b0 ;
        inc[15]=1'b0 ;
        P_7={(~a[63]),a[63],a} ;
        end
      3'b100:
        begin
        inc[14]=1'b0 ;
        inc[15]=1'b1 ;
        P_7={(~a_[63]),a_,1'b0} ;
        end
      3'b101:
        begin
        inc[14]=1'b1 ;
        inc[15]=1'b0 ;
        P_7={(~a_[63]),a_[63],a_} ;
        end
      3'b110:
        begin
        inc[14]=1'b1 ;
        inc[15]=1'b0 ;
        P_7={(~a_[63]),a_[63],a_} ;
        end
      3'b011:
        begin
        inc[14]=1'b0 ;
        inc[15]=1'b0 ;
        P_7={(~a[63]),a,1'b0} ;
        end
    endcase

    case({b[17:15]}) // synopsys full_case parallel_case
      3'b000:
        begin
        inc[16]=1'b0 ;
        inc[17]=1'b0 ;
        P_8={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b111:
        begin
        inc[16]=1'b0 ;
        inc[17]=1'b0 ;
        P_8={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b001:
        begin
        inc[16]=1'b0 ;
        inc[17]=1'b0 ;
        P_8={(~a[63]),a[63],a} ;
        end
      3'b010:
        begin
        inc[16]=1'b0 ;
        inc[17]=1'b0 ;
        P_8={(~a[63]),a[63],a} ;
        end
      3'b100:
        begin
        inc[16]=1'b0 ;
        inc[17]=1'b1 ;
        P_8={(~a_[63]),a_,1'b0} ;
        end
      3'b101:
        begin
        inc[16]=1'b1 ;
        inc[17]=1'b0 ;
        P_8={(~a_[63]),a_[63],a_} ;
        end
      3'b110:
        begin
        inc[16]=1'b1 ;
        inc[17]=1'b0 ;
        P_8={(~a_[63]),a_[63],a_} ;
        end
      3'b011:
        begin
        inc[16]=1'b0 ;
        inc[17]=1'b0 ;
        P_8={(~a[63]),a,1'b0} ;
        end
    endcase

    case({b[19:17]}) // synopsys full_case parallel_case
      3'b000:
        begin
        inc[18]=1'b0 ;
        inc[19]=1'b0 ;
        P_9={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b111:
        begin
        inc[18]=1'b0 ;
        inc[19]=1'b0 ;
        P_9={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b001:
        begin
        inc[18]=1'b0 ;
        inc[19]=1'b0 ;
        P_9={(~a[63]),a[63],a} ;
        end
      3'b010:
        begin
        inc[18]=1'b0 ;
        inc[19]=1'b0 ;
        P_9={(~a[63]),a[63],a} ;
        end
      3'b100:
        begin
        inc[18]=1'b0 ;
        inc[19]=1'b1 ;
        P_9={(~a_[63]),a_,1'b0} ;
        end
      3'b101:
        begin
        inc[18]=1'b1 ;
        inc[19]=1'b0 ;
        P_9={(~a_[63]),a_[63],a_} ;
        end
      3'b110:
        begin
        inc[18]=1'b1 ;
        inc[19]=1'b0 ;
        P_9={(~a_[63]),a_[63],a_} ;
        end
      3'b011:
        begin
        inc[18]=1'b0 ;
        inc[19]=1'b0 ;
        P_9={(~a[63]),a,1'b0} ;
        end
    endcase

    case({b[21:19]}) // synopsys full_case parallel_case
      3'b000:
        begin
        inc[20]=1'b0 ;
        inc[21]=1'b0 ;
        P_10={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b111:
        begin
        inc[20]=1'b0 ;
        inc[21]=1'b0 ;
        P_10={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b001:
        begin
        inc[20]=1'b0 ;
        inc[21]=1'b0 ;
        P_10={(~a[63]),a[63],a} ;
        end
      3'b010:
        begin
        inc[20]=1'b0 ;
        inc[21]=1'b0 ;
        P_10={(~a[63]),a[63],a} ;
        end
      3'b100:
        begin
        inc[20]=1'b0 ;
        inc[21]=1'b1 ;
        P_10={(~a_[63]),a_,1'b0} ;
        end
      3'b101:
        begin
        inc[20]=1'b1 ;
        inc[21]=1'b0 ;
        P_10={(~a_[63]),a_[63],a_} ;
        end
      3'b110:
        begin
        inc[20]=1'b1 ;
        inc[21]=1'b0 ;
        P_10={(~a_[63]),a_[63],a_} ;
        end
      3'b011:
        begin
        inc[20]=1'b0 ;
        inc[21]=1'b0 ;
        P_10={(~a[63]),a,1'b0} ;
        end
    endcase

    case({b[23:21]}) // synopsys full_case parallel_case
      3'b000:
        begin
        inc[22]=1'b0 ;
        inc[23]=1'b0 ;
        P_11={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b111:
        begin
        inc[22]=1'b0 ;
        inc[23]=1'b0 ;
        P_11={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b001:
        begin
        inc[22]=1'b0 ;
        inc[23]=1'b0 ;
        P_11={(~a[63]),a[63],a} ;
        end
      3'b010:
        begin
        inc[22]=1'b0 ;
        inc[23]=1'b0 ;
        P_11={(~a[63]),a[63],a} ;
        end
      3'b100:
        begin
        inc[22]=1'b0 ;
        inc[23]=1'b1 ;
        P_11={(~a_[63]),a_,1'b0} ;
        end
      3'b101:
        begin
        inc[22]=1'b1 ;
        inc[23]=1'b0 ;
        P_11={(~a_[63]),a_[63],a_} ;
        end
      3'b110:
        begin
        inc[22]=1'b1 ;
        inc[23]=1'b0 ;
        P_11={(~a_[63]),a_[63],a_} ;
        end
      3'b011:
        begin
        inc[22]=1'b0 ;
        inc[23]=1'b0 ;
        P_11={(~a[63]),a,1'b0} ;
        end
    endcase

    case({b[25:23]}) // synopsys full_case parallel_case
      3'b000:
        begin
        inc[24]=1'b0 ;
        inc[25]=1'b0 ;
        P_12={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b111:
        begin
        inc[24]=1'b0 ;
        inc[25]=1'b0 ;
        P_12={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b001:
        begin
        inc[24]=1'b0 ;
        inc[25]=1'b0 ;
        P_12={(~a[63]),a[63],a} ;
        end
      3'b010:
        begin
        inc[24]=1'b0 ;
        inc[25]=1'b0 ;
        P_12={(~a[63]),a[63],a} ;
        end
      3'b100:
        begin
        inc[24]=1'b0 ;
        inc[25]=1'b1 ;
        P_12={(~a_[63]),a_,1'b0} ;
        end
      3'b101:
        begin
        inc[24]=1'b1 ;
        inc[25]=1'b0 ;
        P_12={(~a_[63]),a_[63],a_} ;
        end
      3'b110:
        begin
        inc[24]=1'b1 ;
        inc[25]=1'b0 ;
        P_12={(~a_[63]),a_[63],a_} ;
        end
      3'b011:
        begin
        inc[24]=1'b0 ;
        inc[25]=1'b0 ;
        P_12={(~a[63]),a,1'b0} ;
        end
    endcase

    case({b[27:25]}) // synopsys full_case parallel_case
      3'b000:
        begin
        inc[26]=1'b0 ;
        inc[27]=1'b0 ;
        P_13={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b111:
        begin
        inc[26]=1'b0 ;
        inc[27]=1'b0 ;
        P_13={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b001:
        begin
        inc[26]=1'b0 ;
        inc[27]=1'b0 ;
        P_13={(~a[63]),a[63],a} ;
        end
      3'b010:
        begin
        inc[26]=1'b0 ;
        inc[27]=1'b0 ;
        P_13={(~a[63]),a[63],a} ;
        end
      3'b100:
        begin
        inc[26]=1'b0 ;
        inc[27]=1'b1 ;
        P_13={(~a_[63]),a_,1'b0} ;
        end
      3'b101:
        begin
        inc[26]=1'b1 ;
        inc[27]=1'b0 ;
        P_13={(~a_[63]),a_[63],a_} ;
        end
      3'b110:
        begin
        inc[26]=1'b1 ;
        inc[27]=1'b0 ;
        P_13={(~a_[63]),a_[63],a_} ;
        end
      3'b011:
        begin
        inc[26]=1'b0 ;
        inc[27]=1'b0 ;
        P_13={(~a[63]),a,1'b0} ;
        end
    endcase

    case({b[29:27]}) // synopsys full_case parallel_case
      3'b000:
        begin
        inc[28]=1'b0 ;
        inc[29]=1'b0 ;
        P_14={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b111:
        begin
        inc[28]=1'b0 ;
        inc[29]=1'b0 ;
        P_14={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b001:
        begin
        inc[28]=1'b0 ;
        inc[29]=1'b0 ;
        P_14={(~a[63]),a[63],a} ;
        end
      3'b010:
        begin
        inc[28]=1'b0 ;
        inc[29]=1'b0 ;
        P_14={(~a[63]),a[63],a} ;
        end
      3'b100:
        begin
        inc[28]=1'b0 ;
        inc[29]=1'b1 ;
        P_14={(~a_[63]),a_,1'b0} ;
        end
      3'b101:
        begin
        inc[28]=1'b1 ;
        inc[29]=1'b0 ;
        P_14={(~a_[63]),a_[63],a_} ;
        end
      3'b110:
        begin
        inc[28]=1'b1 ;
        inc[29]=1'b0 ;
        P_14={(~a_[63]),a_[63],a_} ;
        end
      3'b011:
        begin
        inc[28]=1'b0 ;
        inc[29]=1'b0 ;
        P_14={(~a[63]),a,1'b0} ;
        end
    endcase

    case({b[31:29]}) // synopsys full_case parallel_case
      3'b000:
        begin
        inc[30]=1'b0 ;
        inc[31]=1'b0 ;
        P_15={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b111:
        begin
        inc[30]=1'b0 ;
        inc[31]=1'b0 ;
        P_15={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b001:
        begin
        inc[30]=1'b0 ;
        inc[31]=1'b0 ;
        P_15={(~a[63]),a[63],a} ;
        end
      3'b010:
        begin
        inc[30]=1'b0 ;
        inc[31]=1'b0 ;
        P_15={(~a[63]),a[63],a} ;
        end
      3'b100:
        begin
        inc[30]=1'b0 ;
        inc[31]=1'b1 ;
        P_15={(~a_[63]),a_,1'b0} ;
        end
      3'b101:
        begin
        inc[30]=1'b1 ;
        inc[31]=1'b0 ;
        P_15={(~a_[63]),a_[63],a_} ;
        end
      3'b110:
        begin
        inc[30]=1'b1 ;
        inc[31]=1'b0 ;
        P_15={(~a_[63]),a_[63],a_} ;
        end
      3'b011:
        begin
        inc[30]=1'b0 ;
        inc[31]=1'b0 ;
        P_15={(~a[63]),a,1'b0} ;
        end
    endcase

    case({b[33:31]}) // synopsys full_case parallel_case
      3'b000:
        begin
        inc[32]=1'b0 ;
        inc[33]=1'b0 ;
        P_16={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b111:
        begin
        inc[32]=1'b0 ;
        inc[33]=1'b0 ;
        P_16={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b001:
        begin
        inc[32]=1'b0 ;
        inc[33]=1'b0 ;
        P_16={(~a[63]),a[63],a} ;
        end
      3'b010:
        begin
        inc[32]=1'b0 ;
        inc[33]=1'b0 ;
        P_16={(~a[63]),a[63],a} ;
        end
      3'b100:
        begin
        inc[32]=1'b0 ;
        inc[33]=1'b1 ;
        P_16={(~a_[63]),a_,1'b0} ;
        end
      3'b101:
        begin
        inc[32]=1'b1 ;
        inc[33]=1'b0 ;
        P_16={(~a_[63]),a_[63],a_} ;
        end
      3'b110:
        begin
        inc[32]=1'b1 ;
        inc[33]=1'b0 ;
        P_16={(~a_[63]),a_[63],a_} ;
        end
      3'b011:
        begin
        inc[32]=1'b0 ;
        inc[33]=1'b0 ;
        P_16={(~a[63]),a,1'b0} ;
        end
    endcase

    case({b[35:33]}) // synopsys full_case parallel_case
      3'b000:
        begin
        inc[34]=1'b0 ;
        inc[35]=1'b0 ;
        P_17={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b111:
        begin
        inc[34]=1'b0 ;
        inc[35]=1'b0 ;
        P_17={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b001:
        begin
        inc[34]=1'b0 ;
        inc[35]=1'b0 ;
        P_17={(~a[63]),a[63],a} ;
        end
      3'b010:
        begin
        inc[34]=1'b0 ;
        inc[35]=1'b0 ;
        P_17={(~a[63]),a[63],a} ;
        end
      3'b100:
        begin
        inc[34]=1'b0 ;
        inc[35]=1'b1 ;
        P_17={(~a_[63]),a_,1'b0} ;
        end
      3'b101:
        begin
        inc[34]=1'b1 ;
        inc[35]=1'b0 ;
        P_17={(~a_[63]),a_[63],a_} ;
        end
      3'b110:
        begin
        inc[34]=1'b1 ;
        inc[35]=1'b0 ;
        P_17={(~a_[63]),a_[63],a_} ;
        end
      3'b011:
        begin
        inc[34]=1'b0 ;
        inc[35]=1'b0 ;
        P_17={(~a[63]),a,1'b0} ;
        end
    endcase

    case({b[37:35]}) // synopsys full_case parallel_case
      3'b000:
        begin
        inc[36]=1'b0 ;
        inc[37]=1'b0 ;
        P_18={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b111:
        begin
        inc[36]=1'b0 ;
        inc[37]=1'b0 ;
        P_18={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b001:
        begin
        inc[36]=1'b0 ;
        inc[37]=1'b0 ;
        P_18={(~a[63]),a[63],a} ;
        end
      3'b010:
        begin
        inc[36]=1'b0 ;
        inc[37]=1'b0 ;
        P_18={(~a[63]),a[63],a} ;
        end
      3'b100:
        begin
        inc[36]=1'b0 ;
        inc[37]=1'b1 ;
        P_18={(~a_[63]),a_,1'b0} ;
        end
      3'b101:
        begin
        inc[36]=1'b1 ;
        inc[37]=1'b0 ;
        P_18={(~a_[63]),a_[63],a_} ;
        end
      3'b110:
        begin
        inc[36]=1'b1 ;
        inc[37]=1'b0 ;
        P_18={(~a_[63]),a_[63],a_} ;
        end
      3'b011:
        begin
        inc[36]=1'b0 ;
        inc[37]=1'b0 ;
        P_18={(~a[63]),a,1'b0} ;
        end
    endcase

    case({b[39:37]}) // synopsys full_case parallel_case
      3'b000:
        begin
        inc[38]=1'b0 ;
        inc[39]=1'b0 ;
        P_19={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b111:
        begin
        inc[38]=1'b0 ;
        inc[39]=1'b0 ;
        P_19={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b001:
        begin
        inc[38]=1'b0 ;
        inc[39]=1'b0 ;
        P_19={(~a[63]),a[63],a} ;
        end
      3'b010:
        begin
        inc[38]=1'b0 ;
        inc[39]=1'b0 ;
        P_19={(~a[63]),a[63],a} ;
        end
      3'b100:
        begin
        inc[38]=1'b0 ;
        inc[39]=1'b1 ;
        P_19={(~a_[63]),a_,1'b0} ;
        end
      3'b101:
        begin
        inc[38]=1'b1 ;
        inc[39]=1'b0 ;
        P_19={(~a_[63]),a_[63],a_} ;
        end
      3'b110:
        begin
        inc[38]=1'b1 ;
        inc[39]=1'b0 ;
        P_19={(~a_[63]),a_[63],a_} ;
        end
      3'b011:
        begin
        inc[38]=1'b0 ;
        inc[39]=1'b0 ;
        P_19={(~a[63]),a,1'b0} ;
        end
    endcase

    case({b[41:39]}) // synopsys full_case parallel_case
      3'b000:
        begin
        inc[40]=1'b0 ;
        inc[41]=1'b0 ;
        P_20={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b111:
        begin
        inc[40]=1'b0 ;
        inc[41]=1'b0 ;
        P_20={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b001:
        begin
        inc[40]=1'b0 ;
        inc[41]=1'b0 ;
        P_20={(~a[63]),a[63],a} ;
        end
      3'b010:
        begin
        inc[40]=1'b0 ;
        inc[41]=1'b0 ;
        P_20={(~a[63]),a[63],a} ;
        end
      3'b100:
        begin
        inc[40]=1'b0 ;
        inc[41]=1'b1 ;
        P_20={(~a_[63]),a_,1'b0} ;
        end
      3'b101:
        begin
        inc[40]=1'b1 ;
        inc[41]=1'b0 ;
        P_20={(~a_[63]),a_[63],a_} ;
        end
      3'b110:
        begin
        inc[40]=1'b1 ;
        inc[41]=1'b0 ;
        P_20={(~a_[63]),a_[63],a_} ;
        end
      3'b011:
        begin
        inc[40]=1'b0 ;
        inc[41]=1'b0 ;
        P_20={(~a[63]),a,1'b0} ;
        end
    endcase

    case({b[43:41]}) // synopsys full_case parallel_case
      3'b000:
        begin
        inc[42]=1'b0 ;
        inc[43]=1'b0 ;
        P_21={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b111:
        begin
        inc[42]=1'b0 ;
        inc[43]=1'b0 ;
        P_21={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b001:
        begin
        inc[42]=1'b0 ;
        inc[43]=1'b0 ;
        P_21={(~a[63]),a[63],a} ;
        end
      3'b010:
        begin
        inc[42]=1'b0 ;
        inc[43]=1'b0 ;
        P_21={(~a[63]),a[63],a} ;
        end
      3'b100:
        begin
        inc[42]=1'b0 ;
        inc[43]=1'b1 ;
        P_21={(~a_[63]),a_,1'b0} ;
        end
      3'b101:
        begin
        inc[42]=1'b1 ;
        inc[43]=1'b0 ;
        P_21={(~a_[63]),a_[63],a_} ;
        end
      3'b110:
        begin
        inc[42]=1'b1 ;
        inc[43]=1'b0 ;
        P_21={(~a_[63]),a_[63],a_} ;
        end
      3'b011:
        begin
        inc[42]=1'b0 ;
        inc[43]=1'b0 ;
        P_21={(~a[63]),a,1'b0} ;
        end
    endcase

    case({b[45:43]}) // synopsys full_case parallel_case
      3'b000:
        begin
        inc[44]=1'b0 ;
        inc[45]=1'b0 ;
        P_22={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b111:
        begin
        inc[44]=1'b0 ;
        inc[45]=1'b0 ;
        P_22={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b001:
        begin
        inc[44]=1'b0 ;
        inc[45]=1'b0 ;
        P_22={(~a[63]),a[63],a} ;
        end
      3'b010:
        begin
        inc[44]=1'b0 ;
        inc[45]=1'b0 ;
        P_22={(~a[63]),a[63],a} ;
        end
      3'b100:
        begin
        inc[44]=1'b0 ;
        inc[45]=1'b1 ;
        P_22={(~a_[63]),a_,1'b0} ;
        end
      3'b101:
        begin
        inc[44]=1'b1 ;
        inc[45]=1'b0 ;
        P_22={(~a_[63]),a_[63],a_} ;
        end
      3'b110:
        begin
        inc[44]=1'b1 ;
        inc[45]=1'b0 ;
        P_22={(~a_[63]),a_[63],a_} ;
        end
      3'b011:
        begin
        inc[44]=1'b0 ;
        inc[45]=1'b0 ;
        P_22={(~a[63]),a,1'b0} ;
        end
    endcase

    case({b[47:45]}) // synopsys full_case parallel_case
      3'b000:
        begin
        inc[46]=1'b0 ;
        inc[47]=1'b0 ;
        P_23={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b111:
        begin
        inc[46]=1'b0 ;
        inc[47]=1'b0 ;
        P_23={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b001:
        begin
        inc[46]=1'b0 ;
        inc[47]=1'b0 ;
        P_23={(~a[63]),a[63],a} ;
        end
      3'b010:
        begin
        inc[46]=1'b0 ;
        inc[47]=1'b0 ;
        P_23={(~a[63]),a[63],a} ;
        end
      3'b100:
        begin
        inc[46]=1'b0 ;
        inc[47]=1'b1 ;
        P_23={(~a_[63]),a_,1'b0} ;
        end
      3'b101:
        begin
        inc[46]=1'b1 ;
        inc[47]=1'b0 ;
        P_23={(~a_[63]),a_[63],a_} ;
        end
      3'b110:
        begin
        inc[46]=1'b1 ;
        inc[47]=1'b0 ;
        P_23={(~a_[63]),a_[63],a_} ;
        end
      3'b011:
        begin
        inc[46]=1'b0 ;
        inc[47]=1'b0 ;
        P_23={(~a[63]),a,1'b0} ;
        end
    endcase

    case({b[49:47]}) // synopsys full_case parallel_case
      3'b000:
        begin
        inc[48]=1'b0 ;
        inc[49]=1'b0 ;
        P_24={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b111:
        begin
        inc[48]=1'b0 ;
        inc[49]=1'b0 ;
        P_24={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b001:
        begin
        inc[48]=1'b0 ;
        inc[49]=1'b0 ;
        P_24={(~a[63]),a[63],a} ;
        end
      3'b010:
        begin
        inc[48]=1'b0 ;
        inc[49]=1'b0 ;
        P_24={(~a[63]),a[63],a} ;
        end
      3'b100:
        begin
        inc[48]=1'b0 ;
        inc[49]=1'b1 ;
        P_24={(~a_[63]),a_,1'b0} ;
        end
      3'b101:
        begin
        inc[48]=1'b1 ;
        inc[49]=1'b0 ;
        P_24={(~a_[63]),a_[63],a_} ;
        end
      3'b110:
        begin
        inc[48]=1'b1 ;
        inc[49]=1'b0 ;
        P_24={(~a_[63]),a_[63],a_} ;
        end
      3'b011:
        begin
        inc[48]=1'b0 ;
        inc[49]=1'b0 ;
        P_24={(~a[63]),a,1'b0} ;
        end
    endcase

    case({b[51:49]}) // synopsys full_case parallel_case
      3'b000:
        begin
        inc[50]=1'b0 ;
        inc[51]=1'b0 ;
        P_25={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b111:
        begin
        inc[50]=1'b0 ;
        inc[51]=1'b0 ;
        P_25={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b001:
        begin
        inc[50]=1'b0 ;
        inc[51]=1'b0 ;
        P_25={(~a[63]),a[63],a} ;
        end
      3'b010:
        begin
        inc[50]=1'b0 ;
        inc[51]=1'b0 ;
        P_25={(~a[63]),a[63],a} ;
        end
      3'b100:
        begin
        inc[50]=1'b0 ;
        inc[51]=1'b1 ;
        P_25={(~a_[63]),a_,1'b0} ;
        end
      3'b101:
        begin
        inc[50]=1'b1 ;
        inc[51]=1'b0 ;
        P_25={(~a_[63]),a_[63],a_} ;
        end
      3'b110:
        begin
        inc[50]=1'b1 ;
        inc[51]=1'b0 ;
        P_25={(~a_[63]),a_[63],a_} ;
        end
      3'b011:
        begin
        inc[50]=1'b0 ;
        inc[51]=1'b0 ;
        P_25={(~a[63]),a,1'b0} ;
        end
    endcase

    case({b[53:51]}) // synopsys full_case parallel_case
      3'b000:
        begin
        inc[52]=1'b0 ;
        inc[53]=1'b0 ;
        P_26={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b111:
        begin
        inc[52]=1'b0 ;
        inc[53]=1'b0 ;
        P_26={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b001:
        begin
        inc[52]=1'b0 ;
        inc[53]=1'b0 ;
        P_26={(~a[63]),a[63],a} ;
        end
      3'b010:
        begin
        inc[52]=1'b0 ;
        inc[53]=1'b0 ;
        P_26={(~a[63]),a[63],a} ;
        end
      3'b100:
        begin
        inc[52]=1'b0 ;
        inc[53]=1'b1 ;
        P_26={(~a_[63]),a_,1'b0} ;
        end
      3'b101:
        begin
        inc[52]=1'b1 ;
        inc[53]=1'b0 ;
        P_26={(~a_[63]),a_[63],a_} ;
        end
      3'b110:
        begin
        inc[52]=1'b1 ;
        inc[53]=1'b0 ;
        P_26={(~a_[63]),a_[63],a_} ;
        end
      3'b011:
        begin
        inc[52]=1'b0 ;
        inc[53]=1'b0 ;
        P_26={(~a[63]),a,1'b0} ;
        end
    endcase

    case({b[55:53]}) // synopsys full_case parallel_case
      3'b000:
        begin
        inc[54]=1'b0 ;
        inc[55]=1'b0 ;
        P_27={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b111:
        begin
        inc[54]=1'b0 ;
        inc[55]=1'b0 ;
        P_27={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b001:
        begin
        inc[54]=1'b0 ;
        inc[55]=1'b0 ;
        P_27={(~a[63]),a[63],a} ;
        end
      3'b010:
        begin
        inc[54]=1'b0 ;
        inc[55]=1'b0 ;
        P_27={(~a[63]),a[63],a} ;
        end
      3'b100:
        begin
        inc[54]=1'b0 ;
        inc[55]=1'b1 ;
        P_27={(~a_[63]),a_,1'b0} ;
        end
      3'b101:
        begin
        inc[54]=1'b1 ;
        inc[55]=1'b0 ;
        P_27={(~a_[63]),a_[63],a_} ;
        end
      3'b110:
        begin
        inc[54]=1'b1 ;
        inc[55]=1'b0 ;
        P_27={(~a_[63]),a_[63],a_} ;
        end
      3'b011:
        begin
        inc[54]=1'b0 ;
        inc[55]=1'b0 ;
        P_27={(~a[63]),a,1'b0} ;
        end
    endcase

    case({b[57:55]}) // synopsys full_case parallel_case
      3'b000:
        begin
        inc[56]=1'b0 ;
        inc[57]=1'b0 ;
        P_28={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b111:
        begin
        inc[56]=1'b0 ;
        inc[57]=1'b0 ;
        P_28={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b001:
        begin
        inc[56]=1'b0 ;
        inc[57]=1'b0 ;
        P_28={(~a[63]),a[63],a} ;
        end
      3'b010:
        begin
        inc[56]=1'b0 ;
        inc[57]=1'b0 ;
        P_28={(~a[63]),a[63],a} ;
        end
      3'b100:
        begin
        inc[56]=1'b0 ;
        inc[57]=1'b1 ;
        P_28={(~a_[63]),a_,1'b0} ;
        end
      3'b101:
        begin
        inc[56]=1'b1 ;
        inc[57]=1'b0 ;
        P_28={(~a_[63]),a_[63],a_} ;
        end
      3'b110:
        begin
        inc[56]=1'b1 ;
        inc[57]=1'b0 ;
        P_28={(~a_[63]),a_[63],a_} ;
        end
      3'b011:
        begin
        inc[56]=1'b0 ;
        inc[57]=1'b0 ;
        P_28={(~a[63]),a,1'b0} ;
        end
    endcase

    case({b[59:57]}) // synopsys full_case parallel_case
      3'b000:
        begin
        inc[58]=1'b0 ;
        inc[59]=1'b0 ;
        P_29={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b111:
        begin
        inc[58]=1'b0 ;
        inc[59]=1'b0 ;
        P_29={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b001:
        begin
        inc[58]=1'b0 ;
        inc[59]=1'b0 ;
        P_29={(~a[63]),a[63],a} ;
        end
      3'b010:
        begin
        inc[58]=1'b0 ;
        inc[59]=1'b0 ;
        P_29={(~a[63]),a[63],a} ;
        end
      3'b100:
        begin
        inc[58]=1'b0 ;
        inc[59]=1'b1 ;
        P_29={(~a_[63]),a_,1'b0} ;
        end
      3'b101:
        begin
        inc[58]=1'b1 ;
        inc[59]=1'b0 ;
        P_29={(~a_[63]),a_[63],a_} ;
        end
      3'b110:
        begin
        inc[58]=1'b1 ;
        inc[59]=1'b0 ;
        P_29={(~a_[63]),a_[63],a_} ;
        end
      3'b011:
        begin
        inc[58]=1'b0 ;
        inc[59]=1'b0 ;
        P_29={(~a[63]),a,1'b0} ;
        end
    endcase

    case({b[61:59]}) // synopsys full_case parallel_case
      3'b000:
        begin
        inc[60]=1'b0 ;
        inc[61]=1'b0 ;
        P_30={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b111:
        begin
        inc[60]=1'b0 ;
        inc[61]=1'b0 ;
        P_30={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b001:
        begin
        inc[60]=1'b0 ;
        inc[61]=1'b0 ;
        P_30={(~a[63]),a[63],a} ;
        end
      3'b010:
        begin
        inc[60]=1'b0 ;
        inc[61]=1'b0 ;
        P_30={(~a[63]),a[63],a} ;
        end
      3'b100:
        begin
        inc[60]=1'b0 ;
        inc[61]=1'b1 ;
        P_30={(~a_[63]),a_,1'b0} ;
        end
      3'b101:
        begin
        inc[60]=1'b1 ;
        inc[61]=1'b0 ;
        P_30={(~a_[63]),a_[63],a_} ;
        end
      3'b110:
        begin
        inc[60]=1'b1 ;
        inc[61]=1'b0 ;
        P_30={(~a_[63]),a_[63],a_} ;
        end
      3'b011:
        begin
        inc[60]=1'b0 ;
        inc[61]=1'b0 ;
        P_30={(~a[63]),a,1'b0} ;
        end
    endcase

    case({b[63:61]}) // synopsys full_case parallel_case
      3'b000:
        begin
        inc[62]=1'b0 ;
        inc[63]=1'b0 ;
        P_31={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b111:
        begin
        inc[62]=1'b0 ;
        inc[63]=1'b0 ;
        P_31={1'b1,{65'b00000000000000000000000000000000000000000000000000000000000000000}} ;
        end
      3'b001:
        begin
        inc[62]=1'b0 ;
        inc[63]=1'b0 ;
        P_31={(~a[63]),a[63],a} ;
        end
      3'b010:
        begin
        inc[62]=1'b0 ;
        inc[63]=1'b0 ;
        P_31={(~a[63]),a[63],a} ;
        end
      3'b100:
        begin
        inc[62]=1'b0 ;
        inc[63]=1'b1 ;
        P_31={(~a_[63]),a_,1'b0} ;
        end
      3'b101:
        begin
        inc[62]=1'b1 ;
        inc[63]=1'b0 ;
        P_31={(~a_[63]),a_[63],a_} ;
        end
      3'b110:
        begin
        inc[62]=1'b1 ;
        inc[63]=1'b0 ;
        P_31={(~a_[63]),a_[63],a_} ;
        end
      3'b011:
        begin
        inc[62]=1'b0 ;
        inc[63]=1'b0 ;
        P_31={(~a[63]),a,1'b0} ;
        end
    endcase

    end


  // ***** Bit 0 ***** //
  Hadder_ A_0_0( .carry(c[0]), .sum(s[0]), .in2(inc[0]), .in1(P_0[0]) );

  // ***** Bit 1 ***** //
  Hadder_ A_1_1( .carry(c[1]), .sum(s[1]), .in2(inc[1]), .in1(P_0[1]) );

  // ***** Bit 2 ***** //
  Fadder_ A_2_2( .carry(c[2]), .sum(s[2]), .in3(inc[2]), .in2(P_1[0]), .in1(P_0[2]) );

  // ***** Bit 3 ***** //
  Fadder_ A_3_3( .carry(c[3]), .sum(s[3]), .in3(inc[3]), .in2(P_1[1]), .in1(P_0[3]) );

  // ***** Bit 4 ***** //
  Hadder_ A_4_4( .carry(c_4_4), .sum(s_4_4), .in2(inc[4]), .in1(P_2[0]) );
  Fadder_ A_4_5( .carry(c[4]), .sum(s[4]), .in3(P_1[2]), .in2(P_0[4]), .in1(s_4_4) );

  // ***** Bit 5 ***** //
  Fadder_ A_5_6( .carry(c_5_6), .sum(s_5_6), .in3(inc[5]), .in2(P_2[1]), .in1(P_1[3]) );
  Fadder_ A_5_7( .carry(c[5]), .sum(s[5]), .in3(P_0[5]), .in2(c_4_4), .in1(s_5_6) );

  // ***** Bit 6 ***** //
  Hadder_ A_6_8( .carry(c_6_8), .sum(s_6_8), .in2(inc[6]), .in1(P_3[0]) );
  Fadder_ A_6_9( .carry(c_6_9), .sum(s_6_9), .in3(P_2[2]), .in2(P_1[4]), .in1(P_0[6]) );
  Fadder_ A_6_10( .carry(c[6]), .sum(s[6]), .in3(c_5_6), .in2(s_6_8), .in1(s_6_9) );

  // ***** Bit 7 ***** //
  Fadder_ A_7_11( .carry(c_7_11), .sum(s_7_11), .in3(inc[7]), .in2(P_3[1]), .in1(P_2[3]) );
  Fadder_ A_7_12( .carry(c_7_12), .sum(s_7_12), .in3(P_1[5]), .in2(P_0[7]), .in1(c_6_8) );
  Fadder_ A_7_13( .carry(c[7]), .sum(s[7]), .in3(c_6_9), .in2(s_7_11), .in1(s_7_12) );

  // ***** Bit 8 ***** //
  Hadder_ A_8_14( .carry(c_8_14), .sum(s_8_14), .in2(inc[8]), .in1(P_4[0]) );
  Fadder_ A_8_15( .carry(c_8_15), .sum(s_8_15), .in3(P_3[2]), .in2(P_2[4]), .in1(P_1[6]) );
  Fadder_ A_8_16( .carry(c_8_16), .sum(s_8_16), .in3(P_0[8]), .in2(c_7_11), .in1(s_8_14) );
  Fadder_ A_8_17( .carry(c[8]), .sum(s[8]), .in3(s_8_15), .in2(c_7_12), .in1(s_8_16) );

  // ***** Bit 9 ***** //
  Fadder_ A_9_18( .carry(c_9_18), .sum(s_9_18), .in3(inc[9]), .in2(P_4[1]), .in1(P_3[3]) );
  Fadder_ A_9_19( .carry(c_9_19), .sum(s_9_19), .in3(P_2[5]), .in2(P_1[7]), .in1(P_0[9]) );
  Fadder_ A_9_20( .carry(c_9_20), .sum(s_9_20), .in3(c_8_14), .in2(c_8_15), .in1(s_9_19) );
  Fadder_ A_9_21( .carry(c[9]), .sum(s[9]), .in3(s_9_18), .in2(c_8_16), .in1(s_9_20) );

  // ***** Bit 10 ***** //
  Hadder_ A_10_22( .carry(c_10_22), .sum(s_10_22), .in2(inc[10]), .in1(P_5[0]) );
  Fadder_ A_10_23( .carry(c_10_23), .sum(s_10_23), .in3(P_4[2]), .in2(P_3[4]), .in1(P_2[6]) );
  Fadder_ A_10_24( .carry(c_10_24), .sum(s_10_24), .in3(P_1[8]), .in2(P_0[10]), .in1(c_9_19) );
  Fadder_ A_10_25( .carry(c_10_25), .sum(s_10_25), .in3(c_9_18), .in2(s_10_22), .in1(s_10_23) );
  Fadder_ A_10_26( .carry(c[10]), .sum(s[10]), .in3(c_9_20), .in2(s_10_24), .in1(s_10_25) );

  // ***** Bit 11 ***** //
  Fadder_ A_11_27( .carry(c_11_27), .sum(s_11_27), .in3(inc[11]), .in2(P_5[1]), .in1(P_4[3]) );
  Fadder_ A_11_28( .carry(c_11_28), .sum(s_11_28), .in3(P_3[5]), .in2(P_2[7]), .in1(P_1[9]) );
  Fadder_ A_11_29( .carry(c_11_29), .sum(s_11_29), .in3(P_0[11]), .in2(c_10_22), .in1(c_10_23) );
  Fadder_ A_11_30( .carry(c_11_30), .sum(s_11_30), .in3(s_11_28), .in2(s_11_27), .in1(c_10_24) );
  Fadder_ A_11_31( .carry(c[11]), .sum(s[11]), .in3(s_11_29), .in2(c_10_25), .in1(s_11_30) );

  // ***** Bit 12 ***** //
  Hadder_ A_12_32( .carry(c_12_32), .sum(s_12_32), .in2(inc[12]), .in1(P_6[0]) );
  Fadder_ A_12_33( .carry(c_12_33), .sum(s_12_33), .in3(P_5[2]), .in2(P_4[4]), .in1(P_3[6]) );
  Fadder_ A_12_34( .carry(c_12_34), .sum(s_12_34), .in3(P_2[8]), .in2(P_1[10]), .in1(P_0[12]) );
  Fadder_ A_12_35( .carry(c_12_35), .sum(s_12_35), .in3(c_11_28), .in2(c_11_27), .in1(s_12_32) );
  Fadder_ A_12_36( .carry(c_12_36), .sum(s_12_36), .in3(s_12_34), .in2(s_12_33), .in1(c_11_29) );
  Fadder_ A_12_37( .carry(c[12]), .sum(s[12]), .in3(s_12_35), .in2(c_11_30), .in1(s_12_36) );

  // ***** Bit 13 ***** //
  Fadder_ A_13_38( .carry(c_13_38), .sum(s_13_38), .in3(inc[13]), .in2(P_6[1]), .in1(P_5[3]) );
  Fadder_ A_13_39( .carry(c_13_39), .sum(s_13_39), .in3(P_4[5]), .in2(P_3[7]), .in1(P_2[9]) );
  Fadder_ A_13_40( .carry(c_13_40), .sum(s_13_40), .in3(P_1[11]), .in2(P_0[13]), .in1(c_12_32) );
  Fadder_ A_13_41( .carry(c_13_41), .sum(s_13_41), .in3(c_12_34), .in2(c_12_33), .in1(s_13_39) );
  Fadder_ A_13_42( .carry(c_13_42), .sum(s_13_42), .in3(s_13_38), .in2(s_13_40), .in1(c_12_35) );
  Fadder_ A_13_43( .carry(c[13]), .sum(s[13]), .in3(s_13_41), .in2(c_12_36), .in1(s_13_42) );

  // ***** Bit 14 ***** //
  Hadder_ A_14_44( .carry(c_14_44), .sum(s_14_44), .in2(inc[14]), .in1(P_7[0]) );
  Fadder_ A_14_45( .carry(c_14_45), .sum(s_14_45), .in3(P_6[2]), .in2(P_5[4]), .in1(P_4[6]) );
  Fadder_ A_14_46( .carry(c_14_46), .sum(s_14_46), .in3(P_3[8]), .in2(P_2[10]), .in1(P_1[12]) );
  Fadder_ A_14_47( .carry(c_14_47), .sum(s_14_47), .in3(P_0[14]), .in2(c_13_39), .in1(c_13_38) );
  Fadder_ A_14_48( .carry(c_14_48), .sum(s_14_48), .in3(s_14_44), .in2(s_14_46), .in1(s_14_45) );
  Fadder_ A_14_49( .carry(c_14_49), .sum(s_14_49), .in3(c_13_40), .in2(c_13_41), .in1(s_14_47) );
  Fadder_ A_14_50( .carry(c[14]), .sum(s[14]), .in3(s_14_48), .in2(c_13_42), .in1(s_14_49) );

  // ***** Bit 15 ***** //
  Fadder_ A_15_51( .carry(c_15_51), .sum(s_15_51), .in3(inc[15]), .in2(P_7[1]), .in1(P_6[3]) );
  Fadder_ A_15_52( .carry(c_15_52), .sum(s_15_52), .in3(P_5[5]), .in2(P_4[7]), .in1(P_3[9]) );
  Fadder_ A_15_53( .carry(c_15_53), .sum(s_15_53), .in3(P_2[11]), .in2(P_1[13]), .in1(P_0[15]) );
  Fadder_ A_15_54( .carry(c_15_54), .sum(s_15_54), .in3(c_14_44), .in2(c_14_46), .in1(c_14_45) );
  Fadder_ A_15_55( .carry(c_15_55), .sum(s_15_55), .in3(s_15_53), .in2(s_15_52), .in1(s_15_51) );
  Fadder_ A_15_56( .carry(c_15_56), .sum(s_15_56), .in3(c_14_47), .in2(s_15_54), .in1(c_14_48) );
  Fadder_ A_15_57( .carry(c[15]), .sum(s[15]), .in3(s_15_55), .in2(c_14_49), .in1(s_15_56) );

  // ***** Bit 16 ***** //
  Hadder_ A_16_58( .carry(c_16_58), .sum(s_16_58), .in2(inc[16]), .in1(P_8[0]) );
  Fadder_ A_16_59( .carry(c_16_59), .sum(s_16_59), .in3(P_7[2]), .in2(P_6[4]), .in1(P_5[6]) );
  Fadder_ A_16_60( .carry(c_16_60), .sum(s_16_60), .in3(P_4[8]), .in2(P_3[10]), .in1(P_2[12]) );
  Fadder_ A_16_61( .carry(c_16_61), .sum(s_16_61), .in3(P_1[14]), .in2(P_0[16]), .in1(c_15_53) );
  Fadder_ A_16_62( .carry(c_16_62), .sum(s_16_62), .in3(c_15_52), .in2(c_15_51), .in1(s_16_58) );
  Fadder_ A_16_63( .carry(c_16_63), .sum(s_16_63), .in3(s_16_60), .in2(s_16_59), .in1(c_15_54) );
  Fadder_ A_16_64( .carry(c_16_64), .sum(s_16_64), .in3(s_16_61), .in2(c_15_55), .in1(s_16_62) );
  Fadder_ A_16_65( .carry(c[16]), .sum(s[16]), .in3(s_16_63), .in2(c_15_56), .in1(s_16_64) );

  // ***** Bit 17 ***** //
  Fadder_ A_17_66( .carry(c_17_66), .sum(s_17_66), .in3(inc[17]), .in2(P_8[1]), .in1(P_7[3]) );
  Fadder_ A_17_67( .carry(c_17_67), .sum(s_17_67), .in3(P_6[5]), .in2(P_5[7]), .in1(P_4[9]) );
  Fadder_ A_17_68( .carry(c_17_68), .sum(s_17_68), .in3(P_3[11]), .in2(P_2[13]), .in1(P_1[15]) );
  Fadder_ A_17_69( .carry(c_17_69), .sum(s_17_69), .in3(P_0[17]), .in2(c_16_58), .in1(c_16_60) );
  Fadder_ A_17_70( .carry(c_17_70), .sum(s_17_70), .in3(c_16_59), .in2(s_17_68), .in1(s_17_67) );
  Fadder_ A_17_71( .carry(c_17_71), .sum(s_17_71), .in3(s_17_66), .in2(c_16_61), .in1(c_16_62) );
  Fadder_ A_17_72( .carry(c_17_72), .sum(s_17_72), .in3(s_17_69), .in2(s_17_70), .in1(c_16_63) );
  Fadder_ A_17_73( .carry(c[17]), .sum(s[17]), .in3(s_17_71), .in2(c_16_64), .in1(s_17_72) );

  // ***** Bit 18 ***** //
  Hadder_ A_18_74( .carry(c_18_74), .sum(s_18_74), .in2(inc[18]), .in1(P_9[0]) );
  Fadder_ A_18_75( .carry(c_18_75), .sum(s_18_75), .in3(P_8[2]), .in2(P_7[4]), .in1(P_6[6]) );
  Fadder_ A_18_76( .carry(c_18_76), .sum(s_18_76), .in3(P_5[8]), .in2(P_4[10]), .in1(P_3[12]) );
  Fadder_ A_18_77( .carry(c_18_77), .sum(s_18_77), .in3(P_2[14]), .in2(P_1[16]), .in1(P_0[18]) );
  Fadder_ A_18_78( .carry(c_18_78), .sum(s_18_78), .in3(c_17_68), .in2(c_17_67), .in1(c_17_66) );
  Fadder_ A_18_79( .carry(c_18_79), .sum(s_18_79), .in3(s_18_74), .in2(s_18_77), .in1(s_18_76) );
  Fadder_ A_18_80( .carry(c_18_80), .sum(s_18_80), .in3(s_18_75), .in2(c_17_69), .in1(s_18_78) );
  Fadder_ A_18_81( .carry(c_18_81), .sum(s_18_81), .in3(c_17_70), .in2(s_18_79), .in1(c_17_71) );
  Fadder_ A_18_82( .carry(c[18]), .sum(s[18]), .in3(s_18_80), .in2(c_17_72), .in1(s_18_81) );

  // ***** Bit 19 ***** //
  Fadder_ A_19_83( .carry(c_19_83), .sum(s_19_83), .in3(inc[19]), .in2(P_9[1]), .in1(P_8[3]) );
  Fadder_ A_19_84( .carry(c_19_84), .sum(s_19_84), .in3(P_7[5]), .in2(P_6[7]), .in1(P_5[9]) );
  Fadder_ A_19_85( .carry(c_19_85), .sum(s_19_85), .in3(P_4[11]), .in2(P_3[13]), .in1(P_2[15]) );
  Fadder_ A_19_86( .carry(c_19_86), .sum(s_19_86), .in3(P_1[17]), .in2(P_0[19]), .in1(c_18_74) );
  Fadder_ A_19_87( .carry(c_19_87), .sum(s_19_87), .in3(c_18_77), .in2(c_18_76), .in1(c_18_75) );
  Fadder_ A_19_88( .carry(c_19_88), .sum(s_19_88), .in3(s_19_85), .in2(s_19_84), .in1(s_19_83) );
  Fadder_ A_19_89( .carry(c_19_89), .sum(s_19_89), .in3(s_19_86), .in2(c_18_78), .in1(s_19_87) );
  Fadder_ A_19_90( .carry(c_19_90), .sum(s_19_90), .in3(c_18_79), .in2(s_19_88), .in1(c_18_80) );
  Fadder_ A_19_91( .carry(c[19]), .sum(s[19]), .in3(s_19_89), .in2(c_18_81), .in1(s_19_90) );

  // ***** Bit 20 ***** //
  Hadder_ A_20_92( .carry(c_20_92), .sum(s_20_92), .in2(inc[20]), .in1(P_10[0]) );
  Fadder_ A_20_93( .carry(c_20_93), .sum(s_20_93), .in3(P_9[2]), .in2(P_8[4]), .in1(P_7[6]) );
  Fadder_ A_20_94( .carry(c_20_94), .sum(s_20_94), .in3(P_6[8]), .in2(P_5[10]), .in1(P_4[12]) );
  Fadder_ A_20_95( .carry(c_20_95), .sum(s_20_95), .in3(P_3[14]), .in2(P_2[16]), .in1(P_1[18]) );
  Fadder_ A_20_96( .carry(c_20_96), .sum(s_20_96), .in3(P_0[20]), .in2(c_19_85), .in1(c_19_84) );
  Fadder_ A_20_97( .carry(c_20_97), .sum(s_20_97), .in3(c_19_83), .in2(s_20_92), .in1(s_20_95) );
  Fadder_ A_20_98( .carry(c_20_98), .sum(s_20_98), .in3(s_20_94), .in2(s_20_93), .in1(c_19_86) );
  Fadder_ A_20_99( .carry(c_20_99), .sum(s_20_99), .in3(c_19_87), .in2(s_20_96), .in1(c_19_88) );
  Fadder_ A_20_100( .carry(c_20_100), .sum(s_20_100), .in3(s_20_97), .in2(s_20_98), .in1(c_19_89) );
  Fadder_ A_20_101( .carry(c[20]), .sum(s[20]), .in3(s_20_99), .in2(c_19_90), .in1(s_20_100) );

  // ***** Bit 21 ***** //
  Fadder_ A_21_102( .carry(c_21_102), .sum(s_21_102), .in3(inc[21]), .in2(P_10[1]), .in1(P_9[3]) );
  Fadder_ A_21_103( .carry(c_21_103), .sum(s_21_103), .in3(P_8[5]), .in2(P_7[7]), .in1(P_6[9]) );
  Fadder_ A_21_104( .carry(c_21_104), .sum(s_21_104), .in3(P_5[11]), .in2(P_4[13]), .in1(P_3[15]) );
  Fadder_ A_21_105( .carry(c_21_105), .sum(s_21_105), .in3(P_2[17]), .in2(P_1[19]), .in1(P_0[21]) );
  Fadder_ A_21_106( .carry(c_21_106), .sum(s_21_106), .in3(c_20_92), .in2(c_20_95), .in1(c_20_94) );
  Fadder_ A_21_107( .carry(c_21_107), .sum(s_21_107), .in3(c_20_93), .in2(s_21_105), .in1(s_21_104) );
  Fadder_ A_21_108( .carry(c_21_108), .sum(s_21_108), .in3(s_21_103), .in2(s_21_102), .in1(c_20_96) );
  Fadder_ A_21_109( .carry(c_21_109), .sum(s_21_109), .in3(s_21_106), .in2(c_20_97), .in1(c_20_98) );
  Fadder_ A_21_110( .carry(c_21_110), .sum(s_21_110), .in3(s_21_107), .in2(s_21_108), .in1(c_20_99) );
  Fadder_ A_21_111( .carry(c[21]), .sum(s[21]), .in3(s_21_109), .in2(c_20_100), .in1(s_21_110) );

  // ***** Bit 22 ***** //
  Hadder_ A_22_112( .carry(c_22_112), .sum(s_22_112), .in2(inc[22]), .in1(P_11[0]) );
  Fadder_ A_22_113( .carry(c_22_113), .sum(s_22_113), .in3(P_10[2]), .in2(P_9[4]), .in1(P_8[6]) );
  Fadder_ A_22_114( .carry(c_22_114), .sum(s_22_114), .in3(P_7[8]), .in2(P_6[10]), .in1(P_5[12]) );
  Fadder_ A_22_115( .carry(c_22_115), .sum(s_22_115), .in3(P_4[14]), .in2(P_3[16]), .in1(P_2[18]) );
  Fadder_ A_22_116( .carry(c_22_116), .sum(s_22_116), .in3(P_1[20]), .in2(P_0[22]), .in1(c_21_105) );
  Fadder_ A_22_117( .carry(c_22_117), .sum(s_22_117), .in3(c_21_104), .in2(c_21_103), .in1(c_21_102) );
  Fadder_ A_22_118( .carry(c_22_118), .sum(s_22_118), .in3(s_22_112), .in2(s_22_115), .in1(s_22_114) );
  Fadder_ A_22_119( .carry(c_22_119), .sum(s_22_119), .in3(s_22_113), .in2(c_21_106), .in1(s_22_116) );
  Fadder_ A_22_120( .carry(c_22_120), .sum(s_22_120), .in3(s_22_117), .in2(c_21_107), .in1(s_22_118) );
  Fadder_ A_22_121( .carry(c_22_121), .sum(s_22_121), .in3(c_21_108), .in2(c_21_109), .in1(s_22_119) );
  Fadder_ A_22_122( .carry(c[22]), .sum(s[22]), .in3(s_22_120), .in2(c_21_110), .in1(s_22_121) );

  // ***** Bit 23 ***** //
  Fadder_ A_23_123( .carry(c_23_123), .sum(s_23_123), .in3(inc[23]), .in2(P_11[1]), .in1(P_10[3]) );
  Fadder_ A_23_124( .carry(c_23_124), .sum(s_23_124), .in3(P_9[5]), .in2(P_8[7]), .in1(P_7[9]) );
  Fadder_ A_23_125( .carry(c_23_125), .sum(s_23_125), .in3(P_6[11]), .in2(P_5[13]), .in1(P_4[15]) );
  Fadder_ A_23_126( .carry(c_23_126), .sum(s_23_126), .in3(P_3[17]), .in2(P_2[19]), .in1(P_1[21]) );
  Fadder_ A_23_127( .carry(c_23_127), .sum(s_23_127), .in3(P_0[23]), .in2(c_22_112), .in1(c_22_115) );
  Fadder_ A_23_128( .carry(c_23_128), .sum(s_23_128), .in3(c_22_114), .in2(c_22_113), .in1(s_23_126) );
  Fadder_ A_23_129( .carry(c_23_129), .sum(s_23_129), .in3(s_23_125), .in2(s_23_124), .in1(s_23_123) );
  Fadder_ A_23_130( .carry(c_23_130), .sum(s_23_130), .in3(c_22_116), .in2(c_22_117), .in1(s_23_127) );
  Fadder_ A_23_131( .carry(c_23_131), .sum(s_23_131), .in3(c_22_118), .in2(s_23_128), .in1(s_23_129) );
  Fadder_ A_23_132( .carry(c_23_132), .sum(s_23_132), .in3(c_22_119), .in2(c_22_120), .in1(s_23_130) );
  Fadder_ A_23_133( .carry(c[23]), .sum(s[23]), .in3(s_23_131), .in2(c_22_121), .in1(s_23_132) );

  // ***** Bit 24 ***** //
  Hadder_ A_24_134( .carry(c_24_134), .sum(s_24_134), .in2(inc[24]), .in1(P_12[0]) );
  Fadder_ A_24_135( .carry(c_24_135), .sum(s_24_135), .in3(P_11[2]), .in2(P_10[4]), .in1(P_9[6]) );
  Fadder_ A_24_136( .carry(c_24_136), .sum(s_24_136), .in3(P_8[8]), .in2(P_7[10]), .in1(P_6[12]) );
  Fadder_ A_24_137( .carry(c_24_137), .sum(s_24_137), .in3(P_5[14]), .in2(P_4[16]), .in1(P_3[18]) );
  Fadder_ A_24_138( .carry(c_24_138), .sum(s_24_138), .in3(P_2[20]), .in2(P_1[22]), .in1(P_0[24]) );
  Fadder_ A_24_139( .carry(c_24_139), .sum(s_24_139), .in3(c_23_126), .in2(c_23_125), .in1(c_23_124) );
  Fadder_ A_24_140( .carry(c_24_140), .sum(s_24_140), .in3(c_23_123), .in2(s_24_134), .in1(s_24_138) );
  Fadder_ A_24_141( .carry(c_24_141), .sum(s_24_141), .in3(s_24_137), .in2(s_24_136), .in1(s_24_135) );
  Fadder_ A_24_142( .carry(c_24_142), .sum(s_24_142), .in3(c_23_127), .in2(c_23_128), .in1(s_24_139) );
  Fadder_ A_24_143( .carry(c_24_143), .sum(s_24_143), .in3(c_23_129), .in2(s_24_140), .in1(s_24_141) );
  Fadder_ A_24_144( .carry(c_24_144), .sum(s_24_144), .in3(c_23_130), .in2(s_24_142), .in1(c_23_131) );
  Fadder_ A_24_145( .carry(c[24]), .sum(s[24]), .in3(s_24_143), .in2(c_23_132), .in1(s_24_144) );

  // ***** Bit 25 ***** //
  Fadder_ A_25_146( .carry(c_25_146), .sum(s_25_146), .in3(inc[25]), .in2(P_12[1]), .in1(P_11[3]) );
  Fadder_ A_25_147( .carry(c_25_147), .sum(s_25_147), .in3(P_10[5]), .in2(P_9[7]), .in1(P_8[9]) );
  Fadder_ A_25_148( .carry(c_25_148), .sum(s_25_148), .in3(P_7[11]), .in2(P_6[13]), .in1(P_5[15]) );
  Fadder_ A_25_149( .carry(c_25_149), .sum(s_25_149), .in3(P_4[17]), .in2(P_3[19]), .in1(P_2[21]) );
  Fadder_ A_25_150( .carry(c_25_150), .sum(s_25_150), .in3(P_1[23]), .in2(P_0[25]), .in1(c_24_134) );
  Fadder_ A_25_151( .carry(c_25_151), .sum(s_25_151), .in3(c_24_138), .in2(c_24_137), .in1(c_24_136) );
  Fadder_ A_25_152( .carry(c_25_152), .sum(s_25_152), .in3(c_24_135), .in2(s_25_149), .in1(s_25_148) );
  Fadder_ A_25_153( .carry(c_25_153), .sum(s_25_153), .in3(s_25_147), .in2(s_25_146), .in1(s_25_150) );
  Fadder_ A_25_154( .carry(c_25_154), .sum(s_25_154), .in3(c_24_139), .in2(c_24_140), .in1(s_25_151) );
  Fadder_ A_25_155( .carry(c_25_155), .sum(s_25_155), .in3(c_24_141), .in2(s_25_152), .in1(s_25_153) );
  Fadder_ A_25_156( .carry(c_25_156), .sum(s_25_156), .in3(c_24_142), .in2(s_25_154), .in1(c_24_143) );
  Fadder_ A_25_157( .carry(c[25]), .sum(s[25]), .in3(s_25_155), .in2(c_24_144), .in1(s_25_156) );

  // ***** Bit 26 ***** //
  Hadder_ A_26_158( .carry(c_26_158), .sum(s_26_158), .in2(inc[26]), .in1(P_13[0]) );
  Fadder_ A_26_159( .carry(c_26_159), .sum(s_26_159), .in3(P_12[2]), .in2(P_11[4]), .in1(P_10[6]) );
  Fadder_ A_26_160( .carry(c_26_160), .sum(s_26_160), .in3(P_9[8]), .in2(P_8[10]), .in1(P_7[12]) );
  Fadder_ A_26_161( .carry(c_26_161), .sum(s_26_161), .in3(P_6[14]), .in2(P_5[16]), .in1(P_4[18]) );
  Fadder_ A_26_162( .carry(c_26_162), .sum(s_26_162), .in3(P_3[20]), .in2(P_2[22]), .in1(P_1[24]) );
  Fadder_ A_26_163( .carry(c_26_163), .sum(s_26_163), .in3(P_0[26]), .in2(c_25_149), .in1(c_25_148) );
  Fadder_ A_26_164( .carry(c_26_164), .sum(s_26_164), .in3(c_25_147), .in2(c_25_146), .in1(s_26_158) );
  Fadder_ A_26_165( .carry(c_26_165), .sum(s_26_165), .in3(s_26_162), .in2(s_26_161), .in1(s_26_160) );
  Fadder_ A_26_166( .carry(c_26_166), .sum(s_26_166), .in3(s_26_159), .in2(c_25_150), .in1(c_25_151) );
  Fadder_ A_26_167( .carry(c_26_167), .sum(s_26_167), .in3(s_26_163), .in2(c_25_152), .in1(s_26_164) );
  Fadder_ A_26_168( .carry(c_26_168), .sum(s_26_168), .in3(s_26_165), .in2(c_25_153), .in1(s_26_166) );
  Fadder_ A_26_169( .carry(c_26_169), .sum(s_26_169), .in3(c_25_154), .in2(s_26_167), .in1(c_25_155) );
  Fadder_ A_26_170( .carry(c[26]), .sum(s[26]), .in3(s_26_168), .in2(c_25_156), .in1(s_26_169) );

  // ***** Bit 27 ***** //
  Fadder_ A_27_171( .carry(c_27_171), .sum(s_27_171), .in3(inc[27]), .in2(P_13[1]), .in1(P_12[3]) );
  Fadder_ A_27_172( .carry(c_27_172), .sum(s_27_172), .in3(P_11[5]), .in2(P_10[7]), .in1(P_9[9]) );
  Fadder_ A_27_173( .carry(c_27_173), .sum(s_27_173), .in3(P_8[11]), .in2(P_7[13]), .in1(P_6[15]) );
  Fadder_ A_27_174( .carry(c_27_174), .sum(s_27_174), .in3(P_5[17]), .in2(P_4[19]), .in1(P_3[21]) );
  Fadder_ A_27_175( .carry(c_27_175), .sum(s_27_175), .in3(P_2[23]), .in2(P_1[25]), .in1(P_0[27]) );
  Fadder_ A_27_176( .carry(c_27_176), .sum(s_27_176), .in3(c_26_158), .in2(c_26_162), .in1(c_26_161) );
  Fadder_ A_27_177( .carry(c_27_177), .sum(s_27_177), .in3(c_26_160), .in2(c_26_159), .in1(s_27_175) );
  Fadder_ A_27_178( .carry(c_27_178), .sum(s_27_178), .in3(s_27_174), .in2(s_27_173), .in1(s_27_172) );
  Fadder_ A_27_179( .carry(c_27_179), .sum(s_27_179), .in3(s_27_171), .in2(c_26_163), .in1(c_26_164) );
  Fadder_ A_27_180( .carry(c_27_180), .sum(s_27_180), .in3(s_27_176), .in2(c_26_165), .in1(s_27_177) );
  Fadder_ A_27_181( .carry(c_27_181), .sum(s_27_181), .in3(s_27_178), .in2(c_26_166), .in1(s_27_179) );
  Fadder_ A_27_182( .carry(c_27_182), .sum(s_27_182), .in3(c_26_167), .in2(s_27_180), .in1(c_26_168) );
  Fadder_ A_27_183( .carry(c[27]), .sum(s[27]), .in3(s_27_181), .in2(c_26_169), .in1(s_27_182) );

  // ***** Bit 28 ***** //
  Hadder_ A_28_184( .carry(c_28_184), .sum(s_28_184), .in2(inc[28]), .in1(P_14[0]) );
  Fadder_ A_28_185( .carry(c_28_185), .sum(s_28_185), .in3(P_13[2]), .in2(P_12[4]), .in1(P_11[6]) );
  Fadder_ A_28_186( .carry(c_28_186), .sum(s_28_186), .in3(P_10[8]), .in2(P_9[10]), .in1(P_8[12]) );
  Fadder_ A_28_187( .carry(c_28_187), .sum(s_28_187), .in3(P_7[14]), .in2(P_6[16]), .in1(P_5[18]) );
  Fadder_ A_28_188( .carry(c_28_188), .sum(s_28_188), .in3(P_4[20]), .in2(P_3[22]), .in1(P_2[24]) );
  Fadder_ A_28_189( .carry(c_28_189), .sum(s_28_189), .in3(P_1[26]), .in2(P_0[28]), .in1(c_27_175) );
  Fadder_ A_28_190( .carry(c_28_190), .sum(s_28_190), .in3(c_27_174), .in2(c_27_173), .in1(c_27_172) );
  Fadder_ A_28_191( .carry(c_28_191), .sum(s_28_191), .in3(c_27_171), .in2(s_28_184), .in1(s_28_188) );
  Fadder_ A_28_192( .carry(c_28_192), .sum(s_28_192), .in3(s_28_187), .in2(s_28_186), .in1(s_28_185) );
  Fadder_ A_28_193( .carry(c_28_193), .sum(s_28_193), .in3(c_27_176), .in2(c_27_177), .in1(s_28_189) );
  Fadder_ A_28_194( .carry(c_28_194), .sum(s_28_194), .in3(s_28_190), .in2(c_27_178), .in1(s_28_191) );
  Fadder_ A_28_195( .carry(c_28_195), .sum(s_28_195), .in3(s_28_192), .in2(c_27_179), .in1(c_27_180) );
  Fadder_ A_28_196( .carry(c_28_196), .sum(s_28_196), .in3(s_28_193), .in2(s_28_194), .in1(c_27_181) );
  Fadder_ A_28_197( .carry(c[28]), .sum(s[28]), .in3(s_28_195), .in2(c_27_182), .in1(s_28_196) );

  // ***** Bit 29 ***** //
  Fadder_ A_29_198( .carry(c_29_198), .sum(s_29_198), .in3(inc[29]), .in2(P_14[1]), .in1(P_13[3]) );
  Fadder_ A_29_199( .carry(c_29_199), .sum(s_29_199), .in3(P_12[5]), .in2(P_11[7]), .in1(P_10[9]) );
  Fadder_ A_29_200( .carry(c_29_200), .sum(s_29_200), .in3(P_9[11]), .in2(P_8[13]), .in1(P_7[15]) );
  Fadder_ A_29_201( .carry(c_29_201), .sum(s_29_201), .in3(P_6[17]), .in2(P_5[19]), .in1(P_4[21]) );
  Fadder_ A_29_202( .carry(c_29_202), .sum(s_29_202), .in3(P_3[23]), .in2(P_2[25]), .in1(P_1[27]) );
  Fadder_ A_29_203( .carry(c_29_203), .sum(s_29_203), .in3(P_0[29]), .in2(c_28_184), .in1(c_28_188) );
  Fadder_ A_29_204( .carry(c_29_204), .sum(s_29_204), .in3(c_28_187), .in2(c_28_186), .in1(c_28_185) );
  Fadder_ A_29_205( .carry(c_29_205), .sum(s_29_205), .in3(s_29_202), .in2(s_29_201), .in1(s_29_200) );
  Fadder_ A_29_206( .carry(c_29_206), .sum(s_29_206), .in3(s_29_199), .in2(s_29_198), .in1(c_28_189) );
  Fadder_ A_29_207( .carry(c_29_207), .sum(s_29_207), .in3(c_28_190), .in2(s_29_203), .in1(c_28_191) );
  Fadder_ A_29_208( .carry(c_29_208), .sum(s_29_208), .in3(s_29_204), .in2(c_28_192), .in1(s_29_205) );
  Fadder_ A_29_209( .carry(c_29_209), .sum(s_29_209), .in3(s_29_206), .in2(c_28_193), .in1(c_28_194) );
  Fadder_ A_29_210( .carry(c_29_210), .sum(s_29_210), .in3(s_29_207), .in2(s_29_208), .in1(c_28_195) );
  Fadder_ A_29_211( .carry(c[29]), .sum(s[29]), .in3(s_29_209), .in2(c_28_196), .in1(s_29_210) );

  // ***** Bit 30 ***** //
  Hadder_ A_30_212( .carry(c_30_212), .sum(s_30_212), .in2(inc[30]), .in1(P_15[0]) );
  Fadder_ A_30_213( .carry(c_30_213), .sum(s_30_213), .in3(P_14[2]), .in2(P_13[4]), .in1(P_12[6]) );
  Fadder_ A_30_214( .carry(c_30_214), .sum(s_30_214), .in3(P_11[8]), .in2(P_10[10]), .in1(P_9[12]) );
  Fadder_ A_30_215( .carry(c_30_215), .sum(s_30_215), .in3(P_8[14]), .in2(P_7[16]), .in1(P_6[18]) );
  Fadder_ A_30_216( .carry(c_30_216), .sum(s_30_216), .in3(P_5[20]), .in2(P_4[22]), .in1(P_3[24]) );
  Fadder_ A_30_217( .carry(c_30_217), .sum(s_30_217), .in3(P_2[26]), .in2(P_1[28]), .in1(P_0[30]) );
  Fadder_ A_30_218( .carry(c_30_218), .sum(s_30_218), .in3(c_29_202), .in2(c_29_201), .in1(c_29_200) );
  Fadder_ A_30_219( .carry(c_30_219), .sum(s_30_219), .in3(c_29_199), .in2(c_29_198), .in1(s_30_212) );
  Fadder_ A_30_220( .carry(c_30_220), .sum(s_30_220), .in3(s_30_217), .in2(s_30_216), .in1(s_30_215) );
  Fadder_ A_30_221( .carry(c_30_221), .sum(s_30_221), .in3(s_30_214), .in2(s_30_213), .in1(c_29_203) );
  Fadder_ A_30_222( .carry(c_30_222), .sum(s_30_222), .in3(c_29_204), .in2(s_30_218), .in1(c_29_205) );
  Fadder_ A_30_223( .carry(c_30_223), .sum(s_30_223), .in3(s_30_219), .in2(s_30_220), .in1(c_29_206) );
  Fadder_ A_30_224( .carry(c_30_224), .sum(s_30_224), .in3(s_30_221), .in2(c_29_207), .in1(c_29_208) );
  Fadder_ A_30_225( .carry(c_30_225), .sum(s_30_225), .in3(s_30_222), .in2(s_30_223), .in1(c_29_209) );
  Fadder_ A_30_226( .carry(c[30]), .sum(s[30]), .in3(s_30_224), .in2(c_29_210), .in1(s_30_225) );

  // ***** Bit 31 ***** //
  Fadder_ A_31_227( .carry(c_31_227), .sum(s_31_227), .in3(inc[31]), .in2(P_15[1]), .in1(P_14[3]) );
  Fadder_ A_31_228( .carry(c_31_228), .sum(s_31_228), .in3(P_13[5]), .in2(P_12[7]), .in1(P_11[9]) );
  Fadder_ A_31_229( .carry(c_31_229), .sum(s_31_229), .in3(P_10[11]), .in2(P_9[13]), .in1(P_8[15]) );
  Fadder_ A_31_230( .carry(c_31_230), .sum(s_31_230), .in3(P_7[17]), .in2(P_6[19]), .in1(P_5[21]) );
  Fadder_ A_31_231( .carry(c_31_231), .sum(s_31_231), .in3(P_4[23]), .in2(P_3[25]), .in1(P_2[27]) );
  Fadder_ A_31_232( .carry(c_31_232), .sum(s_31_232), .in3(P_1[29]), .in2(P_0[31]), .in1(c_30_212) );
  Fadder_ A_31_233( .carry(c_31_233), .sum(s_31_233), .in3(c_30_217), .in2(c_30_216), .in1(c_30_215) );
  Fadder_ A_31_234( .carry(c_31_234), .sum(s_31_234), .in3(c_30_214), .in2(c_30_213), .in1(s_31_231) );
  Fadder_ A_31_235( .carry(c_31_235), .sum(s_31_235), .in3(s_31_230), .in2(s_31_229), .in1(s_31_228) );
  Fadder_ A_31_236( .carry(c_31_236), .sum(s_31_236), .in3(s_31_227), .in2(s_31_232), .in1(c_30_218) );
  Fadder_ A_31_237( .carry(c_31_237), .sum(s_31_237), .in3(c_30_219), .in2(s_31_233), .in1(c_30_220) );
  Fadder_ A_31_238( .carry(c_31_238), .sum(s_31_238), .in3(s_31_234), .in2(s_31_235), .in1(c_30_221) );
  Fadder_ A_31_239( .carry(c_31_239), .sum(s_31_239), .in3(s_31_236), .in2(c_30_222), .in1(s_31_237) );
  Fadder_ A_31_240( .carry(c_31_240), .sum(s_31_240), .in3(c_30_223), .in2(s_31_238), .in1(c_30_224) );
  Fadder_ A_31_241( .carry(c[31]), .sum(s[31]), .in3(s_31_239), .in2(c_30_225), .in1(s_31_240) );

  // ***** Bit 32 ***** //
  Hadder_ A_32_242( .carry(c_32_242), .sum(s_32_242), .in2(inc[32]), .in1(P_16[0]) );
  Fadder_ A_32_243( .carry(c_32_243), .sum(s_32_243), .in3(P_15[2]), .in2(P_14[4]), .in1(P_13[6]) );
  Fadder_ A_32_244( .carry(c_32_244), .sum(s_32_244), .in3(P_12[8]), .in2(P_11[10]), .in1(P_10[12]) );
  Fadder_ A_32_245( .carry(c_32_245), .sum(s_32_245), .in3(P_9[14]), .in2(P_8[16]), .in1(P_7[18]) );
  Fadder_ A_32_246( .carry(c_32_246), .sum(s_32_246), .in3(P_6[20]), .in2(P_5[22]), .in1(P_4[24]) );
  Fadder_ A_32_247( .carry(c_32_247), .sum(s_32_247), .in3(P_3[26]), .in2(P_2[28]), .in1(P_1[30]) );
  Fadder_ A_32_248( .carry(c_32_248), .sum(s_32_248), .in3(P_0[32]), .in2(c_31_231), .in1(c_31_230) );
  Fadder_ A_32_249( .carry(c_32_249), .sum(s_32_249), .in3(c_31_229), .in2(c_31_228), .in1(c_31_227) );
  Fadder_ A_32_250( .carry(c_32_250), .sum(s_32_250), .in3(s_32_242), .in2(s_32_247), .in1(s_32_246) );
  Fadder_ A_32_251( .carry(c_32_251), .sum(s_32_251), .in3(s_32_245), .in2(s_32_244), .in1(s_32_243) );
  Fadder_ A_32_252( .carry(c_32_252), .sum(s_32_252), .in3(c_31_232), .in2(c_31_233), .in1(c_31_234) );
  Fadder_ A_32_253( .carry(c_32_253), .sum(s_32_253), .in3(s_32_248), .in2(s_32_249), .in1(c_31_235) );
  Fadder_ A_32_254( .carry(c_32_254), .sum(s_32_254), .in3(s_32_250), .in2(s_32_251), .in1(c_31_236) );
  Fadder_ A_32_255( .carry(c_32_255), .sum(s_32_255), .in3(c_31_237), .in2(s_32_252), .in1(s_32_253) );
  Fadder_ A_32_256( .carry(c_32_256), .sum(s_32_256), .in3(c_31_238), .in2(s_32_254), .in1(c_31_239) );
  Fadder_ A_32_257( .carry(c[32]), .sum(s[32]), .in3(s_32_255), .in2(c_31_240), .in1(s_32_256) );

  // ***** Bit 33 ***** //
  Fadder_ A_33_258( .carry(c_33_258), .sum(s_33_258), .in3(inc[33]), .in2(P_16[1]), .in1(P_15[3]) );
  Fadder_ A_33_259( .carry(c_33_259), .sum(s_33_259), .in3(P_14[5]), .in2(P_13[7]), .in1(P_12[9]) );
  Fadder_ A_33_260( .carry(c_33_260), .sum(s_33_260), .in3(P_11[11]), .in2(P_10[13]), .in1(P_9[15]) );
  Fadder_ A_33_261( .carry(c_33_261), .sum(s_33_261), .in3(P_8[17]), .in2(P_7[19]), .in1(P_6[21]) );
  Fadder_ A_33_262( .carry(c_33_262), .sum(s_33_262), .in3(P_5[23]), .in2(P_4[25]), .in1(P_3[27]) );
  Fadder_ A_33_263( .carry(c_33_263), .sum(s_33_263), .in3(P_2[29]), .in2(P_1[31]), .in1(P_0[33]) );
  Fadder_ A_33_264( .carry(c_33_264), .sum(s_33_264), .in3(c_32_242), .in2(c_32_247), .in1(c_32_246) );
  Fadder_ A_33_265( .carry(c_33_265), .sum(s_33_265), .in3(c_32_245), .in2(c_32_244), .in1(c_32_243) );
  Fadder_ A_33_266( .carry(c_33_266), .sum(s_33_266), .in3(s_33_263), .in2(s_33_262), .in1(s_33_261) );
  Fadder_ A_33_267( .carry(c_33_267), .sum(s_33_267), .in3(s_33_260), .in2(s_33_259), .in1(s_33_258) );
  Fadder_ A_33_268( .carry(c_33_268), .sum(s_33_268), .in3(c_32_249), .in2(c_32_248), .in1(s_33_264) );
  Fadder_ A_33_269( .carry(c_33_269), .sum(s_33_269), .in3(s_33_265), .in2(c_32_251), .in1(c_32_250) );
  Fadder_ A_33_270( .carry(c_33_270), .sum(s_33_270), .in3(s_33_267), .in2(s_33_266), .in1(c_32_252) );
  Fadder_ A_33_271( .carry(c_33_271), .sum(s_33_271), .in3(c_32_253), .in2(s_33_268), .in1(s_33_269) );
  Fadder_ A_33_272( .carry(c_33_272), .sum(s_33_272), .in3(c_32_254), .in2(s_33_270), .in1(c_32_255) );
  Fadder_ A_33_273( .carry(c[33]), .sum(s[33]), .in3(s_33_271), .in2(c_32_256), .in1(s_33_272) );

  // ***** Bit 34 ***** //
  Hadder_ A_34_274( .carry(c_34_274), .sum(s_34_274), .in2(inc[34]), .in1(P_17[0]) );
  Fadder_ A_34_275( .carry(c_34_275), .sum(s_34_275), .in3(P_16[2]), .in2(P_15[4]), .in1(P_14[6]) );
  Fadder_ A_34_276( .carry(c_34_276), .sum(s_34_276), .in3(P_13[8]), .in2(P_12[10]), .in1(P_11[12]) );
  Fadder_ A_34_277( .carry(c_34_277), .sum(s_34_277), .in3(P_10[14]), .in2(P_9[16]), .in1(P_8[18]) );
  Fadder_ A_34_278( .carry(c_34_278), .sum(s_34_278), .in3(P_7[20]), .in2(P_6[22]), .in1(P_5[24]) );
  Fadder_ A_34_279( .carry(c_34_279), .sum(s_34_279), .in3(P_4[26]), .in2(P_3[28]), .in1(P_2[30]) );
  Fadder_ A_34_280( .carry(c_34_280), .sum(s_34_280), .in3(P_1[32]), .in2(P_0[34]), .in1(c_33_263) );
  Fadder_ A_34_281( .carry(c_34_281), .sum(s_34_281), .in3(c_33_262), .in2(c_33_261), .in1(c_33_260) );
  Fadder_ A_34_282( .carry(c_34_282), .sum(s_34_282), .in3(c_33_259), .in2(c_33_258), .in1(s_34_274) );
  Fadder_ A_34_283( .carry(c_34_283), .sum(s_34_283), .in3(s_34_279), .in2(s_34_278), .in1(s_34_277) );
  Fadder_ A_34_284( .carry(c_34_284), .sum(s_34_284), .in3(s_34_276), .in2(s_34_275), .in1(c_33_265) );
  Fadder_ A_34_285( .carry(c_34_285), .sum(s_34_285), .in3(c_33_264), .in2(s_34_280), .in1(s_34_281) );
  Fadder_ A_34_286( .carry(c_34_286), .sum(s_34_286), .in3(c_33_267), .in2(c_33_266), .in1(s_34_282) );
  Fadder_ A_34_287( .carry(c_34_287), .sum(s_34_287), .in3(s_34_283), .in2(c_33_268), .in1(s_34_284) );
  Fadder_ A_34_288( .carry(c_34_288), .sum(s_34_288), .in3(c_33_269), .in2(s_34_285), .in1(s_34_286) );
  Fadder_ A_34_289( .carry(c_34_289), .sum(s_34_289), .in3(c_33_270), .in2(s_34_287), .in1(c_33_271) );
  Fadder_ A_34_290( .carry(c[34]), .sum(s[34]), .in3(s_34_288), .in2(c_33_272), .in1(s_34_289) );

  // ***** Bit 35 ***** //
  Fadder_ A_35_291( .carry(c_35_291), .sum(s_35_291), .in3(inc[35]), .in2(P_17[1]), .in1(P_16[3]) );
  Fadder_ A_35_292( .carry(c_35_292), .sum(s_35_292), .in3(P_15[5]), .in2(P_14[7]), .in1(P_13[9]) );
  Fadder_ A_35_293( .carry(c_35_293), .sum(s_35_293), .in3(P_12[11]), .in2(P_11[13]), .in1(P_10[15]) );
  Fadder_ A_35_294( .carry(c_35_294), .sum(s_35_294), .in3(P_9[17]), .in2(P_8[19]), .in1(P_7[21]) );
  Fadder_ A_35_295( .carry(c_35_295), .sum(s_35_295), .in3(P_6[23]), .in2(P_5[25]), .in1(P_4[27]) );
  Fadder_ A_35_296( .carry(c_35_296), .sum(s_35_296), .in3(P_3[29]), .in2(P_2[31]), .in1(P_1[33]) );
  Fadder_ A_35_297( .carry(c_35_297), .sum(s_35_297), .in3(P_0[35]), .in2(c_34_274), .in1(c_34_279) );
  Fadder_ A_35_298( .carry(c_35_298), .sum(s_35_298), .in3(c_34_278), .in2(c_34_277), .in1(c_34_276) );
  Fadder_ A_35_299( .carry(c_35_299), .sum(s_35_299), .in3(c_34_275), .in2(s_35_296), .in1(s_35_295) );
  Fadder_ A_35_300( .carry(c_35_300), .sum(s_35_300), .in3(s_35_294), .in2(s_35_293), .in1(s_35_292) );
  Fadder_ A_35_301( .carry(c_35_301), .sum(s_35_301), .in3(s_35_291), .in2(c_34_280), .in1(c_34_281) );
  Fadder_ A_35_302( .carry(c_35_302), .sum(s_35_302), .in3(c_34_282), .in2(s_35_297), .in1(s_35_298) );
  Fadder_ A_35_303( .carry(c_35_303), .sum(s_35_303), .in3(c_34_283), .in2(s_35_299), .in1(s_35_300) );
  Fadder_ A_35_304( .carry(c_35_304), .sum(s_35_304), .in3(c_34_284), .in2(s_35_301), .in1(c_34_285) );
  Fadder_ A_35_305( .carry(c_35_305), .sum(s_35_305), .in3(c_34_286), .in2(s_35_302), .in1(s_35_303) );
  Fadder_ A_35_306( .carry(c_35_306), .sum(s_35_306), .in3(c_34_287), .in2(s_35_304), .in1(c_34_288) );
  Fadder_ A_35_307( .carry(c[35]), .sum(s[35]), .in3(s_35_305), .in2(c_34_289), .in1(s_35_306) );

  // ***** Bit 36 ***** //
  Hadder_ A_36_308( .carry(c_36_308), .sum(s_36_308), .in2(inc[36]), .in1(P_18[0]) );
  Fadder_ A_36_309( .carry(c_36_309), .sum(s_36_309), .in3(P_17[2]), .in2(P_16[4]), .in1(P_15[6]) );
  Fadder_ A_36_310( .carry(c_36_310), .sum(s_36_310), .in3(P_14[8]), .in2(P_13[10]), .in1(P_12[12]) );
  Fadder_ A_36_311( .carry(c_36_311), .sum(s_36_311), .in3(P_11[14]), .in2(P_10[16]), .in1(P_9[18]) );
  Fadder_ A_36_312( .carry(c_36_312), .sum(s_36_312), .in3(P_8[20]), .in2(P_7[22]), .in1(P_6[24]) );
  Fadder_ A_36_313( .carry(c_36_313), .sum(s_36_313), .in3(P_5[26]), .in2(P_4[28]), .in1(P_3[30]) );
  Fadder_ A_36_314( .carry(c_36_314), .sum(s_36_314), .in3(P_2[32]), .in2(P_1[34]), .in1(P_0[36]) );
  Fadder_ A_36_315( .carry(c_36_315), .sum(s_36_315), .in3(c_35_296), .in2(c_35_295), .in1(c_35_294) );
  Fadder_ A_36_316( .carry(c_36_316), .sum(s_36_316), .in3(c_35_293), .in2(c_35_292), .in1(c_35_291) );
  Fadder_ A_36_317( .carry(c_36_317), .sum(s_36_317), .in3(s_36_308), .in2(s_36_314), .in1(s_36_313) );
  Fadder_ A_36_318( .carry(c_36_318), .sum(s_36_318), .in3(s_36_312), .in2(s_36_311), .in1(s_36_310) );
  Fadder_ A_36_319( .carry(c_36_319), .sum(s_36_319), .in3(s_36_309), .in2(c_35_297), .in1(c_35_298) );
  Fadder_ A_36_320( .carry(c_36_320), .sum(s_36_320), .in3(s_36_316), .in2(s_36_315), .in1(c_35_300) );
  Fadder_ A_36_321( .carry(c_36_321), .sum(s_36_321), .in3(c_35_299), .in2(s_36_317), .in1(s_36_318) );
  Fadder_ A_36_322( .carry(c_36_322), .sum(s_36_322), .in3(c_35_301), .in2(s_36_319), .in1(c_35_302) );
  Fadder_ A_36_323( .carry(c_36_323), .sum(s_36_323), .in3(c_35_303), .in2(s_36_320), .in1(s_36_321) );
  Fadder_ A_36_324( .carry(c_36_324), .sum(s_36_324), .in3(c_35_304), .in2(s_36_322), .in1(c_35_305) );
  Fadder_ A_36_325( .carry(c[36]), .sum(s[36]), .in3(s_36_323), .in2(c_35_306), .in1(s_36_324) );

  // ***** Bit 37 ***** //
  Fadder_ A_37_326( .carry(c_37_326), .sum(s_37_326), .in3(inc[37]), .in2(P_18[1]), .in1(P_17[3]) );
  Fadder_ A_37_327( .carry(c_37_327), .sum(s_37_327), .in3(P_16[5]), .in2(P_15[7]), .in1(P_14[9]) );
  Fadder_ A_37_328( .carry(c_37_328), .sum(s_37_328), .in3(P_13[11]), .in2(P_12[13]), .in1(P_11[15]) );
  Fadder_ A_37_329( .carry(c_37_329), .sum(s_37_329), .in3(P_10[17]), .in2(P_9[19]), .in1(P_8[21]) );
  Fadder_ A_37_330( .carry(c_37_330), .sum(s_37_330), .in3(P_7[23]), .in2(P_6[25]), .in1(P_5[27]) );
  Fadder_ A_37_331( .carry(c_37_331), .sum(s_37_331), .in3(P_4[29]), .in2(P_3[31]), .in1(P_2[33]) );
  Fadder_ A_37_332( .carry(c_37_332), .sum(s_37_332), .in3(P_1[35]), .in2(P_0[37]), .in1(c_36_308) );
  Fadder_ A_37_333( .carry(c_37_333), .sum(s_37_333), .in3(c_36_314), .in2(c_36_313), .in1(c_36_312) );
  Fadder_ A_37_334( .carry(c_37_334), .sum(s_37_334), .in3(c_36_311), .in2(c_36_310), .in1(c_36_309) );
  Fadder_ A_37_335( .carry(c_37_335), .sum(s_37_335), .in3(s_37_331), .in2(s_37_330), .in1(s_37_329) );
  Fadder_ A_37_336( .carry(c_37_336), .sum(s_37_336), .in3(s_37_328), .in2(s_37_327), .in1(s_37_326) );
  Fadder_ A_37_337( .carry(c_37_337), .sum(s_37_337), .in3(s_37_332), .in2(c_36_316), .in1(c_36_315) );
  Fadder_ A_37_338( .carry(c_37_338), .sum(s_37_338), .in3(s_37_334), .in2(s_37_333), .in1(c_36_318) );
  Fadder_ A_37_339( .carry(c_37_339), .sum(s_37_339), .in3(c_36_317), .in2(s_37_336), .in1(s_37_335) );
  Fadder_ A_37_340( .carry(c_37_340), .sum(s_37_340), .in3(c_36_319), .in2(s_37_337), .in1(c_36_320) );
  Fadder_ A_37_341( .carry(c_37_341), .sum(s_37_341), .in3(c_36_321), .in2(s_37_338), .in1(s_37_339) );
  Fadder_ A_37_342( .carry(c_37_342), .sum(s_37_342), .in3(c_36_322), .in2(s_37_340), .in1(c_36_323) );
  Fadder_ A_37_343( .carry(c[37]), .sum(s[37]), .in3(s_37_341), .in2(c_36_324), .in1(s_37_342) );

  // ***** Bit 38 ***** //
  Hadder_ A_38_344( .carry(c_38_344), .sum(s_38_344), .in2(inc[38]), .in1(P_19[0]) );
  Fadder_ A_38_345( .carry(c_38_345), .sum(s_38_345), .in3(P_18[2]), .in2(P_17[4]), .in1(P_16[6]) );
  Fadder_ A_38_346( .carry(c_38_346), .sum(s_38_346), .in3(P_15[8]), .in2(P_14[10]), .in1(P_13[12]) );
  Fadder_ A_38_347( .carry(c_38_347), .sum(s_38_347), .in3(P_12[14]), .in2(P_11[16]), .in1(P_10[18]) );
  Fadder_ A_38_348( .carry(c_38_348), .sum(s_38_348), .in3(P_9[20]), .in2(P_8[22]), .in1(P_7[24]) );
  Fadder_ A_38_349( .carry(c_38_349), .sum(s_38_349), .in3(P_6[26]), .in2(P_5[28]), .in1(P_4[30]) );
  Fadder_ A_38_350( .carry(c_38_350), .sum(s_38_350), .in3(P_3[32]), .in2(P_2[34]), .in1(P_1[36]) );
  Fadder_ A_38_351( .carry(c_38_351), .sum(s_38_351), .in3(P_0[38]), .in2(c_37_331), .in1(c_37_330) );
  Fadder_ A_38_352( .carry(c_38_352), .sum(s_38_352), .in3(c_37_329), .in2(c_37_328), .in1(c_37_327) );
  Fadder_ A_38_353( .carry(c_38_353), .sum(s_38_353), .in3(c_37_326), .in2(s_38_344), .in1(s_38_350) );
  Fadder_ A_38_354( .carry(c_38_354), .sum(s_38_354), .in3(s_38_349), .in2(s_38_348), .in1(s_38_347) );
  Fadder_ A_38_355( .carry(c_38_355), .sum(s_38_355), .in3(s_38_346), .in2(s_38_345), .in1(c_37_332) );
  Fadder_ A_38_356( .carry(c_38_356), .sum(s_38_356), .in3(c_37_334), .in2(c_37_333), .in1(s_38_351) );
  Fadder_ A_38_357( .carry(c_38_357), .sum(s_38_357), .in3(s_38_352), .in2(c_37_336), .in1(c_37_335) );
  Fadder_ A_38_358( .carry(c_38_358), .sum(s_38_358), .in3(s_38_353), .in2(s_38_354), .in1(s_38_355) );
  Fadder_ A_38_359( .carry(c_38_359), .sum(s_38_359), .in3(c_37_337), .in2(c_37_338), .in1(s_38_356) );
  Fadder_ A_38_360( .carry(c_38_360), .sum(s_38_360), .in3(s_38_357), .in2(c_37_339), .in1(s_38_358) );
  Fadder_ A_38_361( .carry(c_38_361), .sum(s_38_361), .in3(c_37_340), .in2(c_37_341), .in1(s_38_359) );
  Fadder_ A_38_362( .carry(c[38]), .sum(s[38]), .in3(s_38_360), .in2(c_37_342), .in1(s_38_361) );

  // ***** Bit 39 ***** //
  Fadder_ A_39_363( .carry(c_39_363), .sum(s_39_363), .in3(inc[39]), .in2(P_19[1]), .in1(P_18[3]) );
  Fadder_ A_39_364( .carry(c_39_364), .sum(s_39_364), .in3(P_17[5]), .in2(P_16[7]), .in1(P_15[9]) );
  Fadder_ A_39_365( .carry(c_39_365), .sum(s_39_365), .in3(P_14[11]), .in2(P_13[13]), .in1(P_12[15]) );
  Fadder_ A_39_366( .carry(c_39_366), .sum(s_39_366), .in3(P_11[17]), .in2(P_10[19]), .in1(P_9[21]) );
  Fadder_ A_39_367( .carry(c_39_367), .sum(s_39_367), .in3(P_8[23]), .in2(P_7[25]), .in1(P_6[27]) );
  Fadder_ A_39_368( .carry(c_39_368), .sum(s_39_368), .in3(P_5[29]), .in2(P_4[31]), .in1(P_3[33]) );
  Fadder_ A_39_369( .carry(c_39_369), .sum(s_39_369), .in3(P_2[35]), .in2(P_1[37]), .in1(P_0[39]) );
  Fadder_ A_39_370( .carry(c_39_370), .sum(s_39_370), .in3(c_38_344), .in2(c_38_350), .in1(c_38_349) );
  Fadder_ A_39_371( .carry(c_39_371), .sum(s_39_371), .in3(c_38_348), .in2(c_38_347), .in1(c_38_346) );
  Fadder_ A_39_372( .carry(c_39_372), .sum(s_39_372), .in3(c_38_345), .in2(s_39_369), .in1(s_39_368) );
  Fadder_ A_39_373( .carry(c_39_373), .sum(s_39_373), .in3(s_39_367), .in2(s_39_366), .in1(s_39_365) );
  Fadder_ A_39_374( .carry(c_39_374), .sum(s_39_374), .in3(s_39_364), .in2(s_39_363), .in1(c_38_352) );
  Fadder_ A_39_375( .carry(c_39_375), .sum(s_39_375), .in3(c_38_351), .in2(s_39_370), .in1(c_38_353) );
  Fadder_ A_39_376( .carry(c_39_376), .sum(s_39_376), .in3(s_39_371), .in2(c_38_354), .in1(c_38_355) );
  Fadder_ A_39_377( .carry(c_39_377), .sum(s_39_377), .in3(s_39_372), .in2(s_39_373), .in1(c_38_356) );
  Fadder_ A_39_378( .carry(c_39_378), .sum(s_39_378), .in3(s_39_374), .in2(c_38_357), .in1(s_39_375) );
  Fadder_ A_39_379( .carry(c_39_379), .sum(s_39_379), .in3(s_39_376), .in2(c_38_358), .in1(s_39_377) );
  Fadder_ A_39_380( .carry(c_39_380), .sum(s_39_380), .in3(c_38_359), .in2(s_39_378), .in1(c_38_360) );
  Fadder_ A_39_381( .carry(c[39]), .sum(s[39]), .in3(s_39_379), .in2(c_38_361), .in1(s_39_380) );

  // ***** Bit 40 ***** //
  Hadder_ A_40_382( .carry(c_40_382), .sum(s_40_382), .in2(inc[40]), .in1(P_20[0]) );
  Fadder_ A_40_383( .carry(c_40_383), .sum(s_40_383), .in3(P_19[2]), .in2(P_18[4]), .in1(P_17[6]) );
  Fadder_ A_40_384( .carry(c_40_384), .sum(s_40_384), .in3(P_16[8]), .in2(P_15[10]), .in1(P_14[12]) );
  Fadder_ A_40_385( .carry(c_40_385), .sum(s_40_385), .in3(P_13[14]), .in2(P_12[16]), .in1(P_11[18]) );
  Fadder_ A_40_386( .carry(c_40_386), .sum(s_40_386), .in3(P_10[20]), .in2(P_9[22]), .in1(P_8[24]) );
  Fadder_ A_40_387( .carry(c_40_387), .sum(s_40_387), .in3(P_7[26]), .in2(P_6[28]), .in1(P_5[30]) );
  Fadder_ A_40_388( .carry(c_40_388), .sum(s_40_388), .in3(P_4[32]), .in2(P_3[34]), .in1(P_2[36]) );
  Fadder_ A_40_389( .carry(c_40_389), .sum(s_40_389), .in3(P_1[38]), .in2(P_0[40]), .in1(c_39_369) );
  Fadder_ A_40_390( .carry(c_40_390), .sum(s_40_390), .in3(c_39_368), .in2(c_39_367), .in1(c_39_366) );
  Fadder_ A_40_391( .carry(c_40_391), .sum(s_40_391), .in3(c_39_365), .in2(c_39_364), .in1(c_39_363) );
  Fadder_ A_40_392( .carry(c_40_392), .sum(s_40_392), .in3(s_40_382), .in2(s_40_388), .in1(s_40_387) );
  Fadder_ A_40_393( .carry(c_40_393), .sum(s_40_393), .in3(s_40_386), .in2(s_40_385), .in1(s_40_384) );
  Fadder_ A_40_394( .carry(c_40_394), .sum(s_40_394), .in3(s_40_383), .in2(c_39_371), .in1(c_39_370) );
  Fadder_ A_40_395( .carry(c_40_395), .sum(s_40_395), .in3(s_40_389), .in2(s_40_391), .in1(s_40_390) );
  Fadder_ A_40_396( .carry(c_40_396), .sum(s_40_396), .in3(c_39_373), .in2(c_39_372), .in1(s_40_392) );
  Fadder_ A_40_397( .carry(c_40_397), .sum(s_40_397), .in3(s_40_393), .in2(c_39_374), .in1(s_40_394) );
  Fadder_ A_40_398( .carry(c_40_398), .sum(s_40_398), .in3(c_39_375), .in2(c_39_376), .in1(s_40_395) );
  Fadder_ A_40_399( .carry(c_40_399), .sum(s_40_399), .in3(s_40_396), .in2(c_39_377), .in1(c_39_378) );
  Fadder_ A_40_400( .carry(c_40_400), .sum(s_40_400), .in3(s_40_397), .in2(s_40_398), .in1(c_39_379) );
  Fadder_ A_40_401( .carry(c[40]), .sum(s[40]), .in3(s_40_399), .in2(c_39_380), .in1(s_40_400) );

  // ***** Bit 41 ***** //
  Fadder_ A_41_402( .carry(c_41_402), .sum(s_41_402), .in3(inc[41]), .in2(P_20[1]), .in1(P_19[3]) );
  Fadder_ A_41_403( .carry(c_41_403), .sum(s_41_403), .in3(P_18[5]), .in2(P_17[7]), .in1(P_16[9]) );
  Fadder_ A_41_404( .carry(c_41_404), .sum(s_41_404), .in3(P_15[11]), .in2(P_14[13]), .in1(P_13[15]) );
  Fadder_ A_41_405( .carry(c_41_405), .sum(s_41_405), .in3(P_12[17]), .in2(P_11[19]), .in1(P_10[21]) );
  Fadder_ A_41_406( .carry(c_41_406), .sum(s_41_406), .in3(P_9[23]), .in2(P_8[25]), .in1(P_7[27]) );
  Fadder_ A_41_407( .carry(c_41_407), .sum(s_41_407), .in3(P_6[29]), .in2(P_5[31]), .in1(P_4[33]) );
  Fadder_ A_41_408( .carry(c_41_408), .sum(s_41_408), .in3(P_3[35]), .in2(P_2[37]), .in1(P_1[39]) );
  Fadder_ A_41_409( .carry(c_41_409), .sum(s_41_409), .in3(P_0[41]), .in2(c_40_382), .in1(c_40_388) );
  Fadder_ A_41_410( .carry(c_41_410), .sum(s_41_410), .in3(c_40_387), .in2(c_40_386), .in1(c_40_385) );
  Fadder_ A_41_411( .carry(c_41_411), .sum(s_41_411), .in3(c_40_384), .in2(c_40_383), .in1(s_41_408) );
  Fadder_ A_41_412( .carry(c_41_412), .sum(s_41_412), .in3(s_41_407), .in2(s_41_406), .in1(s_41_405) );
  Fadder_ A_41_413( .carry(c_41_413), .sum(s_41_413), .in3(s_41_404), .in2(s_41_403), .in1(s_41_402) );
  Fadder_ A_41_414( .carry(c_41_414), .sum(s_41_414), .in3(c_40_389), .in2(c_40_391), .in1(c_40_390) );
  Fadder_ A_41_415( .carry(c_41_415), .sum(s_41_415), .in3(s_41_409), .in2(s_41_410), .in1(c_40_393) );
  Fadder_ A_41_416( .carry(c_41_416), .sum(s_41_416), .in3(c_40_392), .in2(s_41_411), .in1(s_41_413) );
  Fadder_ A_41_417( .carry(c_41_417), .sum(s_41_417), .in3(s_41_412), .in2(c_40_394), .in1(s_41_414) );
  Fadder_ A_41_418( .carry(c_41_418), .sum(s_41_418), .in3(c_40_395), .in2(c_40_396), .in1(s_41_415) );
  Fadder_ A_41_419( .carry(c_41_419), .sum(s_41_419), .in3(s_41_416), .in2(c_40_397), .in1(c_40_398) );
  Fadder_ A_41_420( .carry(c_41_420), .sum(s_41_420), .in3(s_41_417), .in2(s_41_418), .in1(c_40_399) );
  Fadder_ A_41_421( .carry(c[41]), .sum(s[41]), .in3(s_41_419), .in2(c_40_400), .in1(s_41_420) );

  // ***** Bit 42 ***** //
  Hadder_ A_42_422( .carry(c_42_422), .sum(s_42_422), .in2(inc[42]), .in1(P_21[0]) );
  Fadder_ A_42_423( .carry(c_42_423), .sum(s_42_423), .in3(P_20[2]), .in2(P_19[4]), .in1(P_18[6]) );
  Fadder_ A_42_424( .carry(c_42_424), .sum(s_42_424), .in3(P_17[8]), .in2(P_16[10]), .in1(P_15[12]) );
  Fadder_ A_42_425( .carry(c_42_425), .sum(s_42_425), .in3(P_14[14]), .in2(P_13[16]), .in1(P_12[18]) );
  Fadder_ A_42_426( .carry(c_42_426), .sum(s_42_426), .in3(P_11[20]), .in2(P_10[22]), .in1(P_9[24]) );
  Fadder_ A_42_427( .carry(c_42_427), .sum(s_42_427), .in3(P_8[26]), .in2(P_7[28]), .in1(P_6[30]) );
  Fadder_ A_42_428( .carry(c_42_428), .sum(s_42_428), .in3(P_5[32]), .in2(P_4[34]), .in1(P_3[36]) );
  Fadder_ A_42_429( .carry(c_42_429), .sum(s_42_429), .in3(P_2[38]), .in2(P_1[40]), .in1(P_0[42]) );
  Fadder_ A_42_430( .carry(c_42_430), .sum(s_42_430), .in3(c_41_408), .in2(c_41_407), .in1(c_41_406) );
  Fadder_ A_42_431( .carry(c_42_431), .sum(s_42_431), .in3(c_41_405), .in2(c_41_404), .in1(c_41_403) );
  Fadder_ A_42_432( .carry(c_42_432), .sum(s_42_432), .in3(c_41_402), .in2(s_42_422), .in1(s_42_429) );
  Fadder_ A_42_433( .carry(c_42_433), .sum(s_42_433), .in3(s_42_428), .in2(s_42_427), .in1(s_42_426) );
  Fadder_ A_42_434( .carry(c_42_434), .sum(s_42_434), .in3(s_42_425), .in2(s_42_424), .in1(s_42_423) );
  Fadder_ A_42_435( .carry(c_42_435), .sum(s_42_435), .in3(c_41_409), .in2(c_41_410), .in1(c_41_411) );
  Fadder_ A_42_436( .carry(c_42_436), .sum(s_42_436), .in3(s_42_431), .in2(s_42_430), .in1(c_41_413) );
  Fadder_ A_42_437( .carry(c_42_437), .sum(s_42_437), .in3(c_41_412), .in2(s_42_432), .in1(s_42_434) );
  Fadder_ A_42_438( .carry(c_42_438), .sum(s_42_438), .in3(s_42_433), .in2(c_41_414), .in1(c_41_415) );
  Fadder_ A_42_439( .carry(c_42_439), .sum(s_42_439), .in3(s_42_435), .in2(c_41_416), .in1(s_42_436) );
  Fadder_ A_42_440( .carry(c_42_440), .sum(s_42_440), .in3(s_42_437), .in2(c_41_417), .in1(c_41_418) );
  Fadder_ A_42_441( .carry(c_42_441), .sum(s_42_441), .in3(s_42_438), .in2(s_42_439), .in1(c_41_419) );
  Fadder_ A_42_442( .carry(c[42]), .sum(s[42]), .in3(s_42_440), .in2(c_41_420), .in1(s_42_441) );

  // ***** Bit 43 ***** //
  Fadder_ A_43_443( .carry(c_43_443), .sum(s_43_443), .in3(inc[43]), .in2(P_21[1]), .in1(P_20[3]) );
  Fadder_ A_43_444( .carry(c_43_444), .sum(s_43_444), .in3(P_19[5]), .in2(P_18[7]), .in1(P_17[9]) );
  Fadder_ A_43_445( .carry(c_43_445), .sum(s_43_445), .in3(P_16[11]), .in2(P_15[13]), .in1(P_14[15]) );
  Fadder_ A_43_446( .carry(c_43_446), .sum(s_43_446), .in3(P_13[17]), .in2(P_12[19]), .in1(P_11[21]) );
  Fadder_ A_43_447( .carry(c_43_447), .sum(s_43_447), .in3(P_10[23]), .in2(P_9[25]), .in1(P_8[27]) );
  Fadder_ A_43_448( .carry(c_43_448), .sum(s_43_448), .in3(P_7[29]), .in2(P_6[31]), .in1(P_5[33]) );
  Fadder_ A_43_449( .carry(c_43_449), .sum(s_43_449), .in3(P_4[35]), .in2(P_3[37]), .in1(P_2[39]) );
  Fadder_ A_43_450( .carry(c_43_450), .sum(s_43_450), .in3(P_1[41]), .in2(P_0[43]), .in1(c_42_422) );
  Fadder_ A_43_451( .carry(c_43_451), .sum(s_43_451), .in3(c_42_429), .in2(c_42_428), .in1(c_42_427) );
  Fadder_ A_43_452( .carry(c_43_452), .sum(s_43_452), .in3(c_42_426), .in2(c_42_425), .in1(c_42_424) );
  Fadder_ A_43_453( .carry(c_43_453), .sum(s_43_453), .in3(c_42_423), .in2(s_43_449), .in1(s_43_448) );
  Fadder_ A_43_454( .carry(c_43_454), .sum(s_43_454), .in3(s_43_447), .in2(s_43_446), .in1(s_43_445) );
  Fadder_ A_43_455( .carry(c_43_455), .sum(s_43_455), .in3(s_43_444), .in2(s_43_443), .in1(s_43_450) );
  Fadder_ A_43_456( .carry(c_43_456), .sum(s_43_456), .in3(c_42_431), .in2(c_42_430), .in1(c_42_432) );
  Fadder_ A_43_457( .carry(c_43_457), .sum(s_43_457), .in3(s_43_452), .in2(s_43_451), .in1(c_42_434) );
  Fadder_ A_43_458( .carry(c_43_458), .sum(s_43_458), .in3(c_42_433), .in2(s_43_453), .in1(s_43_454) );
  Fadder_ A_43_459( .carry(c_43_459), .sum(s_43_459), .in3(s_43_455), .in2(c_42_435), .in1(c_42_436) );
  Fadder_ A_43_460( .carry(c_43_460), .sum(s_43_460), .in3(s_43_456), .in2(c_42_437), .in1(s_43_457) );
  Fadder_ A_43_461( .carry(c_43_461), .sum(s_43_461), .in3(s_43_458), .in2(c_42_438), .in1(s_43_459) );
  Fadder_ A_43_462( .carry(c_43_462), .sum(s_43_462), .in3(c_42_439), .in2(s_43_460), .in1(c_42_440) );
  Fadder_ A_43_463( .carry(c[43]), .sum(s[43]), .in3(s_43_461), .in2(c_42_441), .in1(s_43_462) );

  // ***** Bit 44 ***** //
  Hadder_ A_44_464( .carry(c_44_464), .sum(s_44_464), .in2(inc[44]), .in1(P_22[0]) );
  Fadder_ A_44_465( .carry(c_44_465), .sum(s_44_465), .in3(P_21[2]), .in2(P_20[4]), .in1(P_19[6]) );
  Fadder_ A_44_466( .carry(c_44_466), .sum(s_44_466), .in3(P_18[8]), .in2(P_17[10]), .in1(P_16[12]) );
  Fadder_ A_44_467( .carry(c_44_467), .sum(s_44_467), .in3(P_15[14]), .in2(P_14[16]), .in1(P_13[18]) );
  Fadder_ A_44_468( .carry(c_44_468), .sum(s_44_468), .in3(P_12[20]), .in2(P_11[22]), .in1(P_10[24]) );
  Fadder_ A_44_469( .carry(c_44_469), .sum(s_44_469), .in3(P_9[26]), .in2(P_8[28]), .in1(P_7[30]) );
  Fadder_ A_44_470( .carry(c_44_470), .sum(s_44_470), .in3(P_6[32]), .in2(P_5[34]), .in1(P_4[36]) );
  Fadder_ A_44_471( .carry(c_44_471), .sum(s_44_471), .in3(P_3[38]), .in2(P_2[40]), .in1(P_1[42]) );
  Fadder_ A_44_472( .carry(c_44_472), .sum(s_44_472), .in3(P_0[44]), .in2(c_43_449), .in1(c_43_448) );
  Fadder_ A_44_473( .carry(c_44_473), .sum(s_44_473), .in3(c_43_447), .in2(c_43_446), .in1(c_43_445) );
  Fadder_ A_44_474( .carry(c_44_474), .sum(s_44_474), .in3(c_43_444), .in2(c_43_443), .in1(s_44_464) );
  Fadder_ A_44_475( .carry(c_44_475), .sum(s_44_475), .in3(s_44_471), .in2(s_44_470), .in1(s_44_469) );
  Fadder_ A_44_476( .carry(c_44_476), .sum(s_44_476), .in3(s_44_468), .in2(s_44_467), .in1(s_44_466) );
  Fadder_ A_44_477( .carry(c_44_477), .sum(s_44_477), .in3(s_44_465), .in2(c_43_450), .in1(c_43_452) );
  Fadder_ A_44_478( .carry(c_44_478), .sum(s_44_478), .in3(c_43_451), .in2(s_44_472), .in1(s_44_473) );
  Fadder_ A_44_479( .carry(c_44_479), .sum(s_44_479), .in3(c_43_454), .in2(c_43_453), .in1(s_44_474) );
  Fadder_ A_44_480( .carry(c_44_480), .sum(s_44_480), .in3(s_44_476), .in2(s_44_475), .in1(c_43_455) );
  Fadder_ A_44_481( .carry(c_44_481), .sum(s_44_481), .in3(c_43_456), .in2(s_44_477), .in1(c_43_457) );
  Fadder_ A_44_482( .carry(c_44_482), .sum(s_44_482), .in3(s_44_478), .in2(c_43_458), .in1(s_44_479) );
  Fadder_ A_44_483( .carry(c_44_483), .sum(s_44_483), .in3(s_44_480), .in2(c_43_459), .in1(s_44_481) );
  Fadder_ A_44_484( .carry(c_44_484), .sum(s_44_484), .in3(c_43_460), .in2(s_44_482), .in1(c_43_461) );
  Fadder_ A_44_485( .carry(c[44]), .sum(s[44]), .in3(s_44_483), .in2(c_43_462), .in1(s_44_484) );

  // ***** Bit 45 ***** //
  Fadder_ A_45_486( .carry(c_45_486), .sum(s_45_486), .in3(inc[45]), .in2(P_22[1]), .in1(P_21[3]) );
  Fadder_ A_45_487( .carry(c_45_487), .sum(s_45_487), .in3(P_20[5]), .in2(P_19[7]), .in1(P_18[9]) );
  Fadder_ A_45_488( .carry(c_45_488), .sum(s_45_488), .in3(P_17[11]), .in2(P_16[13]), .in1(P_15[15]) );
  Fadder_ A_45_489( .carry(c_45_489), .sum(s_45_489), .in3(P_14[17]), .in2(P_13[19]), .in1(P_12[21]) );
  Fadder_ A_45_490( .carry(c_45_490), .sum(s_45_490), .in3(P_11[23]), .in2(P_10[25]), .in1(P_9[27]) );
  Fadder_ A_45_491( .carry(c_45_491), .sum(s_45_491), .in3(P_8[29]), .in2(P_7[31]), .in1(P_6[33]) );
  Fadder_ A_45_492( .carry(c_45_492), .sum(s_45_492), .in3(P_5[35]), .in2(P_4[37]), .in1(P_3[39]) );
  Fadder_ A_45_493( .carry(c_45_493), .sum(s_45_493), .in3(P_2[41]), .in2(P_1[43]), .in1(P_0[45]) );
  Fadder_ A_45_494( .carry(c_45_494), .sum(s_45_494), .in3(c_44_464), .in2(c_44_471), .in1(c_44_470) );
  Fadder_ A_45_495( .carry(c_45_495), .sum(s_45_495), .in3(c_44_469), .in2(c_44_468), .in1(c_44_467) );
  Fadder_ A_45_496( .carry(c_45_496), .sum(s_45_496), .in3(c_44_466), .in2(c_44_465), .in1(s_45_493) );
  Fadder_ A_45_497( .carry(c_45_497), .sum(s_45_497), .in3(s_45_492), .in2(s_45_491), .in1(s_45_490) );
  Fadder_ A_45_498( .carry(c_45_498), .sum(s_45_498), .in3(s_45_489), .in2(s_45_488), .in1(s_45_487) );
  Fadder_ A_45_499( .carry(c_45_499), .sum(s_45_499), .in3(s_45_486), .in2(c_44_473), .in1(c_44_472) );
  Fadder_ A_45_500( .carry(c_45_500), .sum(s_45_500), .in3(c_44_474), .in2(s_45_494), .in1(s_45_495) );
  Fadder_ A_45_501( .carry(c_45_501), .sum(s_45_501), .in3(c_44_476), .in2(c_44_475), .in1(s_45_496) );
  Fadder_ A_45_502( .carry(c_45_502), .sum(s_45_502), .in3(s_45_498), .in2(s_45_497), .in1(c_44_477) );
  Fadder_ A_45_503( .carry(c_45_503), .sum(s_45_503), .in3(s_45_499), .in2(c_44_478), .in1(c_44_479) );
  Fadder_ A_45_504( .carry(c_45_504), .sum(s_45_504), .in3(s_45_500), .in2(c_44_480), .in1(s_45_501) );
  Fadder_ A_45_505( .carry(c_45_505), .sum(s_45_505), .in3(s_45_502), .in2(c_44_481), .in1(s_45_503) );
  Fadder_ A_45_506( .carry(c_45_506), .sum(s_45_506), .in3(c_44_482), .in2(s_45_504), .in1(c_44_483) );
  Fadder_ A_45_507( .carry(c[45]), .sum(s[45]), .in3(s_45_505), .in2(c_44_484), .in1(s_45_506) );

  // ***** Bit 46 ***** //
  Hadder_ A_46_508( .carry(c_46_508), .sum(s_46_508), .in2(inc[46]), .in1(P_23[0]) );
  Fadder_ A_46_509( .carry(c_46_509), .sum(s_46_509), .in3(P_22[2]), .in2(P_21[4]), .in1(P_20[6]) );
  Fadder_ A_46_510( .carry(c_46_510), .sum(s_46_510), .in3(P_19[8]), .in2(P_18[10]), .in1(P_17[12]) );
  Fadder_ A_46_511( .carry(c_46_511), .sum(s_46_511), .in3(P_16[14]), .in2(P_15[16]), .in1(P_14[18]) );
  Fadder_ A_46_512( .carry(c_46_512), .sum(s_46_512), .in3(P_13[20]), .in2(P_12[22]), .in1(P_11[24]) );
  Fadder_ A_46_513( .carry(c_46_513), .sum(s_46_513), .in3(P_10[26]), .in2(P_9[28]), .in1(P_8[30]) );
  Fadder_ A_46_514( .carry(c_46_514), .sum(s_46_514), .in3(P_7[32]), .in2(P_6[34]), .in1(P_5[36]) );
  Fadder_ A_46_515( .carry(c_46_515), .sum(s_46_515), .in3(P_4[38]), .in2(P_3[40]), .in1(P_2[42]) );
  Fadder_ A_46_516( .carry(c_46_516), .sum(s_46_516), .in3(P_1[44]), .in2(P_0[46]), .in1(c_45_493) );
  Fadder_ A_46_517( .carry(c_46_517), .sum(s_46_517), .in3(c_45_492), .in2(c_45_491), .in1(c_45_490) );
  Fadder_ A_46_518( .carry(c_46_518), .sum(s_46_518), .in3(c_45_489), .in2(c_45_488), .in1(c_45_487) );
  Fadder_ A_46_519( .carry(c_46_519), .sum(s_46_519), .in3(c_45_486), .in2(s_46_508), .in1(s_46_515) );
  Fadder_ A_46_520( .carry(c_46_520), .sum(s_46_520), .in3(s_46_514), .in2(s_46_513), .in1(s_46_512) );
  Fadder_ A_46_521( .carry(c_46_521), .sum(s_46_521), .in3(s_46_511), .in2(s_46_510), .in1(s_46_509) );
  Fadder_ A_46_522( .carry(c_46_522), .sum(s_46_522), .in3(c_45_495), .in2(c_45_494), .in1(c_45_496) );
  Fadder_ A_46_523( .carry(c_46_523), .sum(s_46_523), .in3(s_46_516), .in2(s_46_518), .in1(s_46_517) );
  Fadder_ A_46_524( .carry(c_46_524), .sum(s_46_524), .in3(c_45_498), .in2(c_45_497), .in1(s_46_519) );
  Fadder_ A_46_525( .carry(c_46_525), .sum(s_46_525), .in3(s_46_521), .in2(s_46_520), .in1(c_45_499) );
  Fadder_ A_46_526( .carry(c_46_526), .sum(s_46_526), .in3(c_45_500), .in2(s_46_522), .in1(c_45_501) );
  Fadder_ A_46_527( .carry(c_46_527), .sum(s_46_527), .in3(s_46_523), .in2(s_46_524), .in1(c_45_502) );
  Fadder_ A_46_528( .carry(c_46_528), .sum(s_46_528), .in3(s_46_525), .in2(c_45_503), .in1(s_46_526) );
  Fadder_ A_46_529( .carry(c_46_529), .sum(s_46_529), .in3(c_45_504), .in2(s_46_527), .in1(c_45_505) );
  Fadder_ A_46_530( .carry(c[46]), .sum(s[46]), .in3(s_46_528), .in2(c_45_506), .in1(s_46_529) );

  // ***** Bit 47 ***** //
  Fadder_ A_47_531( .carry(c_47_531), .sum(s_47_531), .in3(inc[47]), .in2(P_23[1]), .in1(P_22[3]) );
  Fadder_ A_47_532( .carry(c_47_532), .sum(s_47_532), .in3(P_21[5]), .in2(P_20[7]), .in1(P_19[9]) );
  Fadder_ A_47_533( .carry(c_47_533), .sum(s_47_533), .in3(P_18[11]), .in2(P_17[13]), .in1(P_16[15]) );
  Fadder_ A_47_534( .carry(c_47_534), .sum(s_47_534), .in3(P_15[17]), .in2(P_14[19]), .in1(P_13[21]) );
  Fadder_ A_47_535( .carry(c_47_535), .sum(s_47_535), .in3(P_12[23]), .in2(P_11[25]), .in1(P_10[27]) );
  Fadder_ A_47_536( .carry(c_47_536), .sum(s_47_536), .in3(P_9[29]), .in2(P_8[31]), .in1(P_7[33]) );
  Fadder_ A_47_537( .carry(c_47_537), .sum(s_47_537), .in3(P_6[35]), .in2(P_5[37]), .in1(P_4[39]) );
  Fadder_ A_47_538( .carry(c_47_538), .sum(s_47_538), .in3(P_3[41]), .in2(P_2[43]), .in1(P_1[45]) );
  Fadder_ A_47_539( .carry(c_47_539), .sum(s_47_539), .in3(P_0[47]), .in2(c_46_508), .in1(c_46_515) );
  Fadder_ A_47_540( .carry(c_47_540), .sum(s_47_540), .in3(c_46_514), .in2(c_46_513), .in1(c_46_512) );
  Fadder_ A_47_541( .carry(c_47_541), .sum(s_47_541), .in3(c_46_511), .in2(c_46_510), .in1(c_46_509) );
  Fadder_ A_47_542( .carry(c_47_542), .sum(s_47_542), .in3(s_47_538), .in2(s_47_537), .in1(s_47_536) );
  Fadder_ A_47_543( .carry(c_47_543), .sum(s_47_543), .in3(s_47_535), .in2(s_47_534), .in1(s_47_533) );
  Fadder_ A_47_544( .carry(c_47_544), .sum(s_47_544), .in3(s_47_532), .in2(s_47_531), .in1(c_46_516) );
  Fadder_ A_47_545( .carry(c_47_545), .sum(s_47_545), .in3(c_46_518), .in2(c_46_517), .in1(s_47_539) );
  Fadder_ A_47_546( .carry(c_47_546), .sum(s_47_546), .in3(c_46_519), .in2(s_47_541), .in1(s_47_540) );
  Fadder_ A_47_547( .carry(c_47_547), .sum(s_47_547), .in3(c_46_521), .in2(c_46_520), .in1(s_47_543) );
  Fadder_ A_47_548( .carry(c_47_548), .sum(s_47_548), .in3(s_47_542), .in2(c_46_522), .in1(s_47_544) );
  Fadder_ A_47_549( .carry(c_47_549), .sum(s_47_549), .in3(c_46_523), .in2(c_46_524), .in1(s_47_545) );
  Fadder_ A_47_550( .carry(c_47_550), .sum(s_47_550), .in3(s_47_546), .in2(s_47_547), .in1(c_46_525) );
  Fadder_ A_47_551( .carry(c_47_551), .sum(s_47_551), .in3(s_47_548), .in2(c_46_526), .in1(s_47_549) );
  Fadder_ A_47_552( .carry(c_47_552), .sum(s_47_552), .in3(c_46_527), .in2(s_47_550), .in1(c_46_528) );
  Fadder_ A_47_553( .carry(c[47]), .sum(s[47]), .in3(s_47_551), .in2(c_46_529), .in1(s_47_552) );

  // ***** Bit 48 ***** //
  Hadder_ A_48_554( .carry(c_48_554), .sum(s_48_554), .in2(inc[48]), .in1(P_24[0]) );
  Fadder_ A_48_555( .carry(c_48_555), .sum(s_48_555), .in3(P_23[2]), .in2(P_22[4]), .in1(P_21[6]) );
  Fadder_ A_48_556( .carry(c_48_556), .sum(s_48_556), .in3(P_20[8]), .in2(P_19[10]), .in1(P_18[12]) );
  Fadder_ A_48_557( .carry(c_48_557), .sum(s_48_557), .in3(P_17[14]), .in2(P_16[16]), .in1(P_15[18]) );
  Fadder_ A_48_558( .carry(c_48_558), .sum(s_48_558), .in3(P_14[20]), .in2(P_13[22]), .in1(P_12[24]) );
  Fadder_ A_48_559( .carry(c_48_559), .sum(s_48_559), .in3(P_11[26]), .in2(P_10[28]), .in1(P_9[30]) );
  Fadder_ A_48_560( .carry(c_48_560), .sum(s_48_560), .in3(P_8[32]), .in2(P_7[34]), .in1(P_6[36]) );
  Fadder_ A_48_561( .carry(c_48_561), .sum(s_48_561), .in3(P_5[38]), .in2(P_4[40]), .in1(P_3[42]) );
  Fadder_ A_48_562( .carry(c_48_562), .sum(s_48_562), .in3(P_2[44]), .in2(P_1[46]), .in1(P_0[48]) );
  Fadder_ A_48_563( .carry(c_48_563), .sum(s_48_563), .in3(c_47_538), .in2(c_47_537), .in1(c_47_536) );
  Fadder_ A_48_564( .carry(c_48_564), .sum(s_48_564), .in3(c_47_535), .in2(c_47_534), .in1(c_47_533) );
  Fadder_ A_48_565( .carry(c_48_565), .sum(s_48_565), .in3(c_47_532), .in2(c_47_531), .in1(s_48_554) );
  Fadder_ A_48_566( .carry(c_48_566), .sum(s_48_566), .in3(s_48_562), .in2(s_48_561), .in1(s_48_560) );
  Fadder_ A_48_567( .carry(c_48_567), .sum(s_48_567), .in3(s_48_559), .in2(s_48_558), .in1(s_48_557) );
  Fadder_ A_48_568( .carry(c_48_568), .sum(s_48_568), .in3(s_48_556), .in2(s_48_555), .in1(c_47_539) );
  Fadder_ A_48_569( .carry(c_48_569), .sum(s_48_569), .in3(c_47_541), .in2(c_47_540), .in1(s_48_564) );
  Fadder_ A_48_570( .carry(c_48_570), .sum(s_48_570), .in3(s_48_563), .in2(c_47_543), .in1(c_47_542) );
  Fadder_ A_48_571( .carry(c_48_571), .sum(s_48_571), .in3(s_48_565), .in2(s_48_567), .in1(s_48_566) );
  Fadder_ A_48_572( .carry(c_48_572), .sum(s_48_572), .in3(c_47_544), .in2(s_48_568), .in1(c_47_545) );
  Fadder_ A_48_573( .carry(c_48_573), .sum(s_48_573), .in3(c_47_546), .in2(c_47_547), .in1(s_48_569) );
  Fadder_ A_48_574( .carry(c_48_574), .sum(s_48_574), .in3(s_48_570), .in2(s_48_571), .in1(c_47_548) );
  Fadder_ A_48_575( .carry(c_48_575), .sum(s_48_575), .in3(s_48_572), .in2(c_47_549), .in1(s_48_573) );
  Fadder_ A_48_576( .carry(c_48_576), .sum(s_48_576), .in3(c_47_550), .in2(s_48_574), .in1(c_47_551) );
  Fadder_ A_48_577( .carry(c[48]), .sum(s[48]), .in3(s_48_575), .in2(c_47_552), .in1(s_48_576) );

  // ***** Bit 49 ***** //
  Fadder_ A_49_578( .carry(c_49_578), .sum(s_49_578), .in3(inc[49]), .in2(P_24[1]), .in1(P_23[3]) );
  Fadder_ A_49_579( .carry(c_49_579), .sum(s_49_579), .in3(P_22[5]), .in2(P_21[7]), .in1(P_20[9]) );
  Fadder_ A_49_580( .carry(c_49_580), .sum(s_49_580), .in3(P_19[11]), .in2(P_18[13]), .in1(P_17[15]) );
  Fadder_ A_49_581( .carry(c_49_581), .sum(s_49_581), .in3(P_16[17]), .in2(P_15[19]), .in1(P_14[21]) );
  Fadder_ A_49_582( .carry(c_49_582), .sum(s_49_582), .in3(P_13[23]), .in2(P_12[25]), .in1(P_11[27]) );
  Fadder_ A_49_583( .carry(c_49_583), .sum(s_49_583), .in3(P_10[29]), .in2(P_9[31]), .in1(P_8[33]) );
  Fadder_ A_49_584( .carry(c_49_584), .sum(s_49_584), .in3(P_7[35]), .in2(P_6[37]), .in1(P_5[39]) );
  Fadder_ A_49_585( .carry(c_49_585), .sum(s_49_585), .in3(P_4[41]), .in2(P_3[43]), .in1(P_2[45]) );
  Fadder_ A_49_586( .carry(c_49_586), .sum(s_49_586), .in3(P_1[47]), .in2(P_0[49]), .in1(c_48_554) );
  Fadder_ A_49_587( .carry(c_49_587), .sum(s_49_587), .in3(c_48_562), .in2(c_48_561), .in1(c_48_560) );
  Fadder_ A_49_588( .carry(c_49_588), .sum(s_49_588), .in3(c_48_559), .in2(c_48_558), .in1(c_48_557) );
  Fadder_ A_49_589( .carry(c_49_589), .sum(s_49_589), .in3(c_48_556), .in2(c_48_555), .in1(s_49_585) );
  Fadder_ A_49_590( .carry(c_49_590), .sum(s_49_590), .in3(s_49_584), .in2(s_49_583), .in1(s_49_582) );
  Fadder_ A_49_591( .carry(c_49_591), .sum(s_49_591), .in3(s_49_581), .in2(s_49_580), .in1(s_49_579) );
  Fadder_ A_49_592( .carry(c_49_592), .sum(s_49_592), .in3(s_49_578), .in2(s_49_586), .in1(c_48_564) );
  Fadder_ A_49_593( .carry(c_49_593), .sum(s_49_593), .in3(c_48_563), .in2(c_48_565), .in1(s_49_588) );
  Fadder_ A_49_594( .carry(c_49_594), .sum(s_49_594), .in3(s_49_587), .in2(c_48_567), .in1(c_48_566) );
  Fadder_ A_49_595( .carry(c_49_595), .sum(s_49_595), .in3(s_49_589), .in2(s_49_591), .in1(s_49_590) );
  Fadder_ A_49_596( .carry(c_49_596), .sum(s_49_596), .in3(c_48_568), .in2(c_48_569), .in1(s_49_592) );
  Fadder_ A_49_597( .carry(c_49_597), .sum(s_49_597), .in3(c_48_570), .in2(s_49_593), .in1(s_49_594) );
  Fadder_ A_49_598( .carry(c_49_598), .sum(s_49_598), .in3(c_48_571), .in2(s_49_595), .in1(c_48_572) );
  Fadder_ A_49_599( .carry(c_49_599), .sum(s_49_599), .in3(c_48_573), .in2(s_49_596), .in1(s_49_597) );
  Fadder_ A_49_600( .carry(c_49_600), .sum(s_49_600), .in3(c_48_574), .in2(s_49_598), .in1(c_48_575) );
  Fadder_ A_49_601( .carry(c[49]), .sum(s[49]), .in3(s_49_599), .in2(c_48_576), .in1(s_49_600) );

  // ***** Bit 50 ***** //
  Hadder_ A_50_602( .carry(c_50_602), .sum(s_50_602), .in2(inc[50]), .in1(P_25[0]) );
  Fadder_ A_50_603( .carry(c_50_603), .sum(s_50_603), .in3(P_24[2]), .in2(P_23[4]), .in1(P_22[6]) );
  Fadder_ A_50_604( .carry(c_50_604), .sum(s_50_604), .in3(P_21[8]), .in2(P_20[10]), .in1(P_19[12]) );
  Fadder_ A_50_605( .carry(c_50_605), .sum(s_50_605), .in3(P_18[14]), .in2(P_17[16]), .in1(P_16[18]) );
  Fadder_ A_50_606( .carry(c_50_606), .sum(s_50_606), .in3(P_15[20]), .in2(P_14[22]), .in1(P_13[24]) );
  Fadder_ A_50_607( .carry(c_50_607), .sum(s_50_607), .in3(P_12[26]), .in2(P_11[28]), .in1(P_10[30]) );
  Fadder_ A_50_608( .carry(c_50_608), .sum(s_50_608), .in3(P_9[32]), .in2(P_8[34]), .in1(P_7[36]) );
  Fadder_ A_50_609( .carry(c_50_609), .sum(s_50_609), .in3(P_6[38]), .in2(P_5[40]), .in1(P_4[42]) );
  Fadder_ A_50_610( .carry(c_50_610), .sum(s_50_610), .in3(P_3[44]), .in2(P_2[46]), .in1(P_1[48]) );
  Fadder_ A_50_611( .carry(c_50_611), .sum(s_50_611), .in3(P_0[50]), .in2(c_49_585), .in1(c_49_584) );
  Fadder_ A_50_612( .carry(c_50_612), .sum(s_50_612), .in3(c_49_583), .in2(c_49_582), .in1(c_49_581) );
  Fadder_ A_50_613( .carry(c_50_613), .sum(s_50_613), .in3(c_49_580), .in2(c_49_579), .in1(c_49_578) );
  Fadder_ A_50_614( .carry(c_50_614), .sum(s_50_614), .in3(s_50_602), .in2(s_50_610), .in1(s_50_609) );
  Fadder_ A_50_615( .carry(c_50_615), .sum(s_50_615), .in3(s_50_608), .in2(s_50_607), .in1(s_50_606) );
  Fadder_ A_50_616( .carry(c_50_616), .sum(s_50_616), .in3(s_50_605), .in2(s_50_604), .in1(s_50_603) );
  Fadder_ A_50_617( .carry(c_50_617), .sum(s_50_617), .in3(c_49_586), .in2(c_49_588), .in1(c_49_587) );
  Fadder_ A_50_618( .carry(c_50_618), .sum(s_50_618), .in3(c_49_589), .in2(s_50_611), .in1(s_50_613) );
  Fadder_ A_50_619( .carry(c_50_619), .sum(s_50_619), .in3(s_50_612), .in2(c_49_591), .in1(c_49_590) );
  Fadder_ A_50_620( .carry(c_50_620), .sum(s_50_620), .in3(s_50_614), .in2(s_50_616), .in1(s_50_615) );
  Fadder_ A_50_621( .carry(c_50_621), .sum(s_50_621), .in3(c_49_592), .in2(c_49_593), .in1(s_50_617) );
  Fadder_ A_50_622( .carry(c_50_622), .sum(s_50_622), .in3(c_49_594), .in2(s_50_618), .in1(s_50_619) );
  Fadder_ A_50_623( .carry(c_50_623), .sum(s_50_623), .in3(c_49_595), .in2(s_50_620), .in1(c_49_596) );
  Fadder_ A_50_624( .carry(c_50_624), .sum(s_50_624), .in3(s_50_621), .in2(c_49_597), .in1(s_50_622) );
  Fadder_ A_50_625( .carry(c_50_625), .sum(s_50_625), .in3(c_49_598), .in2(s_50_623), .in1(c_49_599) );
  Fadder_ A_50_626( .carry(c[50]), .sum(s[50]), .in3(s_50_624), .in2(c_49_600), .in1(s_50_625) );

  // ***** Bit 51 ***** //
  Fadder_ A_51_627( .carry(c_51_627), .sum(s_51_627), .in3(inc[51]), .in2(P_25[1]), .in1(P_24[3]) );
  Fadder_ A_51_628( .carry(c_51_628), .sum(s_51_628), .in3(P_23[5]), .in2(P_22[7]), .in1(P_21[9]) );
  Fadder_ A_51_629( .carry(c_51_629), .sum(s_51_629), .in3(P_20[11]), .in2(P_19[13]), .in1(P_18[15]) );
  Fadder_ A_51_630( .carry(c_51_630), .sum(s_51_630), .in3(P_17[17]), .in2(P_16[19]), .in1(P_15[21]) );
  Fadder_ A_51_631( .carry(c_51_631), .sum(s_51_631), .in3(P_14[23]), .in2(P_13[25]), .in1(P_12[27]) );
  Fadder_ A_51_632( .carry(c_51_632), .sum(s_51_632), .in3(P_11[29]), .in2(P_10[31]), .in1(P_9[33]) );
  Fadder_ A_51_633( .carry(c_51_633), .sum(s_51_633), .in3(P_8[35]), .in2(P_7[37]), .in1(P_6[39]) );
  Fadder_ A_51_634( .carry(c_51_634), .sum(s_51_634), .in3(P_5[41]), .in2(P_4[43]), .in1(P_3[45]) );
  Fadder_ A_51_635( .carry(c_51_635), .sum(s_51_635), .in3(P_2[47]), .in2(P_1[49]), .in1(P_0[51]) );
  Fadder_ A_51_636( .carry(c_51_636), .sum(s_51_636), .in3(c_50_602), .in2(c_50_610), .in1(c_50_609) );
  Fadder_ A_51_637( .carry(c_51_637), .sum(s_51_637), .in3(c_50_608), .in2(c_50_607), .in1(c_50_606) );
  Fadder_ A_51_638( .carry(c_51_638), .sum(s_51_638), .in3(c_50_605), .in2(c_50_604), .in1(c_50_603) );
  Fadder_ A_51_639( .carry(c_51_639), .sum(s_51_639), .in3(s_51_635), .in2(s_51_634), .in1(s_51_633) );
  Fadder_ A_51_640( .carry(c_51_640), .sum(s_51_640), .in3(s_51_632), .in2(s_51_631), .in1(s_51_630) );
  Fadder_ A_51_641( .carry(c_51_641), .sum(s_51_641), .in3(s_51_629), .in2(s_51_628), .in1(s_51_627) );
  Fadder_ A_51_642( .carry(c_51_642), .sum(s_51_642), .in3(c_50_613), .in2(c_50_612), .in1(c_50_611) );
  Fadder_ A_51_643( .carry(c_51_643), .sum(s_51_643), .in3(s_51_636), .in2(s_51_638), .in1(s_51_637) );
  Fadder_ A_51_644( .carry(c_51_644), .sum(s_51_644), .in3(c_50_616), .in2(c_50_615), .in1(c_50_614) );
  Fadder_ A_51_645( .carry(c_51_645), .sum(s_51_645), .in3(s_51_641), .in2(s_51_640), .in1(s_51_639) );
  Fadder_ A_51_646( .carry(c_51_646), .sum(s_51_646), .in3(c_50_617), .in2(c_50_618), .in1(s_51_642) );
  Fadder_ A_51_647( .carry(c_51_647), .sum(s_51_647), .in3(c_50_619), .in2(s_51_643), .in1(s_51_644) );
  Fadder_ A_51_648( .carry(c_51_648), .sum(s_51_648), .in3(c_50_620), .in2(s_51_645), .in1(c_50_621) );
  Fadder_ A_51_649( .carry(c_51_649), .sum(s_51_649), .in3(s_51_646), .in2(c_50_622), .in1(s_51_647) );
  Fadder_ A_51_650( .carry(c_51_650), .sum(s_51_650), .in3(c_50_623), .in2(s_51_648), .in1(c_50_624) );
  Fadder_ A_51_651( .carry(c[51]), .sum(s[51]), .in3(s_51_649), .in2(c_50_625), .in1(s_51_650) );

  // ***** Bit 52 ***** //
  Hadder_ A_52_652( .carry(c_52_652), .sum(s_52_652), .in2(inc[52]), .in1(P_26[0]) );
  Fadder_ A_52_653( .carry(c_52_653), .sum(s_52_653), .in3(P_25[2]), .in2(P_24[4]), .in1(P_23[6]) );
  Fadder_ A_52_654( .carry(c_52_654), .sum(s_52_654), .in3(P_22[8]), .in2(P_21[10]), .in1(P_20[12]) );
  Fadder_ A_52_655( .carry(c_52_655), .sum(s_52_655), .in3(P_19[14]), .in2(P_18[16]), .in1(P_17[18]) );
  Fadder_ A_52_656( .carry(c_52_656), .sum(s_52_656), .in3(P_16[20]), .in2(P_15[22]), .in1(P_14[24]) );
  Fadder_ A_52_657( .carry(c_52_657), .sum(s_52_657), .in3(P_13[26]), .in2(P_12[28]), .in1(P_11[30]) );
  Fadder_ A_52_658( .carry(c_52_658), .sum(s_52_658), .in3(P_10[32]), .in2(P_9[34]), .in1(P_8[36]) );
  Fadder_ A_52_659( .carry(c_52_659), .sum(s_52_659), .in3(P_7[38]), .in2(P_6[40]), .in1(P_5[42]) );
  Fadder_ A_52_660( .carry(c_52_660), .sum(s_52_660), .in3(P_4[44]), .in2(P_3[46]), .in1(P_2[48]) );
  Fadder_ A_52_661( .carry(c_52_661), .sum(s_52_661), .in3(P_1[50]), .in2(P_0[52]), .in1(c_51_635) );
  Fadder_ A_52_662( .carry(c_52_662), .sum(s_52_662), .in3(c_51_634), .in2(c_51_633), .in1(c_51_632) );
  Fadder_ A_52_663( .carry(c_52_663), .sum(s_52_663), .in3(c_51_631), .in2(c_51_630), .in1(c_51_629) );
  Fadder_ A_52_664( .carry(c_52_664), .sum(s_52_664), .in3(c_51_628), .in2(c_51_627), .in1(s_52_652) );
  Fadder_ A_52_665( .carry(c_52_665), .sum(s_52_665), .in3(s_52_660), .in2(s_52_659), .in1(s_52_658) );
  Fadder_ A_52_666( .carry(c_52_666), .sum(s_52_666), .in3(s_52_657), .in2(s_52_656), .in1(s_52_655) );
  Fadder_ A_52_667( .carry(c_52_667), .sum(s_52_667), .in3(s_52_654), .in2(s_52_653), .in1(c_51_638) );
  Fadder_ A_52_668( .carry(c_52_668), .sum(s_52_668), .in3(c_51_637), .in2(c_51_636), .in1(s_52_661) );
  Fadder_ A_52_669( .carry(c_52_669), .sum(s_52_669), .in3(s_52_663), .in2(s_52_662), .in1(c_51_641) );
  Fadder_ A_52_670( .carry(c_52_670), .sum(s_52_670), .in3(c_51_640), .in2(c_51_639), .in1(s_52_664) );
  Fadder_ A_52_671( .carry(c_52_671), .sum(s_52_671), .in3(s_52_666), .in2(s_52_665), .in1(c_51_642) );
  Fadder_ A_52_672( .carry(c_52_672), .sum(s_52_672), .in3(s_52_667), .in2(c_51_644), .in1(c_51_643) );
  Fadder_ A_52_673( .carry(c_52_673), .sum(s_52_673), .in3(s_52_668), .in2(s_52_669), .in1(c_51_645) );
  Fadder_ A_52_674( .carry(c_52_674), .sum(s_52_674), .in3(s_52_670), .in2(s_52_671), .in1(c_51_646) );
  Fadder_ A_52_675( .carry(c_52_675), .sum(s_52_675), .in3(s_52_672), .in2(c_51_647), .in1(s_52_673) );
  Fadder_ A_52_676( .carry(c_52_676), .sum(s_52_676), .in3(c_51_648), .in2(s_52_674), .in1(c_51_649) );
  Fadder_ A_52_677( .carry(c[52]), .sum(s[52]), .in3(s_52_675), .in2(c_51_650), .in1(s_52_676) );

  // ***** Bit 53 ***** //
  Fadder_ A_53_678( .carry(c_53_678), .sum(s_53_678), .in3(inc[53]), .in2(P_26[1]), .in1(P_25[3]) );
  Fadder_ A_53_679( .carry(c_53_679), .sum(s_53_679), .in3(P_24[5]), .in2(P_23[7]), .in1(P_22[9]) );
  Fadder_ A_53_680( .carry(c_53_680), .sum(s_53_680), .in3(P_21[11]), .in2(P_20[13]), .in1(P_19[15]) );
  Fadder_ A_53_681( .carry(c_53_681), .sum(s_53_681), .in3(P_18[17]), .in2(P_17[19]), .in1(P_16[21]) );
  Fadder_ A_53_682( .carry(c_53_682), .sum(s_53_682), .in3(P_15[23]), .in2(P_14[25]), .in1(P_13[27]) );
  Fadder_ A_53_683( .carry(c_53_683), .sum(s_53_683), .in3(P_12[29]), .in2(P_11[31]), .in1(P_10[33]) );
  Fadder_ A_53_684( .carry(c_53_684), .sum(s_53_684), .in3(P_9[35]), .in2(P_8[37]), .in1(P_7[39]) );
  Fadder_ A_53_685( .carry(c_53_685), .sum(s_53_685), .in3(P_6[41]), .in2(P_5[43]), .in1(P_4[45]) );
  Fadder_ A_53_686( .carry(c_53_686), .sum(s_53_686), .in3(P_3[47]), .in2(P_2[49]), .in1(P_1[51]) );
  Fadder_ A_53_687( .carry(c_53_687), .sum(s_53_687), .in3(P_0[53]), .in2(c_52_652), .in1(c_52_660) );
  Fadder_ A_53_688( .carry(c_53_688), .sum(s_53_688), .in3(c_52_659), .in2(c_52_658), .in1(c_52_657) );
  Fadder_ A_53_689( .carry(c_53_689), .sum(s_53_689), .in3(c_52_656), .in2(c_52_655), .in1(c_52_654) );
  Fadder_ A_53_690( .carry(c_53_690), .sum(s_53_690), .in3(c_52_653), .in2(s_53_686), .in1(s_53_685) );
  Fadder_ A_53_691( .carry(c_53_691), .sum(s_53_691), .in3(s_53_684), .in2(s_53_683), .in1(s_53_682) );
  Fadder_ A_53_692( .carry(c_53_692), .sum(s_53_692), .in3(s_53_681), .in2(s_53_680), .in1(s_53_679) );
  Fadder_ A_53_693( .carry(c_53_693), .sum(s_53_693), .in3(s_53_678), .in2(c_52_661), .in1(c_52_663) );
  Fadder_ A_53_694( .carry(c_53_694), .sum(s_53_694), .in3(c_52_662), .in2(c_52_664), .in1(s_53_687) );
  Fadder_ A_53_695( .carry(c_53_695), .sum(s_53_695), .in3(s_53_689), .in2(s_53_688), .in1(c_52_666) );
  Fadder_ A_53_696( .carry(c_53_696), .sum(s_53_696), .in3(c_52_665), .in2(s_53_690), .in1(s_53_692) );
  Fadder_ A_53_697( .carry(c_53_697), .sum(s_53_697), .in3(s_53_691), .in2(c_52_667), .in1(c_52_668) );
  Fadder_ A_53_698( .carry(c_53_698), .sum(s_53_698), .in3(s_53_693), .in2(c_52_670), .in1(c_52_669) );
  Fadder_ A_53_699( .carry(c_53_699), .sum(s_53_699), .in3(s_53_694), .in2(s_53_695), .in1(s_53_696) );
  Fadder_ A_53_700( .carry(c_53_700), .sum(s_53_700), .in3(c_52_671), .in2(s_53_697), .in1(c_52_672) );
  Fadder_ A_53_701( .carry(c_53_701), .sum(s_53_701), .in3(s_53_698), .in2(c_52_673), .in1(s_53_699) );
  Fadder_ A_53_702( .carry(c_53_702), .sum(s_53_702), .in3(c_52_674), .in2(s_53_700), .in1(c_52_675) );
  Fadder_ A_53_703( .carry(c[53]), .sum(s[53]), .in3(s_53_701), .in2(c_52_676), .in1(s_53_702) );

  // ***** Bit 54 ***** //
  Hadder_ A_54_704( .carry(c_54_704), .sum(s_54_704), .in2(inc[54]), .in1(P_27[0]) );
  Fadder_ A_54_705( .carry(c_54_705), .sum(s_54_705), .in3(P_26[2]), .in2(P_25[4]), .in1(P_24[6]) );
  Fadder_ A_54_706( .carry(c_54_706), .sum(s_54_706), .in3(P_23[8]), .in2(P_22[10]), .in1(P_21[12]) );
  Fadder_ A_54_707( .carry(c_54_707), .sum(s_54_707), .in3(P_20[14]), .in2(P_19[16]), .in1(P_18[18]) );
  Fadder_ A_54_708( .carry(c_54_708), .sum(s_54_708), .in3(P_17[20]), .in2(P_16[22]), .in1(P_15[24]) );
  Fadder_ A_54_709( .carry(c_54_709), .sum(s_54_709), .in3(P_14[26]), .in2(P_13[28]), .in1(P_12[30]) );
  Fadder_ A_54_710( .carry(c_54_710), .sum(s_54_710), .in3(P_11[32]), .in2(P_10[34]), .in1(P_9[36]) );
  Fadder_ A_54_711( .carry(c_54_711), .sum(s_54_711), .in3(P_8[38]), .in2(P_7[40]), .in1(P_6[42]) );
  Fadder_ A_54_712( .carry(c_54_712), .sum(s_54_712), .in3(P_5[44]), .in2(P_4[46]), .in1(P_3[48]) );
  Fadder_ A_54_713( .carry(c_54_713), .sum(s_54_713), .in3(P_2[50]), .in2(P_1[52]), .in1(P_0[54]) );
  Fadder_ A_54_714( .carry(c_54_714), .sum(s_54_714), .in3(c_53_686), .in2(c_53_685), .in1(c_53_684) );
  Fadder_ A_54_715( .carry(c_54_715), .sum(s_54_715), .in3(c_53_683), .in2(c_53_682), .in1(c_53_681) );
  Fadder_ A_54_716( .carry(c_54_716), .sum(s_54_716), .in3(c_53_680), .in2(c_53_679), .in1(c_53_678) );
  Fadder_ A_54_717( .carry(c_54_717), .sum(s_54_717), .in3(s_54_704), .in2(s_54_713), .in1(s_54_712) );
  Fadder_ A_54_718( .carry(c_54_718), .sum(s_54_718), .in3(s_54_711), .in2(s_54_710), .in1(s_54_709) );
  Fadder_ A_54_719( .carry(c_54_719), .sum(s_54_719), .in3(s_54_708), .in2(s_54_707), .in1(s_54_706) );
  Fadder_ A_54_720( .carry(c_54_720), .sum(s_54_720), .in3(s_54_705), .in2(c_53_687), .in1(c_53_689) );
  Fadder_ A_54_721( .carry(c_54_721), .sum(s_54_721), .in3(c_53_688), .in2(s_54_716), .in1(s_54_715) );
  Fadder_ A_54_722( .carry(c_54_722), .sum(s_54_722), .in3(s_54_714), .in2(c_53_692), .in1(c_53_691) );
  Fadder_ A_54_723( .carry(c_54_723), .sum(s_54_723), .in3(c_53_690), .in2(s_54_717), .in1(s_54_719) );
  Fadder_ A_54_724( .carry(c_54_724), .sum(s_54_724), .in3(s_54_718), .in2(c_53_693), .in1(c_53_694) );
  Fadder_ A_54_725( .carry(c_54_725), .sum(s_54_725), .in3(s_54_720), .in2(c_53_695), .in1(s_54_721) );
  Fadder_ A_54_726( .carry(c_54_726), .sum(s_54_726), .in3(c_53_696), .in2(s_54_722), .in1(s_54_723) );
  Fadder_ A_54_727( .carry(c_54_727), .sum(s_54_727), .in3(c_53_697), .in2(s_54_724), .in1(c_53_698) );
  Fadder_ A_54_728( .carry(c_54_728), .sum(s_54_728), .in3(c_53_699), .in2(s_54_725), .in1(s_54_726) );
  Fadder_ A_54_729( .carry(c_54_729), .sum(s_54_729), .in3(c_53_700), .in2(s_54_727), .in1(c_53_701) );
  Fadder_ A_54_730( .carry(c[54]), .sum(s[54]), .in3(s_54_728), .in2(c_53_702), .in1(s_54_729) );

  // ***** Bit 55 ***** //
  Fadder_ A_55_731( .carry(c_55_731), .sum(s_55_731), .in3(inc[55]), .in2(P_27[1]), .in1(P_26[3]) );
  Fadder_ A_55_732( .carry(c_55_732), .sum(s_55_732), .in3(P_25[5]), .in2(P_24[7]), .in1(P_23[9]) );
  Fadder_ A_55_733( .carry(c_55_733), .sum(s_55_733), .in3(P_22[11]), .in2(P_21[13]), .in1(P_20[15]) );
  Fadder_ A_55_734( .carry(c_55_734), .sum(s_55_734), .in3(P_19[17]), .in2(P_18[19]), .in1(P_17[21]) );
  Fadder_ A_55_735( .carry(c_55_735), .sum(s_55_735), .in3(P_16[23]), .in2(P_15[25]), .in1(P_14[27]) );
  Fadder_ A_55_736( .carry(c_55_736), .sum(s_55_736), .in3(P_13[29]), .in2(P_12[31]), .in1(P_11[33]) );
  Fadder_ A_55_737( .carry(c_55_737), .sum(s_55_737), .in3(P_10[35]), .in2(P_9[37]), .in1(P_8[39]) );
  Fadder_ A_55_738( .carry(c_55_738), .sum(s_55_738), .in3(P_7[41]), .in2(P_6[43]), .in1(P_5[45]) );
  Fadder_ A_55_739( .carry(c_55_739), .sum(s_55_739), .in3(P_4[47]), .in2(P_3[49]), .in1(P_2[51]) );
  Fadder_ A_55_740( .carry(c_55_740), .sum(s_55_740), .in3(P_1[53]), .in2(P_0[55]), .in1(c_54_704) );
  Fadder_ A_55_741( .carry(c_55_741), .sum(s_55_741), .in3(c_54_713), .in2(c_54_712), .in1(c_54_711) );
  Fadder_ A_55_742( .carry(c_55_742), .sum(s_55_742), .in3(c_54_710), .in2(c_54_709), .in1(c_54_708) );
  Fadder_ A_55_743( .carry(c_55_743), .sum(s_55_743), .in3(c_54_707), .in2(c_54_706), .in1(c_54_705) );
  Fadder_ A_55_744( .carry(c_55_744), .sum(s_55_744), .in3(s_55_739), .in2(s_55_738), .in1(s_55_737) );
  Fadder_ A_55_745( .carry(c_55_745), .sum(s_55_745), .in3(s_55_736), .in2(s_55_735), .in1(s_55_734) );
  Fadder_ A_55_746( .carry(c_55_746), .sum(s_55_746), .in3(s_55_733), .in2(s_55_732), .in1(s_55_731) );
  Fadder_ A_55_747( .carry(c_55_747), .sum(s_55_747), .in3(s_55_740), .in2(c_54_716), .in1(c_54_715) );
  Fadder_ A_55_748( .carry(c_55_748), .sum(s_55_748), .in3(c_54_714), .in2(s_55_743), .in1(s_55_742) );
  Fadder_ A_55_749( .carry(c_55_749), .sum(s_55_749), .in3(s_55_741), .in2(c_54_719), .in1(c_54_718) );
  Fadder_ A_55_750( .carry(c_55_750), .sum(s_55_750), .in3(c_54_717), .in2(s_55_746), .in1(s_55_745) );
  Fadder_ A_55_751( .carry(c_55_751), .sum(s_55_751), .in3(s_55_744), .in2(c_54_720), .in1(s_55_747) );
  Fadder_ A_55_752( .carry(c_55_752), .sum(s_55_752), .in3(c_54_722), .in2(c_54_721), .in1(s_55_748) );
  Fadder_ A_55_753( .carry(c_55_753), .sum(s_55_753), .in3(c_54_723), .in2(s_55_749), .in1(s_55_750) );
  Fadder_ A_55_754( .carry(c_55_754), .sum(s_55_754), .in3(c_54_724), .in2(c_54_725), .in1(s_55_751) );
  Fadder_ A_55_755( .carry(c_55_755), .sum(s_55_755), .in3(c_54_726), .in2(s_55_752), .in1(s_55_753) );
  Fadder_ A_55_756( .carry(c_55_756), .sum(s_55_756), .in3(c_54_727), .in2(s_55_754), .in1(c_54_728) );
  Fadder_ A_55_757( .carry(c[55]), .sum(s[55]), .in3(s_55_755), .in2(c_54_729), .in1(s_55_756) );

  // ***** Bit 56 ***** //
  Hadder_ A_56_758( .carry(c_56_758), .sum(s_56_758), .in2(inc[56]), .in1(P_28[0]) );
  Fadder_ A_56_759( .carry(c_56_759), .sum(s_56_759), .in3(P_27[2]), .in2(P_26[4]), .in1(P_25[6]) );
  Fadder_ A_56_760( .carry(c_56_760), .sum(s_56_760), .in3(P_24[8]), .in2(P_23[10]), .in1(P_22[12]) );
  Fadder_ A_56_761( .carry(c_56_761), .sum(s_56_761), .in3(P_21[14]), .in2(P_20[16]), .in1(P_19[18]) );
  Fadder_ A_56_762( .carry(c_56_762), .sum(s_56_762), .in3(P_18[20]), .in2(P_17[22]), .in1(P_16[24]) );
  Fadder_ A_56_763( .carry(c_56_763), .sum(s_56_763), .in3(P_15[26]), .in2(P_14[28]), .in1(P_13[30]) );
  Fadder_ A_56_764( .carry(c_56_764), .sum(s_56_764), .in3(P_12[32]), .in2(P_11[34]), .in1(P_10[36]) );
  Fadder_ A_56_765( .carry(c_56_765), .sum(s_56_765), .in3(P_9[38]), .in2(P_8[40]), .in1(P_7[42]) );
  Fadder_ A_56_766( .carry(c_56_766), .sum(s_56_766), .in3(P_6[44]), .in2(P_5[46]), .in1(P_4[48]) );
  Fadder_ A_56_767( .carry(c_56_767), .sum(s_56_767), .in3(P_3[50]), .in2(P_2[52]), .in1(P_1[54]) );
  Fadder_ A_56_768( .carry(c_56_768), .sum(s_56_768), .in3(P_0[56]), .in2(c_55_739), .in1(c_55_738) );
  Fadder_ A_56_769( .carry(c_56_769), .sum(s_56_769), .in3(c_55_737), .in2(c_55_736), .in1(c_55_735) );
  Fadder_ A_56_770( .carry(c_56_770), .sum(s_56_770), .in3(c_55_734), .in2(c_55_733), .in1(c_55_732) );
  Fadder_ A_56_771( .carry(c_56_771), .sum(s_56_771), .in3(c_55_731), .in2(s_56_758), .in1(s_56_767) );
  Fadder_ A_56_772( .carry(c_56_772), .sum(s_56_772), .in3(s_56_766), .in2(s_56_765), .in1(s_56_764) );
  Fadder_ A_56_773( .carry(c_56_773), .sum(s_56_773), .in3(s_56_763), .in2(s_56_762), .in1(s_56_761) );
  Fadder_ A_56_774( .carry(c_56_774), .sum(s_56_774), .in3(s_56_760), .in2(s_56_759), .in1(c_55_740) );
  Fadder_ A_56_775( .carry(c_56_775), .sum(s_56_775), .in3(c_55_743), .in2(c_55_742), .in1(c_55_741) );
  Fadder_ A_56_776( .carry(c_56_776), .sum(s_56_776), .in3(s_56_768), .in2(s_56_770), .in1(s_56_769) );
  Fadder_ A_56_777( .carry(c_56_777), .sum(s_56_777), .in3(c_55_746), .in2(c_55_745), .in1(c_55_744) );
  Fadder_ A_56_778( .carry(c_56_778), .sum(s_56_778), .in3(s_56_771), .in2(s_56_773), .in1(s_56_772) );
  Fadder_ A_56_779( .carry(c_56_779), .sum(s_56_779), .in3(s_56_774), .in2(c_55_747), .in1(s_56_775) );
  Fadder_ A_56_780( .carry(c_56_780), .sum(s_56_780), .in3(c_55_749), .in2(c_55_748), .in1(s_56_776) );
  Fadder_ A_56_781( .carry(c_56_781), .sum(s_56_781), .in3(s_56_777), .in2(c_55_750), .in1(s_56_778) );
  Fadder_ A_56_782( .carry(c_56_782), .sum(s_56_782), .in3(c_55_751), .in2(c_55_752), .in1(s_56_779) );
  Fadder_ A_56_783( .carry(c_56_783), .sum(s_56_783), .in3(c_55_753), .in2(s_56_780), .in1(s_56_781) );
  Fadder_ A_56_784( .carry(c_56_784), .sum(s_56_784), .in3(c_55_754), .in2(s_56_782), .in1(c_55_755) );
  Fadder_ A_56_785( .carry(c[56]), .sum(s[56]), .in3(s_56_783), .in2(c_55_756), .in1(s_56_784) );

  // ***** Bit 57 ***** //
  Fadder_ A_57_786( .carry(c_57_786), .sum(s_57_786), .in3(inc[57]), .in2(P_28[1]), .in1(P_27[3]) );
  Fadder_ A_57_787( .carry(c_57_787), .sum(s_57_787), .in3(P_26[5]), .in2(P_25[7]), .in1(P_24[9]) );
  Fadder_ A_57_788( .carry(c_57_788), .sum(s_57_788), .in3(P_23[11]), .in2(P_22[13]), .in1(P_21[15]) );
  Fadder_ A_57_789( .carry(c_57_789), .sum(s_57_789), .in3(P_20[17]), .in2(P_19[19]), .in1(P_18[21]) );
  Fadder_ A_57_790( .carry(c_57_790), .sum(s_57_790), .in3(P_17[23]), .in2(P_16[25]), .in1(P_15[27]) );
  Fadder_ A_57_791( .carry(c_57_791), .sum(s_57_791), .in3(P_14[29]), .in2(P_13[31]), .in1(P_12[33]) );
  Fadder_ A_57_792( .carry(c_57_792), .sum(s_57_792), .in3(P_11[35]), .in2(P_10[37]), .in1(P_9[39]) );
  Fadder_ A_57_793( .carry(c_57_793), .sum(s_57_793), .in3(P_8[41]), .in2(P_7[43]), .in1(P_6[45]) );
  Fadder_ A_57_794( .carry(c_57_794), .sum(s_57_794), .in3(P_5[47]), .in2(P_4[49]), .in1(P_3[51]) );
  Fadder_ A_57_795( .carry(c_57_795), .sum(s_57_795), .in3(P_2[53]), .in2(P_1[55]), .in1(P_0[57]) );
  Fadder_ A_57_796( .carry(c_57_796), .sum(s_57_796), .in3(c_56_758), .in2(c_56_767), .in1(c_56_766) );
  Fadder_ A_57_797( .carry(c_57_797), .sum(s_57_797), .in3(c_56_765), .in2(c_56_764), .in1(c_56_763) );
  Fadder_ A_57_798( .carry(c_57_798), .sum(s_57_798), .in3(c_56_762), .in2(c_56_761), .in1(c_56_760) );
  Fadder_ A_57_799( .carry(c_57_799), .sum(s_57_799), .in3(c_56_759), .in2(s_57_795), .in1(s_57_794) );
  Fadder_ A_57_800( .carry(c_57_800), .sum(s_57_800), .in3(s_57_793), .in2(s_57_792), .in1(s_57_791) );
  Fadder_ A_57_801( .carry(c_57_801), .sum(s_57_801), .in3(s_57_790), .in2(s_57_789), .in1(s_57_788) );
  Fadder_ A_57_802( .carry(c_57_802), .sum(s_57_802), .in3(s_57_787), .in2(s_57_786), .in1(c_56_770) );
  Fadder_ A_57_803( .carry(c_57_803), .sum(s_57_803), .in3(c_56_769), .in2(c_56_768), .in1(s_57_796) );
  Fadder_ A_57_804( .carry(c_57_804), .sum(s_57_804), .in3(c_56_771), .in2(s_57_798), .in1(s_57_797) );
  Fadder_ A_57_805( .carry(c_57_805), .sum(s_57_805), .in3(c_56_773), .in2(c_56_772), .in1(c_56_774) );
  Fadder_ A_57_806( .carry(c_57_806), .sum(s_57_806), .in3(s_57_799), .in2(s_57_801), .in1(s_57_800) );
  Fadder_ A_57_807( .carry(c_57_807), .sum(s_57_807), .in3(c_56_775), .in2(s_57_802), .in1(c_56_777) );
  Fadder_ A_57_808( .carry(c_57_808), .sum(s_57_808), .in3(c_56_776), .in2(s_57_803), .in1(s_57_804) );
  Fadder_ A_57_809( .carry(c_57_809), .sum(s_57_809), .in3(s_57_805), .in2(c_56_778), .in1(s_57_806) );
  Fadder_ A_57_810( .carry(c_57_810), .sum(s_57_810), .in3(c_56_779), .in2(c_56_780), .in1(s_57_807) );
  Fadder_ A_57_811( .carry(c_57_811), .sum(s_57_811), .in3(c_56_781), .in2(s_57_808), .in1(s_57_809) );
  Fadder_ A_57_812( .carry(c_57_812), .sum(s_57_812), .in3(c_56_782), .in2(s_57_810), .in1(c_56_783) );
  Fadder_ A_57_813( .carry(c[57]), .sum(s[57]), .in3(s_57_811), .in2(c_56_784), .in1(s_57_812) );

  // ***** Bit 58 ***** //
  Hadder_ A_58_814( .carry(c_58_814), .sum(s_58_814), .in2(inc[58]), .in1(P_29[0]) );
  Fadder_ A_58_815( .carry(c_58_815), .sum(s_58_815), .in3(P_28[2]), .in2(P_27[4]), .in1(P_26[6]) );
  Fadder_ A_58_816( .carry(c_58_816), .sum(s_58_816), .in3(P_25[8]), .in2(P_24[10]), .in1(P_23[12]) );
  Fadder_ A_58_817( .carry(c_58_817), .sum(s_58_817), .in3(P_22[14]), .in2(P_21[16]), .in1(P_20[18]) );
  Fadder_ A_58_818( .carry(c_58_818), .sum(s_58_818), .in3(P_19[20]), .in2(P_18[22]), .in1(P_17[24]) );
  Fadder_ A_58_819( .carry(c_58_819), .sum(s_58_819), .in3(P_16[26]), .in2(P_15[28]), .in1(P_14[30]) );
  Fadder_ A_58_820( .carry(c_58_820), .sum(s_58_820), .in3(P_13[32]), .in2(P_12[34]), .in1(P_11[36]) );
  Fadder_ A_58_821( .carry(c_58_821), .sum(s_58_821), .in3(P_10[38]), .in2(P_9[40]), .in1(P_8[42]) );
  Fadder_ A_58_822( .carry(c_58_822), .sum(s_58_822), .in3(P_7[44]), .in2(P_6[46]), .in1(P_5[48]) );
  Fadder_ A_58_823( .carry(c_58_823), .sum(s_58_823), .in3(P_4[50]), .in2(P_3[52]), .in1(P_2[54]) );
  Fadder_ A_58_824( .carry(c_58_824), .sum(s_58_824), .in3(P_1[56]), .in2(P_0[58]), .in1(c_57_795) );
  Fadder_ A_58_825( .carry(c_58_825), .sum(s_58_825), .in3(c_57_794), .in2(c_57_793), .in1(c_57_792) );
  Fadder_ A_58_826( .carry(c_58_826), .sum(s_58_826), .in3(c_57_791), .in2(c_57_790), .in1(c_57_789) );
  Fadder_ A_58_827( .carry(c_58_827), .sum(s_58_827), .in3(c_57_788), .in2(c_57_787), .in1(c_57_786) );
  Fadder_ A_58_828( .carry(c_58_828), .sum(s_58_828), .in3(s_58_814), .in2(s_58_823), .in1(s_58_822) );
  Fadder_ A_58_829( .carry(c_58_829), .sum(s_58_829), .in3(s_58_821), .in2(s_58_820), .in1(s_58_819) );
  Fadder_ A_58_830( .carry(c_58_830), .sum(s_58_830), .in3(s_58_818), .in2(s_58_817), .in1(s_58_816) );
  Fadder_ A_58_831( .carry(c_58_831), .sum(s_58_831), .in3(s_58_815), .in2(c_57_798), .in1(c_57_797) );
  Fadder_ A_58_832( .carry(c_58_832), .sum(s_58_832), .in3(c_57_796), .in2(s_58_824), .in1(s_58_827) );
  Fadder_ A_58_833( .carry(c_58_833), .sum(s_58_833), .in3(s_58_826), .in2(s_58_825), .in1(c_57_801) );
  Fadder_ A_58_834( .carry(c_58_834), .sum(s_58_834), .in3(c_57_800), .in2(c_57_799), .in1(s_58_828) );
  Fadder_ A_58_835( .carry(c_58_835), .sum(s_58_835), .in3(s_58_830), .in2(s_58_829), .in1(c_57_802) );
  Fadder_ A_58_836( .carry(c_58_836), .sum(s_58_836), .in3(c_57_803), .in2(s_58_831), .in1(c_57_805) );
  Fadder_ A_58_837( .carry(c_58_837), .sum(s_58_837), .in3(c_57_804), .in2(s_58_832), .in1(s_58_833) );
  Fadder_ A_58_838( .carry(c_58_838), .sum(s_58_838), .in3(c_57_806), .in2(s_58_834), .in1(s_58_835) );
  Fadder_ A_58_839( .carry(c_58_839), .sum(s_58_839), .in3(c_57_807), .in2(c_57_808), .in1(s_58_836) );
  Fadder_ A_58_840( .carry(c_58_840), .sum(s_58_840), .in3(c_57_809), .in2(s_58_837), .in1(s_58_838) );
  Fadder_ A_58_841( .carry(c_58_841), .sum(s_58_841), .in3(c_57_810), .in2(s_58_839), .in1(c_57_811) );
  Fadder_ A_58_842( .carry(c[58]), .sum(s[58]), .in3(s_58_840), .in2(c_57_812), .in1(s_58_841) );

  // ***** Bit 59 ***** //
  Fadder_ A_59_843( .carry(c_59_843), .sum(s_59_843), .in3(inc[59]), .in2(P_29[1]), .in1(P_28[3]) );
  Fadder_ A_59_844( .carry(c_59_844), .sum(s_59_844), .in3(P_27[5]), .in2(P_26[7]), .in1(P_25[9]) );
  Fadder_ A_59_845( .carry(c_59_845), .sum(s_59_845), .in3(P_24[11]), .in2(P_23[13]), .in1(P_22[15]) );
  Fadder_ A_59_846( .carry(c_59_846), .sum(s_59_846), .in3(P_21[17]), .in2(P_20[19]), .in1(P_19[21]) );
  Fadder_ A_59_847( .carry(c_59_847), .sum(s_59_847), .in3(P_18[23]), .in2(P_17[25]), .in1(P_16[27]) );
  Fadder_ A_59_848( .carry(c_59_848), .sum(s_59_848), .in3(P_15[29]), .in2(P_14[31]), .in1(P_13[33]) );
  Fadder_ A_59_849( .carry(c_59_849), .sum(s_59_849), .in3(P_12[35]), .in2(P_11[37]), .in1(P_10[39]) );
  Fadder_ A_59_850( .carry(c_59_850), .sum(s_59_850), .in3(P_9[41]), .in2(P_8[43]), .in1(P_7[45]) );
  Fadder_ A_59_851( .carry(c_59_851), .sum(s_59_851), .in3(P_6[47]), .in2(P_5[49]), .in1(P_4[51]) );
  Fadder_ A_59_852( .carry(c_59_852), .sum(s_59_852), .in3(P_3[53]), .in2(P_2[55]), .in1(P_1[57]) );
  Fadder_ A_59_853( .carry(c_59_853), .sum(s_59_853), .in3(P_0[59]), .in2(c_58_814), .in1(c_58_823) );
  Fadder_ A_59_854( .carry(c_59_854), .sum(s_59_854), .in3(c_58_822), .in2(c_58_821), .in1(c_58_820) );
  Fadder_ A_59_855( .carry(c_59_855), .sum(s_59_855), .in3(c_58_819), .in2(c_58_818), .in1(c_58_817) );
  Fadder_ A_59_856( .carry(c_59_856), .sum(s_59_856), .in3(c_58_816), .in2(c_58_815), .in1(s_59_852) );
  Fadder_ A_59_857( .carry(c_59_857), .sum(s_59_857), .in3(s_59_851), .in2(s_59_850), .in1(s_59_849) );
  Fadder_ A_59_858( .carry(c_59_858), .sum(s_59_858), .in3(s_59_848), .in2(s_59_847), .in1(s_59_846) );
  Fadder_ A_59_859( .carry(c_59_859), .sum(s_59_859), .in3(s_59_845), .in2(s_59_844), .in1(s_59_843) );
  Fadder_ A_59_860( .carry(c_59_860), .sum(s_59_860), .in3(c_58_824), .in2(c_58_827), .in1(c_58_826) );
  Fadder_ A_59_861( .carry(c_59_861), .sum(s_59_861), .in3(c_58_825), .in2(s_59_853), .in1(s_59_855) );
  Fadder_ A_59_862( .carry(c_59_862), .sum(s_59_862), .in3(s_59_854), .in2(c_58_830), .in1(c_58_829) );
  Fadder_ A_59_863( .carry(c_59_863), .sum(s_59_863), .in3(c_58_828), .in2(s_59_856), .in1(s_59_859) );
  Fadder_ A_59_864( .carry(c_59_864), .sum(s_59_864), .in3(s_59_858), .in2(s_59_857), .in1(c_58_831) );
  Fadder_ A_59_865( .carry(c_59_865), .sum(s_59_865), .in3(s_59_860), .in2(c_58_832), .in1(c_58_833) );
  Fadder_ A_59_866( .carry(c_59_866), .sum(s_59_866), .in3(c_58_834), .in2(s_59_861), .in1(s_59_862) );
  Fadder_ A_59_867( .carry(c_59_867), .sum(s_59_867), .in3(s_59_863), .in2(c_58_835), .in1(s_59_864) );
  Fadder_ A_59_868( .carry(c_59_868), .sum(s_59_868), .in3(c_58_836), .in2(s_59_865), .in1(c_58_837) );
  Fadder_ A_59_869( .carry(c_59_869), .sum(s_59_869), .in3(s_59_866), .in2(c_58_838), .in1(s_59_867) );
  Fadder_ A_59_870( .carry(c_59_870), .sum(s_59_870), .in3(c_58_839), .in2(s_59_868), .in1(c_58_840) );
  Fadder_ A_59_871( .carry(c[59]), .sum(s[59]), .in3(s_59_869), .in2(c_58_841), .in1(s_59_870) );

  // ***** Bit 60 ***** //
  Hadder_ A_60_872( .carry(c_60_872), .sum(s_60_872), .in2(inc[60]), .in1(P_30[0]) );
  Fadder_ A_60_873( .carry(c_60_873), .sum(s_60_873), .in3(P_29[2]), .in2(P_28[4]), .in1(P_27[6]) );
  Fadder_ A_60_874( .carry(c_60_874), .sum(s_60_874), .in3(P_26[8]), .in2(P_25[10]), .in1(P_24[12]) );
  Fadder_ A_60_875( .carry(c_60_875), .sum(s_60_875), .in3(P_23[14]), .in2(P_22[16]), .in1(P_21[18]) );
  Fadder_ A_60_876( .carry(c_60_876), .sum(s_60_876), .in3(P_20[20]), .in2(P_19[22]), .in1(P_18[24]) );
  Fadder_ A_60_877( .carry(c_60_877), .sum(s_60_877), .in3(P_17[26]), .in2(P_16[28]), .in1(P_15[30]) );
  Fadder_ A_60_878( .carry(c_60_878), .sum(s_60_878), .in3(P_14[32]), .in2(P_13[34]), .in1(P_12[36]) );
  Fadder_ A_60_879( .carry(c_60_879), .sum(s_60_879), .in3(P_11[38]), .in2(P_10[40]), .in1(P_9[42]) );
  Fadder_ A_60_880( .carry(c_60_880), .sum(s_60_880), .in3(P_8[44]), .in2(P_7[46]), .in1(P_6[48]) );
  Fadder_ A_60_881( .carry(c_60_881), .sum(s_60_881), .in3(P_5[50]), .in2(P_4[52]), .in1(P_3[54]) );
  Fadder_ A_60_882( .carry(c_60_882), .sum(s_60_882), .in3(P_2[56]), .in2(P_1[58]), .in1(P_0[60]) );
  Fadder_ A_60_883( .carry(c_60_883), .sum(s_60_883), .in3(c_59_852), .in2(c_59_851), .in1(c_59_850) );
  Fadder_ A_60_884( .carry(c_60_884), .sum(s_60_884), .in3(c_59_849), .in2(c_59_848), .in1(c_59_847) );
  Fadder_ A_60_885( .carry(c_60_885), .sum(s_60_885), .in3(c_59_846), .in2(c_59_845), .in1(c_59_844) );
  Fadder_ A_60_886( .carry(c_60_886), .sum(s_60_886), .in3(c_59_843), .in2(s_60_872), .in1(s_60_882) );
  Fadder_ A_60_887( .carry(c_60_887), .sum(s_60_887), .in3(s_60_881), .in2(s_60_880), .in1(s_60_879) );
  Fadder_ A_60_888( .carry(c_60_888), .sum(s_60_888), .in3(s_60_878), .in2(s_60_877), .in1(s_60_876) );
  Fadder_ A_60_889( .carry(c_60_889), .sum(s_60_889), .in3(s_60_875), .in2(s_60_874), .in1(s_60_873) );
  Fadder_ A_60_890( .carry(c_60_890), .sum(s_60_890), .in3(c_59_853), .in2(c_59_855), .in1(c_59_854) );
  Fadder_ A_60_891( .carry(c_60_891), .sum(s_60_891), .in3(c_59_856), .in2(s_60_885), .in1(s_60_884) );
  Fadder_ A_60_892( .carry(c_60_892), .sum(s_60_892), .in3(s_60_883), .in2(c_59_859), .in1(c_59_858) );
  Fadder_ A_60_893( .carry(c_60_893), .sum(s_60_893), .in3(c_59_857), .in2(s_60_886), .in1(s_60_889) );
  Fadder_ A_60_894( .carry(c_60_894), .sum(s_60_894), .in3(s_60_888), .in2(s_60_887), .in1(c_59_860) );
  Fadder_ A_60_895( .carry(c_60_895), .sum(s_60_895), .in3(s_60_890), .in2(c_59_861), .in1(c_59_862) );
  Fadder_ A_60_896( .carry(c_60_896), .sum(s_60_896), .in3(s_60_891), .in2(c_59_863), .in1(s_60_892) );
  Fadder_ A_60_897( .carry(c_60_897), .sum(s_60_897), .in3(s_60_893), .in2(c_59_864), .in1(s_60_894) );
  Fadder_ A_60_898( .carry(c_60_898), .sum(s_60_898), .in3(c_59_865), .in2(s_60_895), .in1(c_59_866) );
  Fadder_ A_60_899( .carry(c_60_899), .sum(s_60_899), .in3(s_60_896), .in2(c_59_867), .in1(s_60_897) );
  Fadder_ A_60_900( .carry(c_60_900), .sum(s_60_900), .in3(c_59_868), .in2(s_60_898), .in1(c_59_869) );
  Fadder_ A_60_901( .carry(c[60]), .sum(s[60]), .in3(s_60_899), .in2(c_59_870), .in1(s_60_900) );

  // ***** Bit 61 ***** //
  Fadder_ A_61_902( .carry(c_61_902), .sum(s_61_902), .in3(inc[61]), .in2(P_30[1]), .in1(P_29[3]) );
  Fadder_ A_61_903( .carry(c_61_903), .sum(s_61_903), .in3(P_28[5]), .in2(P_27[7]), .in1(P_26[9]) );
  Fadder_ A_61_904( .carry(c_61_904), .sum(s_61_904), .in3(P_25[11]), .in2(P_24[13]), .in1(P_23[15]) );
  Fadder_ A_61_905( .carry(c_61_905), .sum(s_61_905), .in3(P_22[17]), .in2(P_21[19]), .in1(P_20[21]) );
  Fadder_ A_61_906( .carry(c_61_906), .sum(s_61_906), .in3(P_19[23]), .in2(P_18[25]), .in1(P_17[27]) );
  Fadder_ A_61_907( .carry(c_61_907), .sum(s_61_907), .in3(P_16[29]), .in2(P_15[31]), .in1(P_14[33]) );
  Fadder_ A_61_908( .carry(c_61_908), .sum(s_61_908), .in3(P_13[35]), .in2(P_12[37]), .in1(P_11[39]) );
  Fadder_ A_61_909( .carry(c_61_909), .sum(s_61_909), .in3(P_10[41]), .in2(P_9[43]), .in1(P_8[45]) );
  Fadder_ A_61_910( .carry(c_61_910), .sum(s_61_910), .in3(P_7[47]), .in2(P_6[49]), .in1(P_5[51]) );
  Fadder_ A_61_911( .carry(c_61_911), .sum(s_61_911), .in3(P_4[53]), .in2(P_3[55]), .in1(P_2[57]) );
  Fadder_ A_61_912( .carry(c_61_912), .sum(s_61_912), .in3(P_1[59]), .in2(P_0[61]), .in1(c_60_872) );
  Fadder_ A_61_913( .carry(c_61_913), .sum(s_61_913), .in3(c_60_882), .in2(c_60_881), .in1(c_60_880) );
  Fadder_ A_61_914( .carry(c_61_914), .sum(s_61_914), .in3(c_60_879), .in2(c_60_878), .in1(c_60_877) );
  Fadder_ A_61_915( .carry(c_61_915), .sum(s_61_915), .in3(c_60_876), .in2(c_60_875), .in1(c_60_874) );
  Fadder_ A_61_916( .carry(c_61_916), .sum(s_61_916), .in3(c_60_873), .in2(s_61_911), .in1(s_61_910) );
  Fadder_ A_61_917( .carry(c_61_917), .sum(s_61_917), .in3(s_61_909), .in2(s_61_908), .in1(s_61_907) );
  Fadder_ A_61_918( .carry(c_61_918), .sum(s_61_918), .in3(s_61_906), .in2(s_61_905), .in1(s_61_904) );
  Fadder_ A_61_919( .carry(c_61_919), .sum(s_61_919), .in3(s_61_903), .in2(s_61_902), .in1(s_61_912) );
  Fadder_ A_61_920( .carry(c_61_920), .sum(s_61_920), .in3(c_60_885), .in2(c_60_884), .in1(c_60_883) );
  Fadder_ A_61_921( .carry(c_61_921), .sum(s_61_921), .in3(c_60_886), .in2(s_61_915), .in1(s_61_914) );
  Fadder_ A_61_922( .carry(c_61_922), .sum(s_61_922), .in3(s_61_913), .in2(c_60_889), .in1(c_60_888) );
  Fadder_ A_61_923( .carry(c_61_923), .sum(s_61_923), .in3(c_60_887), .in2(s_61_916), .in1(s_61_918) );
  Fadder_ A_61_924( .carry(c_61_924), .sum(s_61_924), .in3(s_61_917), .in2(s_61_919), .in1(c_60_890) );
  Fadder_ A_61_925( .carry(c_61_925), .sum(s_61_925), .in3(s_61_920), .in2(c_60_892), .in1(c_60_891) );
  Fadder_ A_61_926( .carry(c_61_926), .sum(s_61_926), .in3(s_61_921), .in2(c_60_893), .in1(s_61_922) );
  Fadder_ A_61_927( .carry(c_61_927), .sum(s_61_927), .in3(s_61_923), .in2(c_60_894), .in1(s_61_924) );
  Fadder_ A_61_928( .carry(c_61_928), .sum(s_61_928), .in3(c_60_895), .in2(c_60_896), .in1(s_61_925) );
  Fadder_ A_61_929( .carry(c_61_929), .sum(s_61_929), .in3(s_61_926), .in2(c_60_897), .in1(s_61_927) );
  Fadder_ A_61_930( .carry(c_61_930), .sum(s_61_930), .in3(c_60_898), .in2(s_61_928), .in1(c_60_899) );
  Fadder_ A_61_931( .carry(c[61]), .sum(s[61]), .in3(s_61_929), .in2(c_60_900), .in1(s_61_930) );

  // ***** Bit 62 ***** //
  Hadder_ A_62_932( .carry(c_62_932), .sum(s_62_932), .in2(inc[62]), .in1(P_31[0]) );
  Fadder_ A_62_933( .carry(c_62_933), .sum(s_62_933), .in3(P_30[2]), .in2(P_29[4]), .in1(P_28[6]) );
  Fadder_ A_62_934( .carry(c_62_934), .sum(s_62_934), .in3(P_27[8]), .in2(P_26[10]), .in1(P_25[12]) );
  Fadder_ A_62_935( .carry(c_62_935), .sum(s_62_935), .in3(P_24[14]), .in2(P_23[16]), .in1(P_22[18]) );
  Fadder_ A_62_936( .carry(c_62_936), .sum(s_62_936), .in3(P_21[20]), .in2(P_20[22]), .in1(P_19[24]) );
  Fadder_ A_62_937( .carry(c_62_937), .sum(s_62_937), .in3(P_18[26]), .in2(P_17[28]), .in1(P_16[30]) );
  Fadder_ A_62_938( .carry(c_62_938), .sum(s_62_938), .in3(P_15[32]), .in2(P_14[34]), .in1(P_13[36]) );
  Fadder_ A_62_939( .carry(c_62_939), .sum(s_62_939), .in3(P_12[38]), .in2(P_11[40]), .in1(P_10[42]) );
  Fadder_ A_62_940( .carry(c_62_940), .sum(s_62_940), .in3(P_9[44]), .in2(P_8[46]), .in1(P_7[48]) );
  Fadder_ A_62_941( .carry(c_62_941), .sum(s_62_941), .in3(P_6[50]), .in2(P_5[52]), .in1(P_4[54]) );
  Fadder_ A_62_942( .carry(c_62_942), .sum(s_62_942), .in3(P_3[56]), .in2(P_2[58]), .in1(P_1[60]) );
  Fadder_ A_62_943( .carry(c_62_943), .sum(s_62_943), .in3(P_0[62]), .in2(c_61_911), .in1(c_61_910) );
  Fadder_ A_62_944( .carry(c_62_944), .sum(s_62_944), .in3(c_61_909), .in2(c_61_908), .in1(c_61_907) );
  Fadder_ A_62_945( .carry(c_62_945), .sum(s_62_945), .in3(c_61_906), .in2(c_61_905), .in1(c_61_904) );
  Fadder_ A_62_946( .carry(c_62_946), .sum(s_62_946), .in3(c_61_903), .in2(c_61_902), .in1(s_62_932) );
  Fadder_ A_62_947( .carry(c_62_947), .sum(s_62_947), .in3(s_62_942), .in2(s_62_941), .in1(s_62_940) );
  Fadder_ A_62_948( .carry(c_62_948), .sum(s_62_948), .in3(s_62_939), .in2(s_62_938), .in1(s_62_937) );
  Fadder_ A_62_949( .carry(c_62_949), .sum(s_62_949), .in3(s_62_936), .in2(s_62_935), .in1(s_62_934) );
  Fadder_ A_62_950( .carry(c_62_950), .sum(s_62_950), .in3(s_62_933), .in2(c_61_912), .in1(c_61_915) );
  Fadder_ A_62_951( .carry(c_62_951), .sum(s_62_951), .in3(c_61_914), .in2(c_61_913), .in1(s_62_943) );
  Fadder_ A_62_952( .carry(c_62_952), .sum(s_62_952), .in3(s_62_945), .in2(s_62_944), .in1(c_61_918) );
  Fadder_ A_62_953( .carry(c_62_953), .sum(s_62_953), .in3(c_61_917), .in2(c_61_916), .in1(s_62_946) );
  Fadder_ A_62_954( .carry(c_62_954), .sum(s_62_954), .in3(s_62_949), .in2(s_62_948), .in1(s_62_947) );
  Fadder_ A_62_955( .carry(c_62_955), .sum(s_62_955), .in3(c_61_919), .in2(c_61_920), .in1(s_62_950) );
  Fadder_ A_62_956( .carry(c_62_956), .sum(s_62_956), .in3(c_61_922), .in2(c_61_921), .in1(s_62_951) );
  Fadder_ A_62_957( .carry(c_62_957), .sum(s_62_957), .in3(c_61_923), .in2(s_62_952), .in1(s_62_953) );
  Fadder_ A_62_958( .carry(c_62_958), .sum(s_62_958), .in3(s_62_954), .in2(c_61_924), .in1(c_61_925) );
  Fadder_ A_62_959( .carry(c_62_959), .sum(s_62_959), .in3(s_62_955), .in2(c_61_926), .in1(s_62_956) );
  Fadder_ A_62_960( .carry(c_62_960), .sum(s_62_960), .in3(s_62_957), .in2(c_61_927), .in1(s_62_958) );
  Fadder_ A_62_961( .carry(c_62_961), .sum(s_62_961), .in3(c_61_928), .in2(s_62_959), .in1(c_61_929) );
  Fadder_ A_62_962( .carry(c[62]), .sum(s[62]), .in3(s_62_960), .in2(c_61_930), .in1(s_62_961) );

  // ***** Bit 63 ***** //
  Fadder_ A_63_963( .carry(c_63_963), .sum(s_63_963), .in3(inc[63]), .in2(P_31[1]), .in1(P_30[3]) );
  Fadder_ A_63_964( .carry(c_63_964), .sum(s_63_964), .in3(P_29[5]), .in2(P_28[7]), .in1(P_27[9]) );
  Fadder_ A_63_965( .carry(c_63_965), .sum(s_63_965), .in3(P_26[11]), .in2(P_25[13]), .in1(P_24[15]) );
  Fadder_ A_63_966( .carry(c_63_966), .sum(s_63_966), .in3(P_23[17]), .in2(P_22[19]), .in1(P_21[21]) );
  Fadder_ A_63_967( .carry(c_63_967), .sum(s_63_967), .in3(P_20[23]), .in2(P_19[25]), .in1(P_18[27]) );
  Fadder_ A_63_968( .carry(c_63_968), .sum(s_63_968), .in3(P_17[29]), .in2(P_16[31]), .in1(P_15[33]) );
  Fadder_ A_63_969( .carry(c_63_969), .sum(s_63_969), .in3(P_14[35]), .in2(P_13[37]), .in1(P_12[39]) );
  Fadder_ A_63_970( .carry(c_63_970), .sum(s_63_970), .in3(P_11[41]), .in2(P_10[43]), .in1(P_9[45]) );
  Fadder_ A_63_971( .carry(c_63_971), .sum(s_63_971), .in3(P_8[47]), .in2(P_7[49]), .in1(P_6[51]) );
  Fadder_ A_63_972( .carry(c_63_972), .sum(s_63_972), .in3(P_5[53]), .in2(P_4[55]), .in1(P_3[57]) );
  Fadder_ A_63_973( .carry(c_63_973), .sum(s_63_973), .in3(P_2[59]), .in2(P_1[61]), .in1(P_0[63]) );
  Fadder_ A_63_974( .carry(c_63_974), .sum(s_63_974), .in3(c_62_932), .in2(c_62_942), .in1(c_62_941) );
  Fadder_ A_63_975( .carry(c_63_975), .sum(s_63_975), .in3(c_62_940), .in2(c_62_939), .in1(c_62_938) );
  Fadder_ A_63_976( .carry(c_63_976), .sum(s_63_976), .in3(c_62_937), .in2(c_62_936), .in1(c_62_935) );
  Fadder_ A_63_977( .carry(c_63_977), .sum(s_63_977), .in3(c_62_934), .in2(c_62_933), .in1(s_63_973) );
  Fadder_ A_63_978( .carry(c_63_978), .sum(s_63_978), .in3(s_63_972), .in2(s_63_971), .in1(s_63_970) );
  Fadder_ A_63_979( .carry(c_63_979), .sum(s_63_979), .in3(s_63_969), .in2(s_63_968), .in1(s_63_967) );
  Fadder_ A_63_980( .carry(c_63_980), .sum(s_63_980), .in3(s_63_966), .in2(s_63_965), .in1(s_63_964) );
  Fadder_ A_63_981( .carry(c_63_981), .sum(s_63_981), .in3(s_63_963), .in2(c_62_945), .in1(c_62_944) );
  Fadder_ A_63_982( .carry(c_63_982), .sum(s_63_982), .in3(c_62_943), .in2(c_62_946), .in1(s_63_974) );
  Fadder_ A_63_983( .carry(c_63_983), .sum(s_63_983), .in3(s_63_976), .in2(s_63_975), .in1(c_62_949) );
  Fadder_ A_63_984( .carry(c_63_984), .sum(s_63_984), .in3(c_62_948), .in2(c_62_947), .in1(s_63_977) );
  Fadder_ A_63_985( .carry(c_63_985), .sum(s_63_985), .in3(s_63_980), .in2(s_63_979), .in1(s_63_978) );
  Fadder_ A_63_986( .carry(c_63_986), .sum(s_63_986), .in3(c_62_950), .in2(c_62_951), .in1(s_63_981) );
  Fadder_ A_63_987( .carry(c_63_987), .sum(s_63_987), .in3(c_62_953), .in2(c_62_952), .in1(s_63_982) );
  Fadder_ A_63_988( .carry(c_63_988), .sum(s_63_988), .in3(s_63_983), .in2(c_62_954), .in1(s_63_984) );
  Fadder_ A_63_989( .carry(c_63_989), .sum(s_63_989), .in3(s_63_985), .in2(c_62_955), .in1(c_62_956) );
  Fadder_ A_63_990( .carry(c_63_990), .sum(s_63_990), .in3(s_63_986), .in2(c_62_957), .in1(s_63_987) );
  Fadder_ A_63_991( .carry(c_63_991), .sum(s_63_991), .in3(s_63_988), .in2(c_62_958), .in1(s_63_989) );
  Fadder_ A_63_992( .carry(c_63_992), .sum(s_63_992), .in3(c_62_959), .in2(s_63_990), .in1(c_62_960) );
  Fadder_ A_63_993( .carry(c[63]), .sum(s[63]), .in3(s_63_991), .in2(c_62_961), .in1(s_63_992) );

  // ***** Bit 64 ***** //
  Hadder_ A_64_994( .carry(c_64_994), .sum(s_64_994), .in2(P_31[2]), .in1(P_30[4]) );
  Fadder_ A_64_995( .carry(c_64_995), .sum(s_64_995), .in3(P_29[6]), .in2(P_28[8]), .in1(P_27[10]) );
  Fadder_ A_64_996( .carry(c_64_996), .sum(s_64_996), .in3(P_26[12]), .in2(P_25[14]), .in1(P_24[16]) );
  Fadder_ A_64_997( .carry(c_64_997), .sum(s_64_997), .in3(P_23[18]), .in2(P_22[20]), .in1(P_21[22]) );
  Fadder_ A_64_998( .carry(c_64_998), .sum(s_64_998), .in3(P_20[24]), .in2(P_19[26]), .in1(P_18[28]) );
  Fadder_ A_64_999( .carry(c_64_999), .sum(s_64_999), .in3(P_17[30]), .in2(P_16[32]), .in1(P_15[34]) );
  Fadder_ A_64_1000( .carry(c_64_1000), .sum(s_64_1000), .in3(P_14[36]), .in2(P_13[38]), .in1(P_12[40]) );
  Fadder_ A_64_1001( .carry(c_64_1001), .sum(s_64_1001), .in3(P_11[42]), .in2(P_10[44]), .in1(P_9[46]) );
  Fadder_ A_64_1002( .carry(c_64_1002), .sum(s_64_1002), .in3(P_8[48]), .in2(P_7[50]), .in1(P_6[52]) );
  Fadder_ A_64_1003( .carry(c_64_1003), .sum(s_64_1003), .in3(P_5[54]), .in2(P_4[56]), .in1(P_3[58]) );
  Fadder_ A_64_1004( .carry(c_64_1004), .sum(s_64_1004), .in3(P_2[60]), .in2(P_1[62]), .in1(P_0[64]) );
  Fadder_ A_64_1005( .carry(c_64_1005), .sum(s_64_1005), .in3(c_63_973), .in2(c_63_972), .in1(c_63_971) );
  Fadder_ A_64_1006( .carry(c_64_1006), .sum(s_64_1006), .in3(c_63_970), .in2(c_63_969), .in1(c_63_968) );
  Fadder_ A_64_1007( .carry(c_64_1007), .sum(s_64_1007), .in3(c_63_967), .in2(c_63_966), .in1(c_63_965) );
  Fadder_ A_64_1008( .carry(c_64_1008), .sum(s_64_1008), .in3(c_63_964), .in2(c_63_963), .in1(s_64_994) );
  Fadder_ A_64_1009( .carry(c_64_1009), .sum(s_64_1009), .in3(s_64_1004), .in2(s_64_1003), .in1(s_64_1002) );
  Fadder_ A_64_1010( .carry(c_64_1010), .sum(s_64_1010), .in3(s_64_1001), .in2(s_64_1000), .in1(s_64_999) );
  Fadder_ A_64_1011( .carry(c_64_1011), .sum(s_64_1011), .in3(s_64_998), .in2(s_64_997), .in1(s_64_996) );
  Fadder_ A_64_1012( .carry(c_64_1012), .sum(s_64_1012), .in3(s_64_995), .in2(c_63_976), .in1(c_63_975) );
  Fadder_ A_64_1013( .carry(c_64_1013), .sum(s_64_1013), .in3(c_63_974), .in2(c_63_977), .in1(s_64_1007) );
  Fadder_ A_64_1014( .carry(c_64_1014), .sum(s_64_1014), .in3(s_64_1006), .in2(s_64_1005), .in1(c_63_980) );
  Fadder_ A_64_1015( .carry(c_64_1015), .sum(s_64_1015), .in3(c_63_979), .in2(c_63_978), .in1(s_64_1008) );
  Fadder_ A_64_1016( .carry(c_64_1016), .sum(s_64_1016), .in3(s_64_1011), .in2(s_64_1010), .in1(s_64_1009) );
  Fadder_ A_64_1017( .carry(c_64_1017), .sum(s_64_1017), .in3(c_63_981), .in2(c_63_982), .in1(s_64_1012) );
  Fadder_ A_64_1018( .carry(c_64_1018), .sum(s_64_1018), .in3(c_63_983), .in2(c_63_984), .in1(s_64_1013) );
  Fadder_ A_64_1019( .carry(c_64_1019), .sum(s_64_1019), .in3(s_64_1014), .in2(c_63_985), .in1(s_64_1015) );
  Fadder_ A_64_1020( .carry(c_64_1020), .sum(s_64_1020), .in3(s_64_1016), .in2(c_63_986), .in1(c_63_987) );
  Fadder_ A_64_1021( .carry(c_64_1021), .sum(s_64_1021), .in3(s_64_1017), .in2(c_63_988), .in1(s_64_1018) );
  Fadder_ A_64_1022( .carry(c_64_1022), .sum(s_64_1022), .in3(s_64_1019), .in2(c_63_989), .in1(s_64_1020) );
  Fadder_ A_64_1023( .carry(c_64_1023), .sum(s_64_1023), .in3(c_63_990), .in2(s_64_1021), .in1(c_63_991) );
  Fadder_ A_64_1024( .carry(c[64]), .sum(s[64]), .in3(s_64_1022), .in2(c_63_992), .in1(s_64_1023) );

  // ***** Bit 65 ***** //
  Fadder_ A_65_1025( .carry(c_65_1025), .sum(s_65_1025), .in3(sign_), .in2(P_31[3]), .in1(P_30[5]) );
  Fadder_ A_65_1026( .carry(c_65_1026), .sum(s_65_1026), .in3(P_29[7]), .in2(P_28[9]), .in1(P_27[11]) );
  Fadder_ A_65_1027( .carry(c_65_1027), .sum(s_65_1027), .in3(P_26[13]), .in2(P_25[15]), .in1(P_24[17]) );
  Fadder_ A_65_1028( .carry(c_65_1028), .sum(s_65_1028), .in3(P_23[19]), .in2(P_22[21]), .in1(P_21[23]) );
  Fadder_ A_65_1029( .carry(c_65_1029), .sum(s_65_1029), .in3(P_20[25]), .in2(P_19[27]), .in1(P_18[29]) );
  Fadder_ A_65_1030( .carry(c_65_1030), .sum(s_65_1030), .in3(P_17[31]), .in2(P_16[33]), .in1(P_15[35]) );
  Fadder_ A_65_1031( .carry(c_65_1031), .sum(s_65_1031), .in3(P_14[37]), .in2(P_13[39]), .in1(P_12[41]) );
  Fadder_ A_65_1032( .carry(c_65_1032), .sum(s_65_1032), .in3(P_11[43]), .in2(P_10[45]), .in1(P_9[47]) );
  Fadder_ A_65_1033( .carry(c_65_1033), .sum(s_65_1033), .in3(P_8[49]), .in2(P_7[51]), .in1(P_6[53]) );
  Fadder_ A_65_1034( .carry(c_65_1034), .sum(s_65_1034), .in3(P_5[55]), .in2(P_4[57]), .in1(P_3[59]) );
  Fadder_ A_65_1035( .carry(c_65_1035), .sum(s_65_1035), .in3(P_2[61]), .in2(P_1[63]), .in1(P_0[65]) );
  Fadder_ A_65_1036( .carry(c_65_1036), .sum(s_65_1036), .in3(c_64_994), .in2(c_64_1004), .in1(c_64_1003) );
  Fadder_ A_65_1037( .carry(c_65_1037), .sum(s_65_1037), .in3(c_64_1002), .in2(c_64_1001), .in1(c_64_1000) );
  Fadder_ A_65_1038( .carry(c_65_1038), .sum(s_65_1038), .in3(c_64_999), .in2(c_64_998), .in1(c_64_997) );
  Fadder_ A_65_1039( .carry(c_65_1039), .sum(s_65_1039), .in3(c_64_996), .in2(c_64_995), .in1(s_65_1025) );
  Fadder_ A_65_1040( .carry(c_65_1040), .sum(s_65_1040), .in3(s_65_1035), .in2(s_65_1034), .in1(s_65_1033) );
  Fadder_ A_65_1041( .carry(c_65_1041), .sum(s_65_1041), .in3(s_65_1032), .in2(s_65_1031), .in1(s_65_1030) );
  Fadder_ A_65_1042( .carry(c_65_1042), .sum(s_65_1042), .in3(s_65_1029), .in2(s_65_1028), .in1(s_65_1027) );
  Fadder_ A_65_1043( .carry(c_65_1043), .sum(s_65_1043), .in3(s_65_1026), .in2(c_64_1007), .in1(c_64_1006) );
  Fadder_ A_65_1044( .carry(c_65_1044), .sum(s_65_1044), .in3(c_64_1005), .in2(c_64_1008), .in1(s_65_1036) );
  Fadder_ A_65_1045( .carry(c_65_1045), .sum(s_65_1045), .in3(s_65_1038), .in2(s_65_1037), .in1(c_64_1011) );
  Fadder_ A_65_1046( .carry(c_65_1046), .sum(s_65_1046), .in3(c_64_1010), .in2(c_64_1009), .in1(s_65_1039) );
  Fadder_ A_65_1047( .carry(c_65_1047), .sum(s_65_1047), .in3(s_65_1042), .in2(s_65_1041), .in1(s_65_1040) );
  Fadder_ A_65_1048( .carry(c_65_1048), .sum(s_65_1048), .in3(c_64_1012), .in2(c_64_1013), .in1(s_65_1043) );
  Fadder_ A_65_1049( .carry(c_65_1049), .sum(s_65_1049), .in3(c_64_1015), .in2(c_64_1014), .in1(s_65_1044) );
  Fadder_ A_65_1050( .carry(c_65_1050), .sum(s_65_1050), .in3(s_65_1045), .in2(c_64_1016), .in1(s_65_1046) );
  Fadder_ A_65_1051( .carry(c_65_1051), .sum(s_65_1051), .in3(s_65_1047), .in2(c_64_1017), .in1(c_64_1018) );
  Fadder_ A_65_1052( .carry(c_65_1052), .sum(s_65_1052), .in3(s_65_1048), .in2(c_64_1019), .in1(s_65_1049) );
  Fadder_ A_65_1053( .carry(c_65_1053), .sum(s_65_1053), .in3(s_65_1050), .in2(c_64_1020), .in1(s_65_1051) );
  Fadder_ A_65_1054( .carry(c_65_1054), .sum(s_65_1054), .in3(c_64_1021), .in2(s_65_1052), .in1(c_64_1022) );
  Fadder_ A_65_1055( .carry(c[65]), .sum(s[65]), .in3(s_65_1053), .in2(c_64_1023), .in1(s_65_1054) );

  // ***** Bit 66 ***** //
  Hadder_ A_66_1056( .carry(c_66_1056), .sum(s_66_1056), .in2(sign_), .in1(P_31[4]) );
  Fadder_ A_66_1057( .carry(c_66_1057), .sum(s_66_1057), .in3(P_30[6]), .in2(P_29[8]), .in1(P_28[10]) );
  Fadder_ A_66_1058( .carry(c_66_1058), .sum(s_66_1058), .in3(P_27[12]), .in2(P_26[14]), .in1(P_25[16]) );
  Fadder_ A_66_1059( .carry(c_66_1059), .sum(s_66_1059), .in3(P_24[18]), .in2(P_23[20]), .in1(P_22[22]) );
  Fadder_ A_66_1060( .carry(c_66_1060), .sum(s_66_1060), .in3(P_21[24]), .in2(P_20[26]), .in1(P_19[28]) );
  Fadder_ A_66_1061( .carry(c_66_1061), .sum(s_66_1061), .in3(P_18[30]), .in2(P_17[32]), .in1(P_16[34]) );
  Fadder_ A_66_1062( .carry(c_66_1062), .sum(s_66_1062), .in3(P_15[36]), .in2(P_14[38]), .in1(P_13[40]) );
  Fadder_ A_66_1063( .carry(c_66_1063), .sum(s_66_1063), .in3(P_12[42]), .in2(P_11[44]), .in1(P_10[46]) );
  Fadder_ A_66_1064( .carry(c_66_1064), .sum(s_66_1064), .in3(P_9[48]), .in2(P_8[50]), .in1(P_7[52]) );
  Fadder_ A_66_1065( .carry(c_66_1065), .sum(s_66_1065), .in3(P_6[54]), .in2(P_5[56]), .in1(P_4[58]) );
  Fadder_ A_66_1066( .carry(c_66_1066), .sum(s_66_1066), .in3(P_3[60]), .in2(P_2[62]), .in1(P_1[64]) );
  Fadder_ A_66_1067( .carry(c_66_1067), .sum(s_66_1067), .in3(c_65_1035), .in2(c_65_1034), .in1(c_65_1033) );
  Fadder_ A_66_1068( .carry(c_66_1068), .sum(s_66_1068), .in3(c_65_1032), .in2(c_65_1031), .in1(c_65_1030) );
  Fadder_ A_66_1069( .carry(c_66_1069), .sum(s_66_1069), .in3(c_65_1029), .in2(c_65_1028), .in1(c_65_1027) );
  Fadder_ A_66_1070( .carry(c_66_1070), .sum(s_66_1070), .in3(c_65_1026), .in2(c_65_1025), .in1(s_66_1056) );
  Fadder_ A_66_1071( .carry(c_66_1071), .sum(s_66_1071), .in3(s_66_1066), .in2(s_66_1065), .in1(s_66_1064) );
  Fadder_ A_66_1072( .carry(c_66_1072), .sum(s_66_1072), .in3(s_66_1063), .in2(s_66_1062), .in1(s_66_1061) );
  Fadder_ A_66_1073( .carry(c_66_1073), .sum(s_66_1073), .in3(s_66_1060), .in2(s_66_1059), .in1(s_66_1058) );
  Fadder_ A_66_1074( .carry(c_66_1074), .sum(s_66_1074), .in3(s_66_1057), .in2(c_65_1038), .in1(c_65_1037) );
  Fadder_ A_66_1075( .carry(c_66_1075), .sum(s_66_1075), .in3(c_65_1036), .in2(c_65_1039), .in1(s_66_1069) );
  Fadder_ A_66_1076( .carry(c_66_1076), .sum(s_66_1076), .in3(s_66_1068), .in2(s_66_1067), .in1(c_65_1042) );
  Fadder_ A_66_1077( .carry(c_66_1077), .sum(s_66_1077), .in3(c_65_1041), .in2(c_65_1040), .in1(s_66_1070) );
  Fadder_ A_66_1078( .carry(c_66_1078), .sum(s_66_1078), .in3(s_66_1073), .in2(s_66_1072), .in1(s_66_1071) );
  Fadder_ A_66_1079( .carry(c_66_1079), .sum(s_66_1079), .in3(c_65_1043), .in2(c_65_1044), .in1(s_66_1074) );
  Fadder_ A_66_1080( .carry(c_66_1080), .sum(s_66_1080), .in3(c_65_1046), .in2(c_65_1045), .in1(s_66_1075) );
  Fadder_ A_66_1081( .carry(c_66_1081), .sum(s_66_1081), .in3(s_66_1076), .in2(c_65_1047), .in1(s_66_1077) );
  Fadder_ A_66_1082( .carry(c_66_1082), .sum(s_66_1082), .in3(s_66_1078), .in2(c_65_1048), .in1(c_65_1049) );
  Fadder_ A_66_1083( .carry(c_66_1083), .sum(s_66_1083), .in3(s_66_1079), .in2(c_65_1050), .in1(s_66_1080) );
  Fadder_ A_66_1084( .carry(c_66_1084), .sum(s_66_1084), .in3(s_66_1081), .in2(c_65_1051), .in1(s_66_1082) );
  Fadder_ A_66_1085( .carry(c_66_1085), .sum(s_66_1085), .in3(c_65_1052), .in2(s_66_1083), .in1(c_65_1053) );
  Fadder_ A_66_1086( .carry(c[66]), .sum(s[66]), .in3(s_66_1084), .in2(c_65_1054), .in1(s_66_1085) );

  // ***** Bit 67 ***** //
  Fadder_ A_67_1087( .carry(c_67_1087), .sum(s_67_1087), .in3(P_31[5]), .in2(P_30[7]), .in1(P_29[9]) );
  Fadder_ A_67_1088( .carry(c_67_1088), .sum(s_67_1088), .in3(P_28[11]), .in2(P_27[13]), .in1(P_26[15]) );
  Fadder_ A_67_1089( .carry(c_67_1089), .sum(s_67_1089), .in3(P_25[17]), .in2(P_24[19]), .in1(P_23[21]) );
  Fadder_ A_67_1090( .carry(c_67_1090), .sum(s_67_1090), .in3(P_22[23]), .in2(P_21[25]), .in1(P_20[27]) );
  Fadder_ A_67_1091( .carry(c_67_1091), .sum(s_67_1091), .in3(P_19[29]), .in2(P_18[31]), .in1(P_17[33]) );
  Fadder_ A_67_1092( .carry(c_67_1092), .sum(s_67_1092), .in3(P_16[35]), .in2(P_15[37]), .in1(P_14[39]) );
  Fadder_ A_67_1093( .carry(c_67_1093), .sum(s_67_1093), .in3(P_13[41]), .in2(P_12[43]), .in1(P_11[45]) );
  Fadder_ A_67_1094( .carry(c_67_1094), .sum(s_67_1094), .in3(P_10[47]), .in2(P_9[49]), .in1(P_8[51]) );
  Fadder_ A_67_1095( .carry(c_67_1095), .sum(s_67_1095), .in3(P_7[53]), .in2(P_6[55]), .in1(P_5[57]) );
  Fadder_ A_67_1096( .carry(c_67_1096), .sum(s_67_1096), .in3(P_4[59]), .in2(P_3[61]), .in1(P_2[63]) );
  Fadder_ A_67_1097( .carry(c_67_1097), .sum(s_67_1097), .in3(P_1[65]), .in2(c_66_1056), .in1(c_66_1066) );
  Fadder_ A_67_1098( .carry(c_67_1098), .sum(s_67_1098), .in3(c_66_1065), .in2(c_66_1064), .in1(c_66_1063) );
  Fadder_ A_67_1099( .carry(c_67_1099), .sum(s_67_1099), .in3(c_66_1062), .in2(c_66_1061), .in1(c_66_1060) );
  Fadder_ A_67_1100( .carry(c_67_1100), .sum(s_67_1100), .in3(c_66_1059), .in2(c_66_1058), .in1(c_66_1057) );
  Fadder_ A_67_1101( .carry(c_67_1101), .sum(s_67_1101), .in3(s_67_1096), .in2(s_67_1095), .in1(s_67_1094) );
  Fadder_ A_67_1102( .carry(c_67_1102), .sum(s_67_1102), .in3(s_67_1093), .in2(s_67_1092), .in1(s_67_1091) );
  Fadder_ A_67_1103( .carry(c_67_1103), .sum(s_67_1103), .in3(s_67_1090), .in2(s_67_1089), .in1(s_67_1088) );
  Fadder_ A_67_1104( .carry(c_67_1104), .sum(s_67_1104), .in3(s_67_1087), .in2(c_66_1070), .in1(c_66_1069) );
  Fadder_ A_67_1105( .carry(c_67_1105), .sum(s_67_1105), .in3(c_66_1068), .in2(c_66_1067), .in1(s_67_1097) );
  Fadder_ A_67_1106( .carry(c_67_1106), .sum(s_67_1106), .in3(s_67_1100), .in2(s_67_1099), .in1(s_67_1098) );
  Fadder_ A_67_1107( .carry(c_67_1107), .sum(s_67_1107), .in3(c_66_1073), .in2(c_66_1072), .in1(c_66_1071) );
  Fadder_ A_67_1108( .carry(c_67_1108), .sum(s_67_1108), .in3(s_67_1103), .in2(s_67_1102), .in1(s_67_1101) );
  Fadder_ A_67_1109( .carry(c_67_1109), .sum(s_67_1109), .in3(c_66_1074), .in2(c_66_1075), .in1(s_67_1104) );
  Fadder_ A_67_1110( .carry(c_67_1110), .sum(s_67_1110), .in3(c_66_1077), .in2(c_66_1076), .in1(s_67_1105) );
  Fadder_ A_67_1111( .carry(c_67_1111), .sum(s_67_1111), .in3(s_67_1107), .in2(s_67_1106), .in1(c_66_1078) );
  Fadder_ A_67_1112( .carry(c_67_1112), .sum(s_67_1112), .in3(s_67_1108), .in2(c_66_1079), .in1(c_66_1080) );
  Fadder_ A_67_1113( .carry(c_67_1113), .sum(s_67_1113), .in3(s_67_1109), .in2(c_66_1081), .in1(s_67_1110) );
  Fadder_ A_67_1114( .carry(c_67_1114), .sum(s_67_1114), .in3(s_67_1111), .in2(c_66_1082), .in1(s_67_1112) );
  Fadder_ A_67_1115( .carry(c_67_1115), .sum(s_67_1115), .in3(c_66_1083), .in2(s_67_1113), .in1(c_66_1084) );
  Fadder_ A_67_1116( .carry(c[67]), .sum(s[67]), .in3(s_67_1114), .in2(c_66_1085), .in1(s_67_1115) );

  // ***** Bit 68 ***** //
  Hadder_ A_68_1117( .carry(c_68_1117), .sum(s_68_1117), .in2(sign_), .in1(P_31[6]) );
  Fadder_ A_68_1118( .carry(c_68_1118), .sum(s_68_1118), .in3(P_30[8]), .in2(P_29[10]), .in1(P_28[12]) );
  Fadder_ A_68_1119( .carry(c_68_1119), .sum(s_68_1119), .in3(P_27[14]), .in2(P_26[16]), .in1(P_25[18]) );
  Fadder_ A_68_1120( .carry(c_68_1120), .sum(s_68_1120), .in3(P_24[20]), .in2(P_23[22]), .in1(P_22[24]) );
  Fadder_ A_68_1121( .carry(c_68_1121), .sum(s_68_1121), .in3(P_21[26]), .in2(P_20[28]), .in1(P_19[30]) );
  Fadder_ A_68_1122( .carry(c_68_1122), .sum(s_68_1122), .in3(P_18[32]), .in2(P_17[34]), .in1(P_16[36]) );
  Fadder_ A_68_1123( .carry(c_68_1123), .sum(s_68_1123), .in3(P_15[38]), .in2(P_14[40]), .in1(P_13[42]) );
  Fadder_ A_68_1124( .carry(c_68_1124), .sum(s_68_1124), .in3(P_12[44]), .in2(P_11[46]), .in1(P_10[48]) );
  Fadder_ A_68_1125( .carry(c_68_1125), .sum(s_68_1125), .in3(P_9[50]), .in2(P_8[52]), .in1(P_7[54]) );
  Fadder_ A_68_1126( .carry(c_68_1126), .sum(s_68_1126), .in3(P_6[56]), .in2(P_5[58]), .in1(P_4[60]) );
  Fadder_ A_68_1127( .carry(c_68_1127), .sum(s_68_1127), .in3(P_3[62]), .in2(P_2[64]), .in1(c_67_1096) );
  Fadder_ A_68_1128( .carry(c_68_1128), .sum(s_68_1128), .in3(c_67_1095), .in2(c_67_1094), .in1(c_67_1093) );
  Fadder_ A_68_1129( .carry(c_68_1129), .sum(s_68_1129), .in3(c_67_1092), .in2(c_67_1091), .in1(c_67_1090) );
  Fadder_ A_68_1130( .carry(c_68_1130), .sum(s_68_1130), .in3(c_67_1089), .in2(c_67_1088), .in1(c_67_1087) );
  Fadder_ A_68_1131( .carry(c_68_1131), .sum(s_68_1131), .in3(s_68_1117), .in2(s_68_1126), .in1(s_68_1125) );
  Fadder_ A_68_1132( .carry(c_68_1132), .sum(s_68_1132), .in3(s_68_1124), .in2(s_68_1123), .in1(s_68_1122) );
  Fadder_ A_68_1133( .carry(c_68_1133), .sum(s_68_1133), .in3(s_68_1121), .in2(s_68_1120), .in1(s_68_1119) );
  Fadder_ A_68_1134( .carry(c_68_1134), .sum(s_68_1134), .in3(s_68_1118), .in2(c_67_1097), .in1(c_67_1100) );
  Fadder_ A_68_1135( .carry(c_68_1135), .sum(s_68_1135), .in3(c_67_1099), .in2(c_67_1098), .in1(s_68_1127) );
  Fadder_ A_68_1136( .carry(c_68_1136), .sum(s_68_1136), .in3(s_68_1130), .in2(s_68_1129), .in1(s_68_1128) );
  Fadder_ A_68_1137( .carry(c_68_1137), .sum(s_68_1137), .in3(c_67_1103), .in2(c_67_1102), .in1(c_67_1101) );
  Fadder_ A_68_1138( .carry(c_68_1138), .sum(s_68_1138), .in3(s_68_1131), .in2(s_68_1133), .in1(s_68_1132) );
  Fadder_ A_68_1139( .carry(c_68_1139), .sum(s_68_1139), .in3(c_67_1104), .in2(c_67_1105), .in1(s_68_1134) );
  Fadder_ A_68_1140( .carry(c_68_1140), .sum(s_68_1140), .in3(c_67_1107), .in2(c_67_1106), .in1(s_68_1135) );
  Fadder_ A_68_1141( .carry(c_68_1141), .sum(s_68_1141), .in3(s_68_1137), .in2(s_68_1136), .in1(c_67_1108) );
  Fadder_ A_68_1142( .carry(c_68_1142), .sum(s_68_1142), .in3(s_68_1138), .in2(c_67_1109), .in1(c_67_1110) );
  Fadder_ A_68_1143( .carry(c_68_1143), .sum(s_68_1143), .in3(s_68_1139), .in2(c_67_1111), .in1(s_68_1140) );
  Fadder_ A_68_1144( .carry(c_68_1144), .sum(s_68_1144), .in3(s_68_1141), .in2(c_67_1112), .in1(s_68_1142) );
  Fadder_ A_68_1145( .carry(c_68_1145), .sum(s_68_1145), .in3(c_67_1113), .in2(s_68_1143), .in1(c_67_1114) );
  Fadder_ A_68_1146( .carry(c[68]), .sum(s[68]), .in3(s_68_1144), .in2(c_67_1115), .in1(s_68_1145) );

  // ***** Bit 69 ***** //
  Fadder_ A_69_1147( .carry(c_69_1147), .sum(s_69_1147), .in3(P_31[7]), .in2(P_30[9]), .in1(P_29[11]) );
  Fadder_ A_69_1148( .carry(c_69_1148), .sum(s_69_1148), .in3(P_28[13]), .in2(P_27[15]), .in1(P_26[17]) );
  Fadder_ A_69_1149( .carry(c_69_1149), .sum(s_69_1149), .in3(P_25[19]), .in2(P_24[21]), .in1(P_23[23]) );
  Fadder_ A_69_1150( .carry(c_69_1150), .sum(s_69_1150), .in3(P_22[25]), .in2(P_21[27]), .in1(P_20[29]) );
  Fadder_ A_69_1151( .carry(c_69_1151), .sum(s_69_1151), .in3(P_19[31]), .in2(P_18[33]), .in1(P_17[35]) );
  Fadder_ A_69_1152( .carry(c_69_1152), .sum(s_69_1152), .in3(P_16[37]), .in2(P_15[39]), .in1(P_14[41]) );
  Fadder_ A_69_1153( .carry(c_69_1153), .sum(s_69_1153), .in3(P_13[43]), .in2(P_12[45]), .in1(P_11[47]) );
  Fadder_ A_69_1154( .carry(c_69_1154), .sum(s_69_1154), .in3(P_10[49]), .in2(P_9[51]), .in1(P_8[53]) );
  Fadder_ A_69_1155( .carry(c_69_1155), .sum(s_69_1155), .in3(P_7[55]), .in2(P_6[57]), .in1(P_5[59]) );
  Fadder_ A_69_1156( .carry(c_69_1156), .sum(s_69_1156), .in3(P_4[61]), .in2(P_3[63]), .in1(P_2[65]) );
  Fadder_ A_69_1157( .carry(c_69_1157), .sum(s_69_1157), .in3(c_68_1117), .in2(c_68_1126), .in1(c_68_1125) );
  Fadder_ A_69_1158( .carry(c_69_1158), .sum(s_69_1158), .in3(c_68_1124), .in2(c_68_1123), .in1(c_68_1122) );
  Fadder_ A_69_1159( .carry(c_69_1159), .sum(s_69_1159), .in3(c_68_1121), .in2(c_68_1120), .in1(c_68_1119) );
  Fadder_ A_69_1160( .carry(c_69_1160), .sum(s_69_1160), .in3(c_68_1118), .in2(s_69_1156), .in1(s_69_1155) );
  Fadder_ A_69_1161( .carry(c_69_1161), .sum(s_69_1161), .in3(s_69_1154), .in2(s_69_1153), .in1(s_69_1152) );
  Fadder_ A_69_1162( .carry(c_69_1162), .sum(s_69_1162), .in3(s_69_1151), .in2(s_69_1150), .in1(s_69_1149) );
  Fadder_ A_69_1163( .carry(c_69_1163), .sum(s_69_1163), .in3(s_69_1148), .in2(s_69_1147), .in1(c_68_1127) );
  Fadder_ A_69_1164( .carry(c_69_1164), .sum(s_69_1164), .in3(c_68_1130), .in2(c_68_1129), .in1(c_68_1128) );
  Fadder_ A_69_1165( .carry(c_69_1165), .sum(s_69_1165), .in3(s_69_1157), .in2(s_69_1159), .in1(s_69_1158) );
  Fadder_ A_69_1166( .carry(c_69_1166), .sum(s_69_1166), .in3(c_68_1133), .in2(c_68_1132), .in1(c_68_1131) );
  Fadder_ A_69_1167( .carry(c_69_1167), .sum(s_69_1167), .in3(s_69_1160), .in2(s_69_1162), .in1(s_69_1161) );
  Fadder_ A_69_1168( .carry(c_69_1168), .sum(s_69_1168), .in3(c_68_1134), .in2(s_69_1163), .in1(c_68_1135) );
  Fadder_ A_69_1169( .carry(c_69_1169), .sum(s_69_1169), .in3(s_69_1164), .in2(c_68_1137), .in1(c_68_1136) );
  Fadder_ A_69_1170( .carry(c_69_1170), .sum(s_69_1170), .in3(s_69_1165), .in2(s_69_1166), .in1(c_68_1138) );
  Fadder_ A_69_1171( .carry(c_69_1171), .sum(s_69_1171), .in3(s_69_1167), .in2(c_68_1139), .in1(s_69_1168) );
  Fadder_ A_69_1172( .carry(c_69_1172), .sum(s_69_1172), .in3(c_68_1140), .in2(s_69_1169), .in1(c_68_1141) );
  Fadder_ A_69_1173( .carry(c_69_1173), .sum(s_69_1173), .in3(s_69_1170), .in2(c_68_1142), .in1(s_69_1171) );
  Fadder_ A_69_1174( .carry(c_69_1174), .sum(s_69_1174), .in3(c_68_1143), .in2(s_69_1172), .in1(c_68_1144) );
  Fadder_ A_69_1175( .carry(c[69]), .sum(s[69]), .in3(s_69_1173), .in2(c_68_1145), .in1(s_69_1174) );

  // ***** Bit 70 ***** //
  Hadder_ A_70_1176( .carry(c_70_1176), .sum(s_70_1176), .in2(sign_), .in1(P_31[8]) );
  Fadder_ A_70_1177( .carry(c_70_1177), .sum(s_70_1177), .in3(P_30[10]), .in2(P_29[12]), .in1(P_28[14]) );
  Fadder_ A_70_1178( .carry(c_70_1178), .sum(s_70_1178), .in3(P_27[16]), .in2(P_26[18]), .in1(P_25[20]) );
  Fadder_ A_70_1179( .carry(c_70_1179), .sum(s_70_1179), .in3(P_24[22]), .in2(P_23[24]), .in1(P_22[26]) );
  Fadder_ A_70_1180( .carry(c_70_1180), .sum(s_70_1180), .in3(P_21[28]), .in2(P_20[30]), .in1(P_19[32]) );
  Fadder_ A_70_1181( .carry(c_70_1181), .sum(s_70_1181), .in3(P_18[34]), .in2(P_17[36]), .in1(P_16[38]) );
  Fadder_ A_70_1182( .carry(c_70_1182), .sum(s_70_1182), .in3(P_15[40]), .in2(P_14[42]), .in1(P_13[44]) );
  Fadder_ A_70_1183( .carry(c_70_1183), .sum(s_70_1183), .in3(P_12[46]), .in2(P_11[48]), .in1(P_10[50]) );
  Fadder_ A_70_1184( .carry(c_70_1184), .sum(s_70_1184), .in3(P_9[52]), .in2(P_8[54]), .in1(P_7[56]) );
  Fadder_ A_70_1185( .carry(c_70_1185), .sum(s_70_1185), .in3(P_6[58]), .in2(P_5[60]), .in1(P_4[62]) );
  Fadder_ A_70_1186( .carry(c_70_1186), .sum(s_70_1186), .in3(P_3[64]), .in2(c_69_1156), .in1(c_69_1155) );
  Fadder_ A_70_1187( .carry(c_70_1187), .sum(s_70_1187), .in3(c_69_1154), .in2(c_69_1153), .in1(c_69_1152) );
  Fadder_ A_70_1188( .carry(c_70_1188), .sum(s_70_1188), .in3(c_69_1151), .in2(c_69_1150), .in1(c_69_1149) );
  Fadder_ A_70_1189( .carry(c_70_1189), .sum(s_70_1189), .in3(c_69_1148), .in2(c_69_1147), .in1(s_70_1176) );
  Fadder_ A_70_1190( .carry(c_70_1190), .sum(s_70_1190), .in3(s_70_1185), .in2(s_70_1184), .in1(s_70_1183) );
  Fadder_ A_70_1191( .carry(c_70_1191), .sum(s_70_1191), .in3(s_70_1182), .in2(s_70_1181), .in1(s_70_1180) );
  Fadder_ A_70_1192( .carry(c_70_1192), .sum(s_70_1192), .in3(s_70_1179), .in2(s_70_1178), .in1(s_70_1177) );
  Fadder_ A_70_1193( .carry(c_70_1193), .sum(s_70_1193), .in3(c_69_1159), .in2(c_69_1158), .in1(c_69_1157) );
  Fadder_ A_70_1194( .carry(c_70_1194), .sum(s_70_1194), .in3(s_70_1186), .in2(s_70_1188), .in1(s_70_1187) );
  Fadder_ A_70_1195( .carry(c_70_1195), .sum(s_70_1195), .in3(c_69_1162), .in2(c_69_1161), .in1(c_69_1160) );
  Fadder_ A_70_1196( .carry(c_70_1196), .sum(s_70_1196), .in3(s_70_1189), .in2(s_70_1192), .in1(s_70_1191) );
  Fadder_ A_70_1197( .carry(c_70_1197), .sum(s_70_1197), .in3(s_70_1190), .in2(c_69_1163), .in1(c_69_1164) );
  Fadder_ A_70_1198( .carry(c_70_1198), .sum(s_70_1198), .in3(s_70_1193), .in2(c_69_1166), .in1(c_69_1165) );
  Fadder_ A_70_1199( .carry(c_70_1199), .sum(s_70_1199), .in3(s_70_1194), .in2(s_70_1195), .in1(c_69_1167) );
  Fadder_ A_70_1200( .carry(c_70_1200), .sum(s_70_1200), .in3(s_70_1196), .in2(c_69_1168), .in1(s_70_1197) );
  Fadder_ A_70_1201( .carry(c_70_1201), .sum(s_70_1201), .in3(c_69_1169), .in2(s_70_1198), .in1(c_69_1170) );
  Fadder_ A_70_1202( .carry(c_70_1202), .sum(s_70_1202), .in3(s_70_1199), .in2(c_69_1171), .in1(s_70_1200) );
  Fadder_ A_70_1203( .carry(c_70_1203), .sum(s_70_1203), .in3(c_69_1172), .in2(s_70_1201), .in1(c_69_1173) );
  Fadder_ A_70_1204( .carry(c[70]), .sum(s[70]), .in3(s_70_1202), .in2(c_69_1174), .in1(s_70_1203) );

  // ***** Bit 71 ***** //
  Fadder_ A_71_1205( .carry(c_71_1205), .sum(s_71_1205), .in3(P_31[9]), .in2(P_30[11]), .in1(P_29[13]) );
  Fadder_ A_71_1206( .carry(c_71_1206), .sum(s_71_1206), .in3(P_28[15]), .in2(P_27[17]), .in1(P_26[19]) );
  Fadder_ A_71_1207( .carry(c_71_1207), .sum(s_71_1207), .in3(P_25[21]), .in2(P_24[23]), .in1(P_23[25]) );
  Fadder_ A_71_1208( .carry(c_71_1208), .sum(s_71_1208), .in3(P_22[27]), .in2(P_21[29]), .in1(P_20[31]) );
  Fadder_ A_71_1209( .carry(c_71_1209), .sum(s_71_1209), .in3(P_19[33]), .in2(P_18[35]), .in1(P_17[37]) );
  Fadder_ A_71_1210( .carry(c_71_1210), .sum(s_71_1210), .in3(P_16[39]), .in2(P_15[41]), .in1(P_14[43]) );
  Fadder_ A_71_1211( .carry(c_71_1211), .sum(s_71_1211), .in3(P_13[45]), .in2(P_12[47]), .in1(P_11[49]) );
  Fadder_ A_71_1212( .carry(c_71_1212), .sum(s_71_1212), .in3(P_10[51]), .in2(P_9[53]), .in1(P_8[55]) );
  Fadder_ A_71_1213( .carry(c_71_1213), .sum(s_71_1213), .in3(P_7[57]), .in2(P_6[59]), .in1(P_5[61]) );
  Fadder_ A_71_1214( .carry(c_71_1214), .sum(s_71_1214), .in3(P_4[63]), .in2(P_3[65]), .in1(c_70_1176) );
  Fadder_ A_71_1215( .carry(c_71_1215), .sum(s_71_1215), .in3(c_70_1185), .in2(c_70_1184), .in1(c_70_1183) );
  Fadder_ A_71_1216( .carry(c_71_1216), .sum(s_71_1216), .in3(c_70_1182), .in2(c_70_1181), .in1(c_70_1180) );
  Fadder_ A_71_1217( .carry(c_71_1217), .sum(s_71_1217), .in3(c_70_1179), .in2(c_70_1178), .in1(c_70_1177) );
  Fadder_ A_71_1218( .carry(c_71_1218), .sum(s_71_1218), .in3(s_71_1213), .in2(s_71_1212), .in1(s_71_1211) );
  Fadder_ A_71_1219( .carry(c_71_1219), .sum(s_71_1219), .in3(s_71_1210), .in2(s_71_1209), .in1(s_71_1208) );
  Fadder_ A_71_1220( .carry(c_71_1220), .sum(s_71_1220), .in3(s_71_1207), .in2(s_71_1206), .in1(s_71_1205) );
  Fadder_ A_71_1221( .carry(c_71_1221), .sum(s_71_1221), .in3(s_71_1214), .in2(c_70_1189), .in1(c_70_1188) );
  Fadder_ A_71_1222( .carry(c_71_1222), .sum(s_71_1222), .in3(c_70_1187), .in2(c_70_1186), .in1(s_71_1217) );
  Fadder_ A_71_1223( .carry(c_71_1223), .sum(s_71_1223), .in3(s_71_1216), .in2(s_71_1215), .in1(c_70_1192) );
  Fadder_ A_71_1224( .carry(c_71_1224), .sum(s_71_1224), .in3(c_70_1191), .in2(c_70_1190), .in1(s_71_1220) );
  Fadder_ A_71_1225( .carry(c_71_1225), .sum(s_71_1225), .in3(s_71_1219), .in2(s_71_1218), .in1(c_70_1193) );
  Fadder_ A_71_1226( .carry(c_71_1226), .sum(s_71_1226), .in3(s_71_1221), .in2(c_70_1195), .in1(c_70_1194) );
  Fadder_ A_71_1227( .carry(c_71_1227), .sum(s_71_1227), .in3(s_71_1222), .in2(s_71_1223), .in1(c_70_1196) );
  Fadder_ A_71_1228( .carry(c_71_1228), .sum(s_71_1228), .in3(s_71_1224), .in2(c_70_1197), .in1(s_71_1225) );
  Fadder_ A_71_1229( .carry(c_71_1229), .sum(s_71_1229), .in3(c_70_1198), .in2(s_71_1226), .in1(c_70_1199) );
  Fadder_ A_71_1230( .carry(c_71_1230), .sum(s_71_1230), .in3(s_71_1227), .in2(c_70_1200), .in1(s_71_1228) );
  Fadder_ A_71_1231( .carry(c_71_1231), .sum(s_71_1231), .in3(c_70_1201), .in2(s_71_1229), .in1(c_70_1202) );
  Fadder_ A_71_1232( .carry(c[71]), .sum(s[71]), .in3(s_71_1230), .in2(c_70_1203), .in1(s_71_1231) );

  // ***** Bit 72 ***** //
  Hadder_ A_72_1233( .carry(c_72_1233), .sum(s_72_1233), .in2(sign_), .in1(P_31[10]) );
  Fadder_ A_72_1234( .carry(c_72_1234), .sum(s_72_1234), .in3(P_30[12]), .in2(P_29[14]), .in1(P_28[16]) );
  Fadder_ A_72_1235( .carry(c_72_1235), .sum(s_72_1235), .in3(P_27[18]), .in2(P_26[20]), .in1(P_25[22]) );
  Fadder_ A_72_1236( .carry(c_72_1236), .sum(s_72_1236), .in3(P_24[24]), .in2(P_23[26]), .in1(P_22[28]) );
  Fadder_ A_72_1237( .carry(c_72_1237), .sum(s_72_1237), .in3(P_21[30]), .in2(P_20[32]), .in1(P_19[34]) );
  Fadder_ A_72_1238( .carry(c_72_1238), .sum(s_72_1238), .in3(P_18[36]), .in2(P_17[38]), .in1(P_16[40]) );
  Fadder_ A_72_1239( .carry(c_72_1239), .sum(s_72_1239), .in3(P_15[42]), .in2(P_14[44]), .in1(P_13[46]) );
  Fadder_ A_72_1240( .carry(c_72_1240), .sum(s_72_1240), .in3(P_12[48]), .in2(P_11[50]), .in1(P_10[52]) );
  Fadder_ A_72_1241( .carry(c_72_1241), .sum(s_72_1241), .in3(P_9[54]), .in2(P_8[56]), .in1(P_7[58]) );
  Fadder_ A_72_1242( .carry(c_72_1242), .sum(s_72_1242), .in3(P_6[60]), .in2(P_5[62]), .in1(P_4[64]) );
  Fadder_ A_72_1243( .carry(c_72_1243), .sum(s_72_1243), .in3(c_71_1213), .in2(c_71_1212), .in1(c_71_1211) );
  Fadder_ A_72_1244( .carry(c_72_1244), .sum(s_72_1244), .in3(c_71_1210), .in2(c_71_1209), .in1(c_71_1208) );
  Fadder_ A_72_1245( .carry(c_72_1245), .sum(s_72_1245), .in3(c_71_1207), .in2(c_71_1206), .in1(c_71_1205) );
  Fadder_ A_72_1246( .carry(c_72_1246), .sum(s_72_1246), .in3(s_72_1233), .in2(s_72_1242), .in1(s_72_1241) );
  Fadder_ A_72_1247( .carry(c_72_1247), .sum(s_72_1247), .in3(s_72_1240), .in2(s_72_1239), .in1(s_72_1238) );
  Fadder_ A_72_1248( .carry(c_72_1248), .sum(s_72_1248), .in3(s_72_1237), .in2(s_72_1236), .in1(s_72_1235) );
  Fadder_ A_72_1249( .carry(c_72_1249), .sum(s_72_1249), .in3(s_72_1234), .in2(c_71_1214), .in1(c_71_1217) );
  Fadder_ A_72_1250( .carry(c_72_1250), .sum(s_72_1250), .in3(c_71_1216), .in2(c_71_1215), .in1(s_72_1245) );
  Fadder_ A_72_1251( .carry(c_72_1251), .sum(s_72_1251), .in3(s_72_1244), .in2(s_72_1243), .in1(c_71_1220) );
  Fadder_ A_72_1252( .carry(c_72_1252), .sum(s_72_1252), .in3(c_71_1219), .in2(c_71_1218), .in1(s_72_1246) );
  Fadder_ A_72_1253( .carry(c_72_1253), .sum(s_72_1253), .in3(s_72_1248), .in2(s_72_1247), .in1(c_71_1221) );
  Fadder_ A_72_1254( .carry(c_72_1254), .sum(s_72_1254), .in3(c_71_1222), .in2(s_72_1249), .in1(c_71_1223) );
  Fadder_ A_72_1255( .carry(c_72_1255), .sum(s_72_1255), .in3(c_71_1224), .in2(s_72_1250), .in1(s_72_1251) );
  Fadder_ A_72_1256( .carry(c_72_1256), .sum(s_72_1256), .in3(s_72_1252), .in2(c_71_1225), .in1(s_72_1253) );
  Fadder_ A_72_1257( .carry(c_72_1257), .sum(s_72_1257), .in3(c_71_1226), .in2(s_72_1254), .in1(c_71_1227) );
  Fadder_ A_72_1258( .carry(c_72_1258), .sum(s_72_1258), .in3(s_72_1255), .in2(c_71_1228), .in1(s_72_1256) );
  Fadder_ A_72_1259( .carry(c_72_1259), .sum(s_72_1259), .in3(c_71_1229), .in2(s_72_1257), .in1(c_71_1230) );
  Fadder_ A_72_1260( .carry(c[72]), .sum(s[72]), .in3(s_72_1258), .in2(c_71_1231), .in1(s_72_1259) );

  // ***** Bit 73 ***** //
  Fadder_ A_73_1261( .carry(c_73_1261), .sum(s_73_1261), .in3(P_31[11]), .in2(P_30[13]), .in1(P_29[15]) );
  Fadder_ A_73_1262( .carry(c_73_1262), .sum(s_73_1262), .in3(P_28[17]), .in2(P_27[19]), .in1(P_26[21]) );
  Fadder_ A_73_1263( .carry(c_73_1263), .sum(s_73_1263), .in3(P_25[23]), .in2(P_24[25]), .in1(P_23[27]) );
  Fadder_ A_73_1264( .carry(c_73_1264), .sum(s_73_1264), .in3(P_22[29]), .in2(P_21[31]), .in1(P_20[33]) );
  Fadder_ A_73_1265( .carry(c_73_1265), .sum(s_73_1265), .in3(P_19[35]), .in2(P_18[37]), .in1(P_17[39]) );
  Fadder_ A_73_1266( .carry(c_73_1266), .sum(s_73_1266), .in3(P_16[41]), .in2(P_15[43]), .in1(P_14[45]) );
  Fadder_ A_73_1267( .carry(c_73_1267), .sum(s_73_1267), .in3(P_13[47]), .in2(P_12[49]), .in1(P_11[51]) );
  Fadder_ A_73_1268( .carry(c_73_1268), .sum(s_73_1268), .in3(P_10[53]), .in2(P_9[55]), .in1(P_8[57]) );
  Fadder_ A_73_1269( .carry(c_73_1269), .sum(s_73_1269), .in3(P_7[59]), .in2(P_6[61]), .in1(P_5[63]) );
  Fadder_ A_73_1270( .carry(c_73_1270), .sum(s_73_1270), .in3(P_4[65]), .in2(c_72_1233), .in1(c_72_1242) );
  Fadder_ A_73_1271( .carry(c_73_1271), .sum(s_73_1271), .in3(c_72_1241), .in2(c_72_1240), .in1(c_72_1239) );
  Fadder_ A_73_1272( .carry(c_73_1272), .sum(s_73_1272), .in3(c_72_1238), .in2(c_72_1237), .in1(c_72_1236) );
  Fadder_ A_73_1273( .carry(c_73_1273), .sum(s_73_1273), .in3(c_72_1235), .in2(c_72_1234), .in1(s_73_1269) );
  Fadder_ A_73_1274( .carry(c_73_1274), .sum(s_73_1274), .in3(s_73_1268), .in2(s_73_1267), .in1(s_73_1266) );
  Fadder_ A_73_1275( .carry(c_73_1275), .sum(s_73_1275), .in3(s_73_1265), .in2(s_73_1264), .in1(s_73_1263) );
  Fadder_ A_73_1276( .carry(c_73_1276), .sum(s_73_1276), .in3(s_73_1262), .in2(s_73_1261), .in1(c_72_1245) );
  Fadder_ A_73_1277( .carry(c_73_1277), .sum(s_73_1277), .in3(c_72_1244), .in2(c_72_1243), .in1(s_73_1270) );
  Fadder_ A_73_1278( .carry(c_73_1278), .sum(s_73_1278), .in3(s_73_1272), .in2(s_73_1271), .in1(c_72_1248) );
  Fadder_ A_73_1279( .carry(c_73_1279), .sum(s_73_1279), .in3(c_72_1247), .in2(c_72_1246), .in1(s_73_1273) );
  Fadder_ A_73_1280( .carry(c_73_1280), .sum(s_73_1280), .in3(s_73_1275), .in2(s_73_1274), .in1(c_72_1249) );
  Fadder_ A_73_1281( .carry(c_73_1281), .sum(s_73_1281), .in3(c_72_1250), .in2(s_73_1276), .in1(c_72_1251) );
  Fadder_ A_73_1282( .carry(c_73_1282), .sum(s_73_1282), .in3(c_72_1252), .in2(s_73_1277), .in1(s_73_1278) );
  Fadder_ A_73_1283( .carry(c_73_1283), .sum(s_73_1283), .in3(s_73_1279), .in2(c_72_1253), .in1(s_73_1280) );
  Fadder_ A_73_1284( .carry(c_73_1284), .sum(s_73_1284), .in3(c_72_1254), .in2(s_73_1281), .in1(c_72_1255) );
  Fadder_ A_73_1285( .carry(c_73_1285), .sum(s_73_1285), .in3(s_73_1282), .in2(c_72_1256), .in1(s_73_1283) );
  Fadder_ A_73_1286( .carry(c_73_1286), .sum(s_73_1286), .in3(c_72_1257), .in2(s_73_1284), .in1(c_72_1258) );
  Fadder_ A_73_1287( .carry(c[73]), .sum(s[73]), .in3(s_73_1285), .in2(c_72_1259), .in1(s_73_1286) );

  // ***** Bit 74 ***** //
  Hadder_ A_74_1288( .carry(c_74_1288), .sum(s_74_1288), .in2(sign_), .in1(P_31[12]) );
  Fadder_ A_74_1289( .carry(c_74_1289), .sum(s_74_1289), .in3(P_30[14]), .in2(P_29[16]), .in1(P_28[18]) );
  Fadder_ A_74_1290( .carry(c_74_1290), .sum(s_74_1290), .in3(P_27[20]), .in2(P_26[22]), .in1(P_25[24]) );
  Fadder_ A_74_1291( .carry(c_74_1291), .sum(s_74_1291), .in3(P_24[26]), .in2(P_23[28]), .in1(P_22[30]) );
  Fadder_ A_74_1292( .carry(c_74_1292), .sum(s_74_1292), .in3(P_21[32]), .in2(P_20[34]), .in1(P_19[36]) );
  Fadder_ A_74_1293( .carry(c_74_1293), .sum(s_74_1293), .in3(P_18[38]), .in2(P_17[40]), .in1(P_16[42]) );
  Fadder_ A_74_1294( .carry(c_74_1294), .sum(s_74_1294), .in3(P_15[44]), .in2(P_14[46]), .in1(P_13[48]) );
  Fadder_ A_74_1295( .carry(c_74_1295), .sum(s_74_1295), .in3(P_12[50]), .in2(P_11[52]), .in1(P_10[54]) );
  Fadder_ A_74_1296( .carry(c_74_1296), .sum(s_74_1296), .in3(P_9[56]), .in2(P_8[58]), .in1(P_7[60]) );
  Fadder_ A_74_1297( .carry(c_74_1297), .sum(s_74_1297), .in3(P_6[62]), .in2(P_5[64]), .in1(c_73_1269) );
  Fadder_ A_74_1298( .carry(c_74_1298), .sum(s_74_1298), .in3(c_73_1268), .in2(c_73_1267), .in1(c_73_1266) );
  Fadder_ A_74_1299( .carry(c_74_1299), .sum(s_74_1299), .in3(c_73_1265), .in2(c_73_1264), .in1(c_73_1263) );
  Fadder_ A_74_1300( .carry(c_74_1300), .sum(s_74_1300), .in3(c_73_1262), .in2(c_73_1261), .in1(s_74_1288) );
  Fadder_ A_74_1301( .carry(c_74_1301), .sum(s_74_1301), .in3(s_74_1296), .in2(s_74_1295), .in1(s_74_1294) );
  Fadder_ A_74_1302( .carry(c_74_1302), .sum(s_74_1302), .in3(s_74_1293), .in2(s_74_1292), .in1(s_74_1291) );
  Fadder_ A_74_1303( .carry(c_74_1303), .sum(s_74_1303), .in3(s_74_1290), .in2(s_74_1289), .in1(c_73_1270) );
  Fadder_ A_74_1304( .carry(c_74_1304), .sum(s_74_1304), .in3(c_73_1272), .in2(c_73_1271), .in1(c_73_1273) );
  Fadder_ A_74_1305( .carry(c_74_1305), .sum(s_74_1305), .in3(s_74_1297), .in2(s_74_1299), .in1(s_74_1298) );
  Fadder_ A_74_1306( .carry(c_74_1306), .sum(s_74_1306), .in3(c_73_1275), .in2(c_73_1274), .in1(s_74_1300) );
  Fadder_ A_74_1307( .carry(c_74_1307), .sum(s_74_1307), .in3(s_74_1302), .in2(s_74_1301), .in1(c_73_1276) );
  Fadder_ A_74_1308( .carry(c_74_1308), .sum(s_74_1308), .in3(s_74_1303), .in2(c_73_1277), .in1(c_73_1278) );
  Fadder_ A_74_1309( .carry(c_74_1309), .sum(s_74_1309), .in3(s_74_1304), .in2(c_73_1279), .in1(s_74_1305) );
  Fadder_ A_74_1310( .carry(c_74_1310), .sum(s_74_1310), .in3(s_74_1306), .in2(c_73_1280), .in1(s_74_1307) );
  Fadder_ A_74_1311( .carry(c_74_1311), .sum(s_74_1311), .in3(c_73_1281), .in2(c_73_1282), .in1(s_74_1308) );
  Fadder_ A_74_1312( .carry(c_74_1312), .sum(s_74_1312), .in3(s_74_1309), .in2(c_73_1283), .in1(s_74_1310) );
  Fadder_ A_74_1313( .carry(c_74_1313), .sum(s_74_1313), .in3(c_73_1284), .in2(s_74_1311), .in1(c_73_1285) );
  Fadder_ A_74_1314( .carry(c[74]), .sum(s[74]), .in3(s_74_1312), .in2(c_73_1286), .in1(s_74_1313) );

  // ***** Bit 75 ***** //
  Fadder_ A_75_1315( .carry(c_75_1315), .sum(s_75_1315), .in3(P_31[13]), .in2(P_30[15]), .in1(P_29[17]) );
  Fadder_ A_75_1316( .carry(c_75_1316), .sum(s_75_1316), .in3(P_28[19]), .in2(P_27[21]), .in1(P_26[23]) );
  Fadder_ A_75_1317( .carry(c_75_1317), .sum(s_75_1317), .in3(P_25[25]), .in2(P_24[27]), .in1(P_23[29]) );
  Fadder_ A_75_1318( .carry(c_75_1318), .sum(s_75_1318), .in3(P_22[31]), .in2(P_21[33]), .in1(P_20[35]) );
  Fadder_ A_75_1319( .carry(c_75_1319), .sum(s_75_1319), .in3(P_19[37]), .in2(P_18[39]), .in1(P_17[41]) );
  Fadder_ A_75_1320( .carry(c_75_1320), .sum(s_75_1320), .in3(P_16[43]), .in2(P_15[45]), .in1(P_14[47]) );
  Fadder_ A_75_1321( .carry(c_75_1321), .sum(s_75_1321), .in3(P_13[49]), .in2(P_12[51]), .in1(P_11[53]) );
  Fadder_ A_75_1322( .carry(c_75_1322), .sum(s_75_1322), .in3(P_10[55]), .in2(P_9[57]), .in1(P_8[59]) );
  Fadder_ A_75_1323( .carry(c_75_1323), .sum(s_75_1323), .in3(P_7[61]), .in2(P_6[63]), .in1(P_5[65]) );
  Fadder_ A_75_1324( .carry(c_75_1324), .sum(s_75_1324), .in3(c_74_1288), .in2(c_74_1296), .in1(c_74_1295) );
  Fadder_ A_75_1325( .carry(c_75_1325), .sum(s_75_1325), .in3(c_74_1294), .in2(c_74_1293), .in1(c_74_1292) );
  Fadder_ A_75_1326( .carry(c_75_1326), .sum(s_75_1326), .in3(c_74_1291), .in2(c_74_1290), .in1(c_74_1289) );
  Fadder_ A_75_1327( .carry(c_75_1327), .sum(s_75_1327), .in3(s_75_1323), .in2(s_75_1322), .in1(s_75_1321) );
  Fadder_ A_75_1328( .carry(c_75_1328), .sum(s_75_1328), .in3(s_75_1320), .in2(s_75_1319), .in1(s_75_1318) );
  Fadder_ A_75_1329( .carry(c_75_1329), .sum(s_75_1329), .in3(s_75_1317), .in2(s_75_1316), .in1(s_75_1315) );
  Fadder_ A_75_1330( .carry(c_75_1330), .sum(s_75_1330), .in3(c_74_1297), .in2(c_74_1300), .in1(c_74_1299) );
  Fadder_ A_75_1331( .carry(c_75_1331), .sum(s_75_1331), .in3(c_74_1298), .in2(s_75_1324), .in1(s_75_1326) );
  Fadder_ A_75_1332( .carry(c_75_1332), .sum(s_75_1332), .in3(s_75_1325), .in2(c_74_1302), .in1(c_74_1301) );
  Fadder_ A_75_1333( .carry(c_75_1333), .sum(s_75_1333), .in3(s_75_1329), .in2(s_75_1328), .in1(s_75_1327) );
  Fadder_ A_75_1334( .carry(c_75_1334), .sum(s_75_1334), .in3(c_74_1303), .in2(c_74_1304), .in1(s_75_1330) );
  Fadder_ A_75_1335( .carry(c_75_1335), .sum(s_75_1335), .in3(c_74_1306), .in2(c_74_1305), .in1(s_75_1331) );
  Fadder_ A_75_1336( .carry(c_75_1336), .sum(s_75_1336), .in3(s_75_1332), .in2(s_75_1333), .in1(c_74_1307) );
  Fadder_ A_75_1337( .carry(c_75_1337), .sum(s_75_1337), .in3(c_74_1308), .in2(c_74_1309), .in1(s_75_1334) );
  Fadder_ A_75_1338( .carry(c_75_1338), .sum(s_75_1338), .in3(s_75_1335), .in2(s_75_1336), .in1(c_74_1310) );
  Fadder_ A_75_1339( .carry(c_75_1339), .sum(s_75_1339), .in3(c_74_1311), .in2(s_75_1337), .in1(c_74_1312) );
  Fadder_ A_75_1340( .carry(c[75]), .sum(s[75]), .in3(s_75_1338), .in2(c_74_1313), .in1(s_75_1339) );

  // ***** Bit 76 ***** //
  Hadder_ A_76_1341( .carry(c_76_1341), .sum(s_76_1341), .in2(sign_), .in1(P_31[14]) );
  Fadder_ A_76_1342( .carry(c_76_1342), .sum(s_76_1342), .in3(P_30[16]), .in2(P_29[18]), .in1(P_28[20]) );
  Fadder_ A_76_1343( .carry(c_76_1343), .sum(s_76_1343), .in3(P_27[22]), .in2(P_26[24]), .in1(P_25[26]) );
  Fadder_ A_76_1344( .carry(c_76_1344), .sum(s_76_1344), .in3(P_24[28]), .in2(P_23[30]), .in1(P_22[32]) );
  Fadder_ A_76_1345( .carry(c_76_1345), .sum(s_76_1345), .in3(P_21[34]), .in2(P_20[36]), .in1(P_19[38]) );
  Fadder_ A_76_1346( .carry(c_76_1346), .sum(s_76_1346), .in3(P_18[40]), .in2(P_17[42]), .in1(P_16[44]) );
  Fadder_ A_76_1347( .carry(c_76_1347), .sum(s_76_1347), .in3(P_15[46]), .in2(P_14[48]), .in1(P_13[50]) );
  Fadder_ A_76_1348( .carry(c_76_1348), .sum(s_76_1348), .in3(P_12[52]), .in2(P_11[54]), .in1(P_10[56]) );
  Fadder_ A_76_1349( .carry(c_76_1349), .sum(s_76_1349), .in3(P_9[58]), .in2(P_8[60]), .in1(P_7[62]) );
  Fadder_ A_76_1350( .carry(c_76_1350), .sum(s_76_1350), .in3(P_6[64]), .in2(c_75_1323), .in1(c_75_1322) );
  Fadder_ A_76_1351( .carry(c_76_1351), .sum(s_76_1351), .in3(c_75_1321), .in2(c_75_1320), .in1(c_75_1319) );
  Fadder_ A_76_1352( .carry(c_76_1352), .sum(s_76_1352), .in3(c_75_1318), .in2(c_75_1317), .in1(c_75_1316) );
  Fadder_ A_76_1353( .carry(c_76_1353), .sum(s_76_1353), .in3(c_75_1315), .in2(s_76_1341), .in1(s_76_1349) );
  Fadder_ A_76_1354( .carry(c_76_1354), .sum(s_76_1354), .in3(s_76_1348), .in2(s_76_1347), .in1(s_76_1346) );
  Fadder_ A_76_1355( .carry(c_76_1355), .sum(s_76_1355), .in3(s_76_1345), .in2(s_76_1344), .in1(s_76_1343) );
  Fadder_ A_76_1356( .carry(c_76_1356), .sum(s_76_1356), .in3(s_76_1342), .in2(c_75_1326), .in1(c_75_1325) );
  Fadder_ A_76_1357( .carry(c_76_1357), .sum(s_76_1357), .in3(c_75_1324), .in2(s_76_1350), .in1(s_76_1352) );
  Fadder_ A_76_1358( .carry(c_76_1358), .sum(s_76_1358), .in3(s_76_1351), .in2(c_75_1329), .in1(c_75_1328) );
  Fadder_ A_76_1359( .carry(c_76_1359), .sum(s_76_1359), .in3(c_75_1327), .in2(s_76_1353), .in1(s_76_1355) );
  Fadder_ A_76_1360( .carry(c_76_1360), .sum(s_76_1360), .in3(s_76_1354), .in2(c_75_1330), .in1(s_76_1356) );
  Fadder_ A_76_1361( .carry(c_76_1361), .sum(s_76_1361), .in3(c_75_1331), .in2(c_75_1332), .in1(s_76_1357) );
  Fadder_ A_76_1362( .carry(c_76_1362), .sum(s_76_1362), .in3(s_76_1358), .in2(c_75_1333), .in1(s_76_1359) );
  Fadder_ A_76_1363( .carry(c_76_1363), .sum(s_76_1363), .in3(c_75_1334), .in2(c_75_1335), .in1(s_76_1360) );
  Fadder_ A_76_1364( .carry(c_76_1364), .sum(s_76_1364), .in3(s_76_1361), .in2(c_75_1336), .in1(s_76_1362) );
  Fadder_ A_76_1365( .carry(c_76_1365), .sum(s_76_1365), .in3(c_75_1337), .in2(s_76_1363), .in1(c_75_1338) );
  Fadder_ A_76_1366( .carry(c[76]), .sum(s[76]), .in3(s_76_1364), .in2(c_75_1339), .in1(s_76_1365) );

  // ***** Bit 77 ***** //
  Fadder_ A_77_1367( .carry(c_77_1367), .sum(s_77_1367), .in3(P_31[15]), .in2(P_30[17]), .in1(P_29[19]) );
  Fadder_ A_77_1368( .carry(c_77_1368), .sum(s_77_1368), .in3(P_28[21]), .in2(P_27[23]), .in1(P_26[25]) );
  Fadder_ A_77_1369( .carry(c_77_1369), .sum(s_77_1369), .in3(P_25[27]), .in2(P_24[29]), .in1(P_23[31]) );
  Fadder_ A_77_1370( .carry(c_77_1370), .sum(s_77_1370), .in3(P_22[33]), .in2(P_21[35]), .in1(P_20[37]) );
  Fadder_ A_77_1371( .carry(c_77_1371), .sum(s_77_1371), .in3(P_19[39]), .in2(P_18[41]), .in1(P_17[43]) );
  Fadder_ A_77_1372( .carry(c_77_1372), .sum(s_77_1372), .in3(P_16[45]), .in2(P_15[47]), .in1(P_14[49]) );
  Fadder_ A_77_1373( .carry(c_77_1373), .sum(s_77_1373), .in3(P_13[51]), .in2(P_12[53]), .in1(P_11[55]) );
  Fadder_ A_77_1374( .carry(c_77_1374), .sum(s_77_1374), .in3(P_10[57]), .in2(P_9[59]), .in1(P_8[61]) );
  Fadder_ A_77_1375( .carry(c_77_1375), .sum(s_77_1375), .in3(P_7[63]), .in2(P_6[65]), .in1(c_76_1341) );
  Fadder_ A_77_1376( .carry(c_77_1376), .sum(s_77_1376), .in3(c_76_1349), .in2(c_76_1348), .in1(c_76_1347) );
  Fadder_ A_77_1377( .carry(c_77_1377), .sum(s_77_1377), .in3(c_76_1346), .in2(c_76_1345), .in1(c_76_1344) );
  Fadder_ A_77_1378( .carry(c_77_1378), .sum(s_77_1378), .in3(c_76_1343), .in2(c_76_1342), .in1(s_77_1374) );
  Fadder_ A_77_1379( .carry(c_77_1379), .sum(s_77_1379), .in3(s_77_1373), .in2(s_77_1372), .in1(s_77_1371) );
  Fadder_ A_77_1380( .carry(c_77_1380), .sum(s_77_1380), .in3(s_77_1370), .in2(s_77_1369), .in1(s_77_1368) );
  Fadder_ A_77_1381( .carry(c_77_1381), .sum(s_77_1381), .in3(s_77_1367), .in2(s_77_1375), .in1(c_76_1352) );
  Fadder_ A_77_1382( .carry(c_77_1382), .sum(s_77_1382), .in3(c_76_1351), .in2(c_76_1350), .in1(c_76_1353) );
  Fadder_ A_77_1383( .carry(c_77_1383), .sum(s_77_1383), .in3(s_77_1377), .in2(s_77_1376), .in1(c_76_1355) );
  Fadder_ A_77_1384( .carry(c_77_1384), .sum(s_77_1384), .in3(c_76_1354), .in2(s_77_1378), .in1(s_77_1380) );
  Fadder_ A_77_1385( .carry(c_77_1385), .sum(s_77_1385), .in3(s_77_1379), .in2(c_76_1356), .in1(s_77_1381) );
  Fadder_ A_77_1386( .carry(c_77_1386), .sum(s_77_1386), .in3(c_76_1357), .in2(c_76_1358), .in1(s_77_1382) );
  Fadder_ A_77_1387( .carry(c_77_1387), .sum(s_77_1387), .in3(c_76_1359), .in2(s_77_1383), .in1(s_77_1384) );
  Fadder_ A_77_1388( .carry(c_77_1388), .sum(s_77_1388), .in3(c_76_1360), .in2(c_76_1361), .in1(s_77_1385) );
  Fadder_ A_77_1389( .carry(c_77_1389), .sum(s_77_1389), .in3(s_77_1386), .in2(c_76_1362), .in1(s_77_1387) );
  Fadder_ A_77_1390( .carry(c_77_1390), .sum(s_77_1390), .in3(c_76_1363), .in2(s_77_1388), .in1(c_76_1364) );
  Fadder_ A_77_1391( .carry(c[77]), .sum(s[77]), .in3(s_77_1389), .in2(c_76_1365), .in1(s_77_1390) );

  // ***** Bit 78 ***** //
  Hadder_ A_78_1392( .carry(c_78_1392), .sum(s_78_1392), .in2(sign_), .in1(P_31[16]) );
  Fadder_ A_78_1393( .carry(c_78_1393), .sum(s_78_1393), .in3(P_30[18]), .in2(P_29[20]), .in1(P_28[22]) );
  Fadder_ A_78_1394( .carry(c_78_1394), .sum(s_78_1394), .in3(P_27[24]), .in2(P_26[26]), .in1(P_25[28]) );
  Fadder_ A_78_1395( .carry(c_78_1395), .sum(s_78_1395), .in3(P_24[30]), .in2(P_23[32]), .in1(P_22[34]) );
  Fadder_ A_78_1396( .carry(c_78_1396), .sum(s_78_1396), .in3(P_21[36]), .in2(P_20[38]), .in1(P_19[40]) );
  Fadder_ A_78_1397( .carry(c_78_1397), .sum(s_78_1397), .in3(P_18[42]), .in2(P_17[44]), .in1(P_16[46]) );
  Fadder_ A_78_1398( .carry(c_78_1398), .sum(s_78_1398), .in3(P_15[48]), .in2(P_14[50]), .in1(P_13[52]) );
  Fadder_ A_78_1399( .carry(c_78_1399), .sum(s_78_1399), .in3(P_12[54]), .in2(P_11[56]), .in1(P_10[58]) );
  Fadder_ A_78_1400( .carry(c_78_1400), .sum(s_78_1400), .in3(P_9[60]), .in2(P_8[62]), .in1(P_7[64]) );
  Fadder_ A_78_1401( .carry(c_78_1401), .sum(s_78_1401), .in3(c_77_1374), .in2(c_77_1373), .in1(c_77_1372) );
  Fadder_ A_78_1402( .carry(c_78_1402), .sum(s_78_1402), .in3(c_77_1371), .in2(c_77_1370), .in1(c_77_1369) );
  Fadder_ A_78_1403( .carry(c_78_1403), .sum(s_78_1403), .in3(c_77_1368), .in2(c_77_1367), .in1(s_78_1392) );
  Fadder_ A_78_1404( .carry(c_78_1404), .sum(s_78_1404), .in3(s_78_1400), .in2(s_78_1399), .in1(s_78_1398) );
  Fadder_ A_78_1405( .carry(c_78_1405), .sum(s_78_1405), .in3(s_78_1397), .in2(s_78_1396), .in1(s_78_1395) );
  Fadder_ A_78_1406( .carry(c_78_1406), .sum(s_78_1406), .in3(s_78_1394), .in2(s_78_1393), .in1(c_77_1375) );
  Fadder_ A_78_1407( .carry(c_78_1407), .sum(s_78_1407), .in3(c_77_1377), .in2(c_77_1376), .in1(c_77_1378) );
  Fadder_ A_78_1408( .carry(c_78_1408), .sum(s_78_1408), .in3(s_78_1402), .in2(s_78_1401), .in1(c_77_1380) );
  Fadder_ A_78_1409( .carry(c_78_1409), .sum(s_78_1409), .in3(c_77_1379), .in2(s_78_1403), .in1(s_78_1405) );
  Fadder_ A_78_1410( .carry(c_78_1410), .sum(s_78_1410), .in3(s_78_1404), .in2(s_78_1406), .in1(c_77_1381) );
  Fadder_ A_78_1411( .carry(c_78_1411), .sum(s_78_1411), .in3(c_77_1382), .in2(c_77_1383), .in1(s_78_1407) );
  Fadder_ A_78_1412( .carry(c_78_1412), .sum(s_78_1412), .in3(c_77_1384), .in2(s_78_1408), .in1(s_78_1409) );
  Fadder_ A_78_1413( .carry(c_78_1413), .sum(s_78_1413), .in3(s_78_1410), .in2(c_77_1385), .in1(c_77_1386) );
  Fadder_ A_78_1414( .carry(c_78_1414), .sum(s_78_1414), .in3(s_78_1411), .in2(c_77_1387), .in1(s_78_1412) );
  Fadder_ A_78_1415( .carry(c_78_1415), .sum(s_78_1415), .in3(c_77_1388), .in2(s_78_1413), .in1(c_77_1389) );
  Fadder_ A_78_1416( .carry(c[78]), .sum(s[78]), .in3(s_78_1414), .in2(c_77_1390), .in1(s_78_1415) );

  // ***** Bit 79 ***** //
  Fadder_ A_79_1417( .carry(c_79_1417), .sum(s_79_1417), .in3(P_31[17]), .in2(P_30[19]), .in1(P_29[21]) );
  Fadder_ A_79_1418( .carry(c_79_1418), .sum(s_79_1418), .in3(P_28[23]), .in2(P_27[25]), .in1(P_26[27]) );
  Fadder_ A_79_1419( .carry(c_79_1419), .sum(s_79_1419), .in3(P_25[29]), .in2(P_24[31]), .in1(P_23[33]) );
  Fadder_ A_79_1420( .carry(c_79_1420), .sum(s_79_1420), .in3(P_22[35]), .in2(P_21[37]), .in1(P_20[39]) );
  Fadder_ A_79_1421( .carry(c_79_1421), .sum(s_79_1421), .in3(P_19[41]), .in2(P_18[43]), .in1(P_17[45]) );
  Fadder_ A_79_1422( .carry(c_79_1422), .sum(s_79_1422), .in3(P_16[47]), .in2(P_15[49]), .in1(P_14[51]) );
  Fadder_ A_79_1423( .carry(c_79_1423), .sum(s_79_1423), .in3(P_13[53]), .in2(P_12[55]), .in1(P_11[57]) );
  Fadder_ A_79_1424( .carry(c_79_1424), .sum(s_79_1424), .in3(P_10[59]), .in2(P_9[61]), .in1(P_8[63]) );
  Fadder_ A_79_1425( .carry(c_79_1425), .sum(s_79_1425), .in3(P_7[65]), .in2(c_78_1392), .in1(c_78_1400) );
  Fadder_ A_79_1426( .carry(c_79_1426), .sum(s_79_1426), .in3(c_78_1399), .in2(c_78_1398), .in1(c_78_1397) );
  Fadder_ A_79_1427( .carry(c_79_1427), .sum(s_79_1427), .in3(c_78_1396), .in2(c_78_1395), .in1(c_78_1394) );
  Fadder_ A_79_1428( .carry(c_79_1428), .sum(s_79_1428), .in3(c_78_1393), .in2(s_79_1424), .in1(s_79_1423) );
  Fadder_ A_79_1429( .carry(c_79_1429), .sum(s_79_1429), .in3(s_79_1422), .in2(s_79_1421), .in1(s_79_1420) );
  Fadder_ A_79_1430( .carry(c_79_1430), .sum(s_79_1430), .in3(s_79_1419), .in2(s_79_1418), .in1(s_79_1417) );
  Fadder_ A_79_1431( .carry(c_79_1431), .sum(s_79_1431), .in3(c_78_1403), .in2(c_78_1402), .in1(c_78_1401) );
  Fadder_ A_79_1432( .carry(c_79_1432), .sum(s_79_1432), .in3(s_79_1425), .in2(s_79_1427), .in1(s_79_1426) );
  Fadder_ A_79_1433( .carry(c_79_1433), .sum(s_79_1433), .in3(c_78_1405), .in2(c_78_1404), .in1(c_78_1406) );
  Fadder_ A_79_1434( .carry(c_79_1434), .sum(s_79_1434), .in3(s_79_1428), .in2(s_79_1430), .in1(s_79_1429) );
  Fadder_ A_79_1435( .carry(c_79_1435), .sum(s_79_1435), .in3(c_78_1407), .in2(s_79_1431), .in1(c_78_1408) );
  Fadder_ A_79_1436( .carry(c_79_1436), .sum(s_79_1436), .in3(c_78_1409), .in2(s_79_1432), .in1(s_79_1433) );
  Fadder_ A_79_1437( .carry(c_79_1437), .sum(s_79_1437), .in3(s_79_1434), .in2(c_78_1410), .in1(c_78_1411) );
  Fadder_ A_79_1438( .carry(c_79_1438), .sum(s_79_1438), .in3(s_79_1435), .in2(c_78_1412), .in1(s_79_1436) );
  Fadder_ A_79_1439( .carry(c_79_1439), .sum(s_79_1439), .in3(c_78_1413), .in2(s_79_1437), .in1(c_78_1414) );
  Fadder_ A_79_1440( .carry(c[79]), .sum(s[79]), .in3(s_79_1438), .in2(c_78_1415), .in1(s_79_1439) );

  // ***** Bit 80 ***** //
  Hadder_ A_80_1441( .carry(c_80_1441), .sum(s_80_1441), .in2(sign_), .in1(P_31[18]) );
  Fadder_ A_80_1442( .carry(c_80_1442), .sum(s_80_1442), .in3(P_30[20]), .in2(P_29[22]), .in1(P_28[24]) );
  Fadder_ A_80_1443( .carry(c_80_1443), .sum(s_80_1443), .in3(P_27[26]), .in2(P_26[28]), .in1(P_25[30]) );
  Fadder_ A_80_1444( .carry(c_80_1444), .sum(s_80_1444), .in3(P_24[32]), .in2(P_23[34]), .in1(P_22[36]) );
  Fadder_ A_80_1445( .carry(c_80_1445), .sum(s_80_1445), .in3(P_21[38]), .in2(P_20[40]), .in1(P_19[42]) );
  Fadder_ A_80_1446( .carry(c_80_1446), .sum(s_80_1446), .in3(P_18[44]), .in2(P_17[46]), .in1(P_16[48]) );
  Fadder_ A_80_1447( .carry(c_80_1447), .sum(s_80_1447), .in3(P_15[50]), .in2(P_14[52]), .in1(P_13[54]) );
  Fadder_ A_80_1448( .carry(c_80_1448), .sum(s_80_1448), .in3(P_12[56]), .in2(P_11[58]), .in1(P_10[60]) );
  Fadder_ A_80_1449( .carry(c_80_1449), .sum(s_80_1449), .in3(P_9[62]), .in2(P_8[64]), .in1(c_79_1424) );
  Fadder_ A_80_1450( .carry(c_80_1450), .sum(s_80_1450), .in3(c_79_1423), .in2(c_79_1422), .in1(c_79_1421) );
  Fadder_ A_80_1451( .carry(c_80_1451), .sum(s_80_1451), .in3(c_79_1420), .in2(c_79_1419), .in1(c_79_1418) );
  Fadder_ A_80_1452( .carry(c_80_1452), .sum(s_80_1452), .in3(c_79_1417), .in2(s_80_1441), .in1(s_80_1448) );
  Fadder_ A_80_1453( .carry(c_80_1453), .sum(s_80_1453), .in3(s_80_1447), .in2(s_80_1446), .in1(s_80_1445) );
  Fadder_ A_80_1454( .carry(c_80_1454), .sum(s_80_1454), .in3(s_80_1444), .in2(s_80_1443), .in1(s_80_1442) );
  Fadder_ A_80_1455( .carry(c_80_1455), .sum(s_80_1455), .in3(c_79_1425), .in2(c_79_1427), .in1(c_79_1426) );
  Fadder_ A_80_1456( .carry(c_80_1456), .sum(s_80_1456), .in3(s_80_1449), .in2(s_80_1451), .in1(s_80_1450) );
  Fadder_ A_80_1457( .carry(c_80_1457), .sum(s_80_1457), .in3(c_79_1430), .in2(c_79_1429), .in1(c_79_1428) );
  Fadder_ A_80_1458( .carry(c_80_1458), .sum(s_80_1458), .in3(s_80_1452), .in2(s_80_1454), .in1(s_80_1453) );
  Fadder_ A_80_1459( .carry(c_80_1459), .sum(s_80_1459), .in3(c_79_1431), .in2(s_80_1455), .in1(c_79_1433) );
  Fadder_ A_80_1460( .carry(c_80_1460), .sum(s_80_1460), .in3(c_79_1432), .in2(s_80_1456), .in1(s_80_1457) );
  Fadder_ A_80_1461( .carry(c_80_1461), .sum(s_80_1461), .in3(c_79_1434), .in2(s_80_1458), .in1(c_79_1435) );
  Fadder_ A_80_1462( .carry(c_80_1462), .sum(s_80_1462), .in3(s_80_1459), .in2(c_79_1436), .in1(s_80_1460) );
  Fadder_ A_80_1463( .carry(c_80_1463), .sum(s_80_1463), .in3(c_79_1437), .in2(s_80_1461), .in1(c_79_1438) );
  Fadder_ A_80_1464( .carry(c[80]), .sum(s[80]), .in3(s_80_1462), .in2(c_79_1439), .in1(s_80_1463) );

  // ***** Bit 81 ***** //
  Fadder_ A_81_1465( .carry(c_81_1465), .sum(s_81_1465), .in3(P_31[19]), .in2(P_30[21]), .in1(P_29[23]) );
  Fadder_ A_81_1466( .carry(c_81_1466), .sum(s_81_1466), .in3(P_28[25]), .in2(P_27[27]), .in1(P_26[29]) );
  Fadder_ A_81_1467( .carry(c_81_1467), .sum(s_81_1467), .in3(P_25[31]), .in2(P_24[33]), .in1(P_23[35]) );
  Fadder_ A_81_1468( .carry(c_81_1468), .sum(s_81_1468), .in3(P_22[37]), .in2(P_21[39]), .in1(P_20[41]) );
  Fadder_ A_81_1469( .carry(c_81_1469), .sum(s_81_1469), .in3(P_19[43]), .in2(P_18[45]), .in1(P_17[47]) );
  Fadder_ A_81_1470( .carry(c_81_1470), .sum(s_81_1470), .in3(P_16[49]), .in2(P_15[51]), .in1(P_14[53]) );
  Fadder_ A_81_1471( .carry(c_81_1471), .sum(s_81_1471), .in3(P_13[55]), .in2(P_12[57]), .in1(P_11[59]) );
  Fadder_ A_81_1472( .carry(c_81_1472), .sum(s_81_1472), .in3(P_10[61]), .in2(P_9[63]), .in1(P_8[65]) );
  Fadder_ A_81_1473( .carry(c_81_1473), .sum(s_81_1473), .in3(c_80_1441), .in2(c_80_1448), .in1(c_80_1447) );
  Fadder_ A_81_1474( .carry(c_81_1474), .sum(s_81_1474), .in3(c_80_1446), .in2(c_80_1445), .in1(c_80_1444) );
  Fadder_ A_81_1475( .carry(c_81_1475), .sum(s_81_1475), .in3(c_80_1443), .in2(c_80_1442), .in1(s_81_1472) );
  Fadder_ A_81_1476( .carry(c_81_1476), .sum(s_81_1476), .in3(s_81_1471), .in2(s_81_1470), .in1(s_81_1469) );
  Fadder_ A_81_1477( .carry(c_81_1477), .sum(s_81_1477), .in3(s_81_1468), .in2(s_81_1467), .in1(s_81_1466) );
  Fadder_ A_81_1478( .carry(c_81_1478), .sum(s_81_1478), .in3(s_81_1465), .in2(c_80_1449), .in1(c_80_1451) );
  Fadder_ A_81_1479( .carry(c_81_1479), .sum(s_81_1479), .in3(c_80_1450), .in2(c_80_1452), .in1(s_81_1473) );
  Fadder_ A_81_1480( .carry(c_81_1480), .sum(s_81_1480), .in3(s_81_1474), .in2(c_80_1454), .in1(c_80_1453) );
  Fadder_ A_81_1481( .carry(c_81_1481), .sum(s_81_1481), .in3(s_81_1475), .in2(s_81_1477), .in1(s_81_1476) );
  Fadder_ A_81_1482( .carry(c_81_1482), .sum(s_81_1482), .in3(c_80_1455), .in2(s_81_1478), .in1(c_80_1457) );
  Fadder_ A_81_1483( .carry(c_81_1483), .sum(s_81_1483), .in3(c_80_1456), .in2(s_81_1479), .in1(s_81_1480) );
  Fadder_ A_81_1484( .carry(c_81_1484), .sum(s_81_1484), .in3(c_80_1458), .in2(s_81_1481), .in1(c_80_1459) );
  Fadder_ A_81_1485( .carry(c_81_1485), .sum(s_81_1485), .in3(s_81_1482), .in2(c_80_1460), .in1(s_81_1483) );
  Fadder_ A_81_1486( .carry(c_81_1486), .sum(s_81_1486), .in3(c_80_1461), .in2(s_81_1484), .in1(c_80_1462) );
  Fadder_ A_81_1487( .carry(c[81]), .sum(s[81]), .in3(s_81_1485), .in2(c_80_1463), .in1(s_81_1486) );

  // ***** Bit 82 ***** //
  Hadder_ A_82_1488( .carry(c_82_1488), .sum(s_82_1488), .in2(sign_), .in1(P_31[20]) );
  Fadder_ A_82_1489( .carry(c_82_1489), .sum(s_82_1489), .in3(P_30[22]), .in2(P_29[24]), .in1(P_28[26]) );
  Fadder_ A_82_1490( .carry(c_82_1490), .sum(s_82_1490), .in3(P_27[28]), .in2(P_26[30]), .in1(P_25[32]) );
  Fadder_ A_82_1491( .carry(c_82_1491), .sum(s_82_1491), .in3(P_24[34]), .in2(P_23[36]), .in1(P_22[38]) );
  Fadder_ A_82_1492( .carry(c_82_1492), .sum(s_82_1492), .in3(P_21[40]), .in2(P_20[42]), .in1(P_19[44]) );
  Fadder_ A_82_1493( .carry(c_82_1493), .sum(s_82_1493), .in3(P_18[46]), .in2(P_17[48]), .in1(P_16[50]) );
  Fadder_ A_82_1494( .carry(c_82_1494), .sum(s_82_1494), .in3(P_15[52]), .in2(P_14[54]), .in1(P_13[56]) );
  Fadder_ A_82_1495( .carry(c_82_1495), .sum(s_82_1495), .in3(P_12[58]), .in2(P_11[60]), .in1(P_10[62]) );
  Fadder_ A_82_1496( .carry(c_82_1496), .sum(s_82_1496), .in3(P_9[64]), .in2(c_81_1472), .in1(c_81_1471) );
  Fadder_ A_82_1497( .carry(c_82_1497), .sum(s_82_1497), .in3(c_81_1470), .in2(c_81_1469), .in1(c_81_1468) );
  Fadder_ A_82_1498( .carry(c_82_1498), .sum(s_82_1498), .in3(c_81_1467), .in2(c_81_1466), .in1(c_81_1465) );
  Fadder_ A_82_1499( .carry(c_82_1499), .sum(s_82_1499), .in3(s_82_1488), .in2(s_82_1495), .in1(s_82_1494) );
  Fadder_ A_82_1500( .carry(c_82_1500), .sum(s_82_1500), .in3(s_82_1493), .in2(s_82_1492), .in1(s_82_1491) );
  Fadder_ A_82_1501( .carry(c_82_1501), .sum(s_82_1501), .in3(s_82_1490), .in2(s_82_1489), .in1(c_81_1474) );
  Fadder_ A_82_1502( .carry(c_82_1502), .sum(s_82_1502), .in3(c_81_1473), .in2(c_81_1475), .in1(s_82_1496) );
  Fadder_ A_82_1503( .carry(c_82_1503), .sum(s_82_1503), .in3(s_82_1498), .in2(s_82_1497), .in1(c_81_1477) );
  Fadder_ A_82_1504( .carry(c_82_1504), .sum(s_82_1504), .in3(c_81_1476), .in2(s_82_1499), .in1(s_82_1500) );
  Fadder_ A_82_1505( .carry(c_82_1505), .sum(s_82_1505), .in3(c_81_1478), .in2(c_81_1479), .in1(s_82_1501) );
  Fadder_ A_82_1506( .carry(c_82_1506), .sum(s_82_1506), .in3(c_81_1480), .in2(s_82_1502), .in1(s_82_1503) );
  Fadder_ A_82_1507( .carry(c_82_1507), .sum(s_82_1507), .in3(c_81_1481), .in2(s_82_1504), .in1(c_81_1482) );
  Fadder_ A_82_1508( .carry(c_82_1508), .sum(s_82_1508), .in3(s_82_1505), .in2(c_81_1483), .in1(s_82_1506) );
  Fadder_ A_82_1509( .carry(c_82_1509), .sum(s_82_1509), .in3(c_81_1484), .in2(s_82_1507), .in1(c_81_1485) );
  Fadder_ A_82_1510( .carry(c[82]), .sum(s[82]), .in3(s_82_1508), .in2(c_81_1486), .in1(s_82_1509) );

  // ***** Bit 83 ***** //
  Fadder_ A_83_1511( .carry(c_83_1511), .sum(s_83_1511), .in3(P_31[21]), .in2(P_30[23]), .in1(P_29[25]) );
  Fadder_ A_83_1512( .carry(c_83_1512), .sum(s_83_1512), .in3(P_28[27]), .in2(P_27[29]), .in1(P_26[31]) );
  Fadder_ A_83_1513( .carry(c_83_1513), .sum(s_83_1513), .in3(P_25[33]), .in2(P_24[35]), .in1(P_23[37]) );
  Fadder_ A_83_1514( .carry(c_83_1514), .sum(s_83_1514), .in3(P_22[39]), .in2(P_21[41]), .in1(P_20[43]) );
  Fadder_ A_83_1515( .carry(c_83_1515), .sum(s_83_1515), .in3(P_19[45]), .in2(P_18[47]), .in1(P_17[49]) );
  Fadder_ A_83_1516( .carry(c_83_1516), .sum(s_83_1516), .in3(P_16[51]), .in2(P_15[53]), .in1(P_14[55]) );
  Fadder_ A_83_1517( .carry(c_83_1517), .sum(s_83_1517), .in3(P_13[57]), .in2(P_12[59]), .in1(P_11[61]) );
  Fadder_ A_83_1518( .carry(c_83_1518), .sum(s_83_1518), .in3(P_10[63]), .in2(P_9[65]), .in1(c_82_1488) );
  Fadder_ A_83_1519( .carry(c_83_1519), .sum(s_83_1519), .in3(c_82_1495), .in2(c_82_1494), .in1(c_82_1493) );
  Fadder_ A_83_1520( .carry(c_83_1520), .sum(s_83_1520), .in3(c_82_1492), .in2(c_82_1491), .in1(c_82_1490) );
  Fadder_ A_83_1521( .carry(c_83_1521), .sum(s_83_1521), .in3(c_82_1489), .in2(s_83_1517), .in1(s_83_1516) );
  Fadder_ A_83_1522( .carry(c_83_1522), .sum(s_83_1522), .in3(s_83_1515), .in2(s_83_1514), .in1(s_83_1513) );
  Fadder_ A_83_1523( .carry(c_83_1523), .sum(s_83_1523), .in3(s_83_1512), .in2(s_83_1511), .in1(s_83_1518) );
  Fadder_ A_83_1524( .carry(c_83_1524), .sum(s_83_1524), .in3(c_82_1498), .in2(c_82_1497), .in1(c_82_1496) );
  Fadder_ A_83_1525( .carry(c_83_1525), .sum(s_83_1525), .in3(s_83_1520), .in2(s_83_1519), .in1(c_82_1500) );
  Fadder_ A_83_1526( .carry(c_83_1526), .sum(s_83_1526), .in3(c_82_1499), .in2(s_83_1521), .in1(s_83_1522) );
  Fadder_ A_83_1527( .carry(c_83_1527), .sum(s_83_1527), .in3(s_83_1523), .in2(c_82_1501), .in1(c_82_1502) );
  Fadder_ A_83_1528( .carry(c_83_1528), .sum(s_83_1528), .in3(s_83_1524), .in2(c_82_1503), .in1(c_82_1504) );
  Fadder_ A_83_1529( .carry(c_83_1529), .sum(s_83_1529), .in3(s_83_1525), .in2(s_83_1526), .in1(c_82_1505) );
  Fadder_ A_83_1530( .carry(c_83_1530), .sum(s_83_1530), .in3(s_83_1527), .in2(c_82_1506), .in1(s_83_1528) );
  Fadder_ A_83_1531( .carry(c_83_1531), .sum(s_83_1531), .in3(c_82_1507), .in2(s_83_1529), .in1(c_82_1508) );
  Fadder_ A_83_1532( .carry(c[83]), .sum(s[83]), .in3(s_83_1530), .in2(c_82_1509), .in1(s_83_1531) );

  // ***** Bit 84 ***** //
  Hadder_ A_84_1533( .carry(c_84_1533), .sum(s_84_1533), .in2(sign_), .in1(P_31[22]) );
  Fadder_ A_84_1534( .carry(c_84_1534), .sum(s_84_1534), .in3(P_30[24]), .in2(P_29[26]), .in1(P_28[28]) );
  Fadder_ A_84_1535( .carry(c_84_1535), .sum(s_84_1535), .in3(P_27[30]), .in2(P_26[32]), .in1(P_25[34]) );
  Fadder_ A_84_1536( .carry(c_84_1536), .sum(s_84_1536), .in3(P_24[36]), .in2(P_23[38]), .in1(P_22[40]) );
  Fadder_ A_84_1537( .carry(c_84_1537), .sum(s_84_1537), .in3(P_21[42]), .in2(P_20[44]), .in1(P_19[46]) );
  Fadder_ A_84_1538( .carry(c_84_1538), .sum(s_84_1538), .in3(P_18[48]), .in2(P_17[50]), .in1(P_16[52]) );
  Fadder_ A_84_1539( .carry(c_84_1539), .sum(s_84_1539), .in3(P_15[54]), .in2(P_14[56]), .in1(P_13[58]) );
  Fadder_ A_84_1540( .carry(c_84_1540), .sum(s_84_1540), .in3(P_12[60]), .in2(P_11[62]), .in1(P_10[64]) );
  Fadder_ A_84_1541( .carry(c_84_1541), .sum(s_84_1541), .in3(c_83_1517), .in2(c_83_1516), .in1(c_83_1515) );
  Fadder_ A_84_1542( .carry(c_84_1542), .sum(s_84_1542), .in3(c_83_1514), .in2(c_83_1513), .in1(c_83_1512) );
  Fadder_ A_84_1543( .carry(c_84_1543), .sum(s_84_1543), .in3(c_83_1511), .in2(s_84_1533), .in1(s_84_1540) );
  Fadder_ A_84_1544( .carry(c_84_1544), .sum(s_84_1544), .in3(s_84_1539), .in2(s_84_1538), .in1(s_84_1537) );
  Fadder_ A_84_1545( .carry(c_84_1545), .sum(s_84_1545), .in3(s_84_1536), .in2(s_84_1535), .in1(s_84_1534) );
  Fadder_ A_84_1546( .carry(c_84_1546), .sum(s_84_1546), .in3(c_83_1518), .in2(c_83_1520), .in1(c_83_1519) );
  Fadder_ A_84_1547( .carry(c_84_1547), .sum(s_84_1547), .in3(s_84_1542), .in2(s_84_1541), .in1(c_83_1522) );
  Fadder_ A_84_1548( .carry(c_84_1548), .sum(s_84_1548), .in3(c_83_1521), .in2(s_84_1543), .in1(s_84_1545) );
  Fadder_ A_84_1549( .carry(c_84_1549), .sum(s_84_1549), .in3(s_84_1544), .in2(c_83_1523), .in1(c_83_1524) );
  Fadder_ A_84_1550( .carry(c_84_1550), .sum(s_84_1550), .in3(s_84_1546), .in2(c_83_1525), .in1(c_83_1526) );
  Fadder_ A_84_1551( .carry(c_84_1551), .sum(s_84_1551), .in3(s_84_1547), .in2(s_84_1548), .in1(c_83_1527) );
  Fadder_ A_84_1552( .carry(c_84_1552), .sum(s_84_1552), .in3(s_84_1549), .in2(c_83_1528), .in1(s_84_1550) );
  Fadder_ A_84_1553( .carry(c_84_1553), .sum(s_84_1553), .in3(c_83_1529), .in2(s_84_1551), .in1(c_83_1530) );
  Fadder_ A_84_1554( .carry(c[84]), .sum(s[84]), .in3(s_84_1552), .in2(c_83_1531), .in1(s_84_1553) );

  // ***** Bit 85 ***** //
  Fadder_ A_85_1555( .carry(c_85_1555), .sum(s_85_1555), .in3(P_31[23]), .in2(P_30[25]), .in1(P_29[27]) );
  Fadder_ A_85_1556( .carry(c_85_1556), .sum(s_85_1556), .in3(P_28[29]), .in2(P_27[31]), .in1(P_26[33]) );
  Fadder_ A_85_1557( .carry(c_85_1557), .sum(s_85_1557), .in3(P_25[35]), .in2(P_24[37]), .in1(P_23[39]) );
  Fadder_ A_85_1558( .carry(c_85_1558), .sum(s_85_1558), .in3(P_22[41]), .in2(P_21[43]), .in1(P_20[45]) );
  Fadder_ A_85_1559( .carry(c_85_1559), .sum(s_85_1559), .in3(P_19[47]), .in2(P_18[49]), .in1(P_17[51]) );
  Fadder_ A_85_1560( .carry(c_85_1560), .sum(s_85_1560), .in3(P_16[53]), .in2(P_15[55]), .in1(P_14[57]) );
  Fadder_ A_85_1561( .carry(c_85_1561), .sum(s_85_1561), .in3(P_13[59]), .in2(P_12[61]), .in1(P_11[63]) );
  Fadder_ A_85_1562( .carry(c_85_1562), .sum(s_85_1562), .in3(P_10[65]), .in2(c_84_1533), .in1(c_84_1540) );
  Fadder_ A_85_1563( .carry(c_85_1563), .sum(s_85_1563), .in3(c_84_1539), .in2(c_84_1538), .in1(c_84_1537) );
  Fadder_ A_85_1564( .carry(c_85_1564), .sum(s_85_1564), .in3(c_84_1536), .in2(c_84_1535), .in1(c_84_1534) );
  Fadder_ A_85_1565( .carry(c_85_1565), .sum(s_85_1565), .in3(s_85_1561), .in2(s_85_1560), .in1(s_85_1559) );
  Fadder_ A_85_1566( .carry(c_85_1566), .sum(s_85_1566), .in3(s_85_1558), .in2(s_85_1557), .in1(s_85_1556) );
  Fadder_ A_85_1567( .carry(c_85_1567), .sum(s_85_1567), .in3(s_85_1555), .in2(c_84_1542), .in1(c_84_1541) );
  Fadder_ A_85_1568( .carry(c_85_1568), .sum(s_85_1568), .in3(c_84_1543), .in2(s_85_1562), .in1(s_85_1564) );
  Fadder_ A_85_1569( .carry(c_85_1569), .sum(s_85_1569), .in3(s_85_1563), .in2(c_84_1545), .in1(c_84_1544) );
  Fadder_ A_85_1570( .carry(c_85_1570), .sum(s_85_1570), .in3(s_85_1566), .in2(s_85_1565), .in1(c_84_1546) );
  Fadder_ A_85_1571( .carry(c_85_1571), .sum(s_85_1571), .in3(s_85_1567), .in2(c_84_1547), .in1(s_85_1568) );
  Fadder_ A_85_1572( .carry(c_85_1572), .sum(s_85_1572), .in3(c_84_1548), .in2(s_85_1569), .in1(c_84_1549) );
  Fadder_ A_85_1573( .carry(c_85_1573), .sum(s_85_1573), .in3(s_85_1570), .in2(c_84_1550), .in1(s_85_1571) );
  Fadder_ A_85_1574( .carry(c_85_1574), .sum(s_85_1574), .in3(c_84_1551), .in2(s_85_1572), .in1(c_84_1552) );
  Fadder_ A_85_1575( .carry(c[85]), .sum(s[85]), .in3(s_85_1573), .in2(c_84_1553), .in1(s_85_1574) );

  // ***** Bit 86 ***** //
  Hadder_ A_86_1576( .carry(c_86_1576), .sum(s_86_1576), .in2(sign_), .in1(P_31[24]) );
  Fadder_ A_86_1577( .carry(c_86_1577), .sum(s_86_1577), .in3(P_30[26]), .in2(P_29[28]), .in1(P_28[30]) );
  Fadder_ A_86_1578( .carry(c_86_1578), .sum(s_86_1578), .in3(P_27[32]), .in2(P_26[34]), .in1(P_25[36]) );
  Fadder_ A_86_1579( .carry(c_86_1579), .sum(s_86_1579), .in3(P_24[38]), .in2(P_23[40]), .in1(P_22[42]) );
  Fadder_ A_86_1580( .carry(c_86_1580), .sum(s_86_1580), .in3(P_21[44]), .in2(P_20[46]), .in1(P_19[48]) );
  Fadder_ A_86_1581( .carry(c_86_1581), .sum(s_86_1581), .in3(P_18[50]), .in2(P_17[52]), .in1(P_16[54]) );
  Fadder_ A_86_1582( .carry(c_86_1582), .sum(s_86_1582), .in3(P_15[56]), .in2(P_14[58]), .in1(P_13[60]) );
  Fadder_ A_86_1583( .carry(c_86_1583), .sum(s_86_1583), .in3(P_12[62]), .in2(P_11[64]), .in1(c_85_1561) );
  Fadder_ A_86_1584( .carry(c_86_1584), .sum(s_86_1584), .in3(c_85_1560), .in2(c_85_1559), .in1(c_85_1558) );
  Fadder_ A_86_1585( .carry(c_86_1585), .sum(s_86_1585), .in3(c_85_1557), .in2(c_85_1556), .in1(c_85_1555) );
  Fadder_ A_86_1586( .carry(c_86_1586), .sum(s_86_1586), .in3(s_86_1576), .in2(s_86_1582), .in1(s_86_1581) );
  Fadder_ A_86_1587( .carry(c_86_1587), .sum(s_86_1587), .in3(s_86_1580), .in2(s_86_1579), .in1(s_86_1578) );
  Fadder_ A_86_1588( .carry(c_86_1588), .sum(s_86_1588), .in3(s_86_1577), .in2(c_85_1562), .in1(c_85_1564) );
  Fadder_ A_86_1589( .carry(c_86_1589), .sum(s_86_1589), .in3(c_85_1563), .in2(s_86_1583), .in1(s_86_1585) );
  Fadder_ A_86_1590( .carry(c_86_1590), .sum(s_86_1590), .in3(s_86_1584), .in2(c_85_1566), .in1(c_85_1565) );
  Fadder_ A_86_1591( .carry(c_86_1591), .sum(s_86_1591), .in3(s_86_1586), .in2(s_86_1587), .in1(c_85_1567) );
  Fadder_ A_86_1592( .carry(c_86_1592), .sum(s_86_1592), .in3(s_86_1588), .in2(c_85_1568), .in1(c_85_1569) );
  Fadder_ A_86_1593( .carry(c_86_1593), .sum(s_86_1593), .in3(s_86_1589), .in2(s_86_1590), .in1(c_85_1570) );
  Fadder_ A_86_1594( .carry(c_86_1594), .sum(s_86_1594), .in3(s_86_1591), .in2(c_85_1571), .in1(s_86_1592) );
  Fadder_ A_86_1595( .carry(c_86_1595), .sum(s_86_1595), .in3(c_85_1572), .in2(s_86_1593), .in1(c_85_1573) );
  Fadder_ A_86_1596( .carry(c[86]), .sum(s[86]), .in3(s_86_1594), .in2(c_85_1574), .in1(s_86_1595) );

  // ***** Bit 87 ***** //
  Fadder_ A_87_1597( .carry(c_87_1597), .sum(s_87_1597), .in3(P_31[25]), .in2(P_30[27]), .in1(P_29[29]) );
  Fadder_ A_87_1598( .carry(c_87_1598), .sum(s_87_1598), .in3(P_28[31]), .in2(P_27[33]), .in1(P_26[35]) );
  Fadder_ A_87_1599( .carry(c_87_1599), .sum(s_87_1599), .in3(P_25[37]), .in2(P_24[39]), .in1(P_23[41]) );
  Fadder_ A_87_1600( .carry(c_87_1600), .sum(s_87_1600), .in3(P_22[43]), .in2(P_21[45]), .in1(P_20[47]) );
  Fadder_ A_87_1601( .carry(c_87_1601), .sum(s_87_1601), .in3(P_19[49]), .in2(P_18[51]), .in1(P_17[53]) );
  Fadder_ A_87_1602( .carry(c_87_1602), .sum(s_87_1602), .in3(P_16[55]), .in2(P_15[57]), .in1(P_14[59]) );
  Fadder_ A_87_1603( .carry(c_87_1603), .sum(s_87_1603), .in3(P_13[61]), .in2(P_12[63]), .in1(P_11[65]) );
  Fadder_ A_87_1604( .carry(c_87_1604), .sum(s_87_1604), .in3(c_86_1576), .in2(c_86_1582), .in1(c_86_1581) );
  Fadder_ A_87_1605( .carry(c_87_1605), .sum(s_87_1605), .in3(c_86_1580), .in2(c_86_1579), .in1(c_86_1578) );
  Fadder_ A_87_1606( .carry(c_87_1606), .sum(s_87_1606), .in3(c_86_1577), .in2(s_87_1603), .in1(s_87_1602) );
  Fadder_ A_87_1607( .carry(c_87_1607), .sum(s_87_1607), .in3(s_87_1601), .in2(s_87_1600), .in1(s_87_1599) );
  Fadder_ A_87_1608( .carry(c_87_1608), .sum(s_87_1608), .in3(s_87_1598), .in2(s_87_1597), .in1(c_86_1583) );
  Fadder_ A_87_1609( .carry(c_87_1609), .sum(s_87_1609), .in3(c_86_1585), .in2(c_86_1584), .in1(s_87_1604) );
  Fadder_ A_87_1610( .carry(c_87_1610), .sum(s_87_1610), .in3(s_87_1605), .in2(c_86_1587), .in1(c_86_1586) );
  Fadder_ A_87_1611( .carry(c_87_1611), .sum(s_87_1611), .in3(s_87_1606), .in2(s_87_1607), .in1(c_86_1588) );
  Fadder_ A_87_1612( .carry(c_87_1612), .sum(s_87_1612), .in3(s_87_1608), .in2(c_86_1589), .in1(c_86_1590) );
  Fadder_ A_87_1613( .carry(c_87_1613), .sum(s_87_1613), .in3(s_87_1609), .in2(s_87_1610), .in1(c_86_1591) );
  Fadder_ A_87_1614( .carry(c_87_1614), .sum(s_87_1614), .in3(s_87_1611), .in2(c_86_1592), .in1(s_87_1612) );
  Fadder_ A_87_1615( .carry(c_87_1615), .sum(s_87_1615), .in3(c_86_1593), .in2(s_87_1613), .in1(c_86_1594) );
  Fadder_ A_87_1616( .carry(c[87]), .sum(s[87]), .in3(s_87_1614), .in2(c_86_1595), .in1(s_87_1615) );

  // ***** Bit 88 ***** //
  Hadder_ A_88_1617( .carry(c_88_1617), .sum(s_88_1617), .in2(sign_), .in1(P_31[26]) );
  Fadder_ A_88_1618( .carry(c_88_1618), .sum(s_88_1618), .in3(P_30[28]), .in2(P_29[30]), .in1(P_28[32]) );
  Fadder_ A_88_1619( .carry(c_88_1619), .sum(s_88_1619), .in3(P_27[34]), .in2(P_26[36]), .in1(P_25[38]) );
  Fadder_ A_88_1620( .carry(c_88_1620), .sum(s_88_1620), .in3(P_24[40]), .in2(P_23[42]), .in1(P_22[44]) );
  Fadder_ A_88_1621( .carry(c_88_1621), .sum(s_88_1621), .in3(P_21[46]), .in2(P_20[48]), .in1(P_19[50]) );
  Fadder_ A_88_1622( .carry(c_88_1622), .sum(s_88_1622), .in3(P_18[52]), .in2(P_17[54]), .in1(P_16[56]) );
  Fadder_ A_88_1623( .carry(c_88_1623), .sum(s_88_1623), .in3(P_15[58]), .in2(P_14[60]), .in1(P_13[62]) );
  Fadder_ A_88_1624( .carry(c_88_1624), .sum(s_88_1624), .in3(P_12[64]), .in2(c_87_1603), .in1(c_87_1602) );
  Fadder_ A_88_1625( .carry(c_88_1625), .sum(s_88_1625), .in3(c_87_1601), .in2(c_87_1600), .in1(c_87_1599) );
  Fadder_ A_88_1626( .carry(c_88_1626), .sum(s_88_1626), .in3(c_87_1598), .in2(c_87_1597), .in1(s_88_1617) );
  Fadder_ A_88_1627( .carry(c_88_1627), .sum(s_88_1627), .in3(s_88_1623), .in2(s_88_1622), .in1(s_88_1621) );
  Fadder_ A_88_1628( .carry(c_88_1628), .sum(s_88_1628), .in3(s_88_1620), .in2(s_88_1619), .in1(s_88_1618) );
  Fadder_ A_88_1629( .carry(c_88_1629), .sum(s_88_1629), .in3(c_87_1605), .in2(c_87_1604), .in1(s_88_1624) );
  Fadder_ A_88_1630( .carry(c_88_1630), .sum(s_88_1630), .in3(s_88_1625), .in2(c_87_1607), .in1(c_87_1606) );
  Fadder_ A_88_1631( .carry(c_88_1631), .sum(s_88_1631), .in3(s_88_1626), .in2(s_88_1628), .in1(s_88_1627) );
  Fadder_ A_88_1632( .carry(c_88_1632), .sum(s_88_1632), .in3(c_87_1608), .in2(c_87_1609), .in1(c_87_1610) );
  Fadder_ A_88_1633( .carry(c_88_1633), .sum(s_88_1633), .in3(s_88_1629), .in2(s_88_1630), .in1(s_88_1631) );
  Fadder_ A_88_1634( .carry(c_88_1634), .sum(s_88_1634), .in3(c_87_1611), .in2(c_87_1612), .in1(s_88_1632) );
  Fadder_ A_88_1635( .carry(c_88_1635), .sum(s_88_1635), .in3(c_87_1613), .in2(s_88_1633), .in1(c_87_1614) );
  Fadder_ A_88_1636( .carry(c[88]), .sum(s[88]), .in3(s_88_1634), .in2(c_87_1615), .in1(s_88_1635) );

  // ***** Bit 89 ***** //
  Fadder_ A_89_1637( .carry(c_89_1637), .sum(s_89_1637), .in3(P_31[27]), .in2(P_30[29]), .in1(P_29[31]) );
  Fadder_ A_89_1638( .carry(c_89_1638), .sum(s_89_1638), .in3(P_28[33]), .in2(P_27[35]), .in1(P_26[37]) );
  Fadder_ A_89_1639( .carry(c_89_1639), .sum(s_89_1639), .in3(P_25[39]), .in2(P_24[41]), .in1(P_23[43]) );
  Fadder_ A_89_1640( .carry(c_89_1640), .sum(s_89_1640), .in3(P_22[45]), .in2(P_21[47]), .in1(P_20[49]) );
  Fadder_ A_89_1641( .carry(c_89_1641), .sum(s_89_1641), .in3(P_19[51]), .in2(P_18[53]), .in1(P_17[55]) );
  Fadder_ A_89_1642( .carry(c_89_1642), .sum(s_89_1642), .in3(P_16[57]), .in2(P_15[59]), .in1(P_14[61]) );
  Fadder_ A_89_1643( .carry(c_89_1643), .sum(s_89_1643), .in3(P_13[63]), .in2(P_12[65]), .in1(c_88_1617) );
  Fadder_ A_89_1644( .carry(c_89_1644), .sum(s_89_1644), .in3(c_88_1623), .in2(c_88_1622), .in1(c_88_1621) );
  Fadder_ A_89_1645( .carry(c_89_1645), .sum(s_89_1645), .in3(c_88_1620), .in2(c_88_1619), .in1(c_88_1618) );
  Fadder_ A_89_1646( .carry(c_89_1646), .sum(s_89_1646), .in3(s_89_1642), .in2(s_89_1641), .in1(s_89_1640) );
  Fadder_ A_89_1647( .carry(c_89_1647), .sum(s_89_1647), .in3(s_89_1639), .in2(s_89_1638), .in1(s_89_1637) );
  Fadder_ A_89_1648( .carry(c_89_1648), .sum(s_89_1648), .in3(s_89_1643), .in2(c_88_1626), .in1(c_88_1625) );
  Fadder_ A_89_1649( .carry(c_89_1649), .sum(s_89_1649), .in3(c_88_1624), .in2(s_89_1645), .in1(s_89_1644) );
  Fadder_ A_89_1650( .carry(c_89_1650), .sum(s_89_1650), .in3(c_88_1628), .in2(c_88_1627), .in1(s_89_1647) );
  Fadder_ A_89_1651( .carry(c_89_1651), .sum(s_89_1651), .in3(s_89_1646), .in2(c_88_1629), .in1(s_89_1648) );
  Fadder_ A_89_1652( .carry(c_89_1652), .sum(s_89_1652), .in3(c_88_1630), .in2(s_89_1649), .in1(c_88_1631) );
  Fadder_ A_89_1653( .carry(c_89_1653), .sum(s_89_1653), .in3(s_89_1650), .in2(c_88_1632), .in1(s_89_1651) );
  Fadder_ A_89_1654( .carry(c_89_1654), .sum(s_89_1654), .in3(c_88_1633), .in2(s_89_1652), .in1(c_88_1634) );
  Fadder_ A_89_1655( .carry(c[89]), .sum(s[89]), .in3(s_89_1653), .in2(c_88_1635), .in1(s_89_1654) );

  // ***** Bit 90 ***** //
  Hadder_ A_90_1656( .carry(c_90_1656), .sum(s_90_1656), .in2(sign_), .in1(P_31[28]) );
  Fadder_ A_90_1657( .carry(c_90_1657), .sum(s_90_1657), .in3(P_30[30]), .in2(P_29[32]), .in1(P_28[34]) );
  Fadder_ A_90_1658( .carry(c_90_1658), .sum(s_90_1658), .in3(P_27[36]), .in2(P_26[38]), .in1(P_25[40]) );
  Fadder_ A_90_1659( .carry(c_90_1659), .sum(s_90_1659), .in3(P_24[42]), .in2(P_23[44]), .in1(P_22[46]) );
  Fadder_ A_90_1660( .carry(c_90_1660), .sum(s_90_1660), .in3(P_21[48]), .in2(P_20[50]), .in1(P_19[52]) );
  Fadder_ A_90_1661( .carry(c_90_1661), .sum(s_90_1661), .in3(P_18[54]), .in2(P_17[56]), .in1(P_16[58]) );
  Fadder_ A_90_1662( .carry(c_90_1662), .sum(s_90_1662), .in3(P_15[60]), .in2(P_14[62]), .in1(P_13[64]) );
  Fadder_ A_90_1663( .carry(c_90_1663), .sum(s_90_1663), .in3(c_89_1642), .in2(c_89_1641), .in1(c_89_1640) );
  Fadder_ A_90_1664( .carry(c_90_1664), .sum(s_90_1664), .in3(c_89_1639), .in2(c_89_1638), .in1(c_89_1637) );
  Fadder_ A_90_1665( .carry(c_90_1665), .sum(s_90_1665), .in3(s_90_1656), .in2(s_90_1662), .in1(s_90_1661) );
  Fadder_ A_90_1666( .carry(c_90_1666), .sum(s_90_1666), .in3(s_90_1660), .in2(s_90_1659), .in1(s_90_1658) );
  Fadder_ A_90_1667( .carry(c_90_1667), .sum(s_90_1667), .in3(s_90_1657), .in2(c_89_1643), .in1(c_89_1645) );
  Fadder_ A_90_1668( .carry(c_90_1668), .sum(s_90_1668), .in3(c_89_1644), .in2(s_90_1664), .in1(s_90_1663) );
  Fadder_ A_90_1669( .carry(c_90_1669), .sum(s_90_1669), .in3(c_89_1647), .in2(c_89_1646), .in1(s_90_1665) );
  Fadder_ A_90_1670( .carry(c_90_1670), .sum(s_90_1670), .in3(s_90_1666), .in2(c_89_1648), .in1(s_90_1667) );
  Fadder_ A_90_1671( .carry(c_90_1671), .sum(s_90_1671), .in3(c_89_1649), .in2(c_89_1650), .in1(s_90_1668) );
  Fadder_ A_90_1672( .carry(c_90_1672), .sum(s_90_1672), .in3(s_90_1669), .in2(c_89_1651), .in1(s_90_1670) );
  Fadder_ A_90_1673( .carry(c_90_1673), .sum(s_90_1673), .in3(c_89_1652), .in2(s_90_1671), .in1(c_89_1653) );
  Fadder_ A_90_1674( .carry(c[90]), .sum(s[90]), .in3(s_90_1672), .in2(c_89_1654), .in1(s_90_1673) );

  // ***** Bit 91 ***** //
  Fadder_ A_91_1675( .carry(c_91_1675), .sum(s_91_1675), .in3(P_31[29]), .in2(P_30[31]), .in1(P_29[33]) );
  Fadder_ A_91_1676( .carry(c_91_1676), .sum(s_91_1676), .in3(P_28[35]), .in2(P_27[37]), .in1(P_26[39]) );
  Fadder_ A_91_1677( .carry(c_91_1677), .sum(s_91_1677), .in3(P_25[41]), .in2(P_24[43]), .in1(P_23[45]) );
  Fadder_ A_91_1678( .carry(c_91_1678), .sum(s_91_1678), .in3(P_22[47]), .in2(P_21[49]), .in1(P_20[51]) );
  Fadder_ A_91_1679( .carry(c_91_1679), .sum(s_91_1679), .in3(P_19[53]), .in2(P_18[55]), .in1(P_17[57]) );
  Fadder_ A_91_1680( .carry(c_91_1680), .sum(s_91_1680), .in3(P_16[59]), .in2(P_15[61]), .in1(P_14[63]) );
  Fadder_ A_91_1681( .carry(c_91_1681), .sum(s_91_1681), .in3(P_13[65]), .in2(c_90_1656), .in1(c_90_1662) );
  Fadder_ A_91_1682( .carry(c_91_1682), .sum(s_91_1682), .in3(c_90_1661), .in2(c_90_1660), .in1(c_90_1659) );
  Fadder_ A_91_1683( .carry(c_91_1683), .sum(s_91_1683), .in3(c_90_1658), .in2(c_90_1657), .in1(s_91_1680) );
  Fadder_ A_91_1684( .carry(c_91_1684), .sum(s_91_1684), .in3(s_91_1679), .in2(s_91_1678), .in1(s_91_1677) );
  Fadder_ A_91_1685( .carry(c_91_1685), .sum(s_91_1685), .in3(s_91_1676), .in2(s_91_1675), .in1(c_90_1664) );
  Fadder_ A_91_1686( .carry(c_91_1686), .sum(s_91_1686), .in3(c_90_1663), .in2(s_91_1681), .in1(s_91_1682) );
  Fadder_ A_91_1687( .carry(c_91_1687), .sum(s_91_1687), .in3(c_90_1666), .in2(c_90_1665), .in1(s_91_1683) );
  Fadder_ A_91_1688( .carry(c_91_1688), .sum(s_91_1688), .in3(s_91_1684), .in2(c_90_1667), .in1(s_91_1685) );
  Fadder_ A_91_1689( .carry(c_91_1689), .sum(s_91_1689), .in3(c_90_1668), .in2(c_90_1669), .in1(s_91_1686) );
  Fadder_ A_91_1690( .carry(c_91_1690), .sum(s_91_1690), .in3(s_91_1687), .in2(c_90_1670), .in1(c_90_1671) );
  Fadder_ A_91_1691( .carry(c_91_1691), .sum(s_91_1691), .in3(s_91_1688), .in2(s_91_1689), .in1(c_90_1672) );
  Fadder_ A_91_1692( .carry(c[91]), .sum(s[91]), .in3(s_91_1690), .in2(c_90_1673), .in1(s_91_1691) );

  // ***** Bit 92 ***** //
  Hadder_ A_92_1693( .carry(c_92_1693), .sum(s_92_1693), .in2(sign_), .in1(P_31[30]) );
  Fadder_ A_92_1694( .carry(c_92_1694), .sum(s_92_1694), .in3(P_30[32]), .in2(P_29[34]), .in1(P_28[36]) );
  Fadder_ A_92_1695( .carry(c_92_1695), .sum(s_92_1695), .in3(P_27[38]), .in2(P_26[40]), .in1(P_25[42]) );
  Fadder_ A_92_1696( .carry(c_92_1696), .sum(s_92_1696), .in3(P_24[44]), .in2(P_23[46]), .in1(P_22[48]) );
  Fadder_ A_92_1697( .carry(c_92_1697), .sum(s_92_1697), .in3(P_21[50]), .in2(P_20[52]), .in1(P_19[54]) );
  Fadder_ A_92_1698( .carry(c_92_1698), .sum(s_92_1698), .in3(P_18[56]), .in2(P_17[58]), .in1(P_16[60]) );
  Fadder_ A_92_1699( .carry(c_92_1699), .sum(s_92_1699), .in3(P_15[62]), .in2(P_14[64]), .in1(c_91_1680) );
  Fadder_ A_92_1700( .carry(c_92_1700), .sum(s_92_1700), .in3(c_91_1679), .in2(c_91_1678), .in1(c_91_1677) );
  Fadder_ A_92_1701( .carry(c_92_1701), .sum(s_92_1701), .in3(c_91_1676), .in2(c_91_1675), .in1(s_92_1693) );
  Fadder_ A_92_1702( .carry(c_92_1702), .sum(s_92_1702), .in3(s_92_1698), .in2(s_92_1697), .in1(s_92_1696) );
  Fadder_ A_92_1703( .carry(c_92_1703), .sum(s_92_1703), .in3(s_92_1695), .in2(s_92_1694), .in1(c_91_1681) );
  Fadder_ A_92_1704( .carry(c_92_1704), .sum(s_92_1704), .in3(c_91_1682), .in2(c_91_1683), .in1(s_92_1699) );
  Fadder_ A_92_1705( .carry(c_92_1705), .sum(s_92_1705), .in3(s_92_1700), .in2(c_91_1684), .in1(s_92_1701) );
  Fadder_ A_92_1706( .carry(c_92_1706), .sum(s_92_1706), .in3(s_92_1702), .in2(c_91_1685), .in1(s_92_1703) );
  Fadder_ A_92_1707( .carry(c_92_1707), .sum(s_92_1707), .in3(c_91_1686), .in2(c_91_1687), .in1(s_92_1704) );
  Fadder_ A_92_1708( .carry(c_92_1708), .sum(s_92_1708), .in3(s_92_1705), .in2(c_91_1688), .in1(s_92_1706) );
  Fadder_ A_92_1709( .carry(c_92_1709), .sum(s_92_1709), .in3(c_91_1689), .in2(s_92_1707), .in1(c_91_1690) );
  Fadder_ A_92_1710( .carry(c[92]), .sum(s[92]), .in3(s_92_1708), .in2(c_91_1691), .in1(s_92_1709) );

  // ***** Bit 93 ***** //
  Fadder_ A_93_1711( .carry(c_93_1711), .sum(s_93_1711), .in3(P_31[31]), .in2(P_30[33]), .in1(P_29[35]) );
  Fadder_ A_93_1712( .carry(c_93_1712), .sum(s_93_1712), .in3(P_28[37]), .in2(P_27[39]), .in1(P_26[41]) );
  Fadder_ A_93_1713( .carry(c_93_1713), .sum(s_93_1713), .in3(P_25[43]), .in2(P_24[45]), .in1(P_23[47]) );
  Fadder_ A_93_1714( .carry(c_93_1714), .sum(s_93_1714), .in3(P_22[49]), .in2(P_21[51]), .in1(P_20[53]) );
  Fadder_ A_93_1715( .carry(c_93_1715), .sum(s_93_1715), .in3(P_19[55]), .in2(P_18[57]), .in1(P_17[59]) );
  Fadder_ A_93_1716( .carry(c_93_1716), .sum(s_93_1716), .in3(P_16[61]), .in2(P_15[63]), .in1(P_14[65]) );
  Fadder_ A_93_1717( .carry(c_93_1717), .sum(s_93_1717), .in3(c_92_1693), .in2(c_92_1698), .in1(c_92_1697) );
  Fadder_ A_93_1718( .carry(c_93_1718), .sum(s_93_1718), .in3(c_92_1696), .in2(c_92_1695), .in1(c_92_1694) );
  Fadder_ A_93_1719( .carry(c_93_1719), .sum(s_93_1719), .in3(s_93_1716), .in2(s_93_1715), .in1(s_93_1714) );
  Fadder_ A_93_1720( .carry(c_93_1720), .sum(s_93_1720), .in3(s_93_1713), .in2(s_93_1712), .in1(s_93_1711) );
  Fadder_ A_93_1721( .carry(c_93_1721), .sum(s_93_1721), .in3(c_92_1699), .in2(c_92_1701), .in1(c_92_1700) );
  Fadder_ A_93_1722( .carry(c_93_1722), .sum(s_93_1722), .in3(s_93_1717), .in2(s_93_1718), .in1(c_92_1702) );
  Fadder_ A_93_1723( .carry(c_93_1723), .sum(s_93_1723), .in3(s_93_1720), .in2(s_93_1719), .in1(c_92_1703) );
  Fadder_ A_93_1724( .carry(c_93_1724), .sum(s_93_1724), .in3(c_92_1704), .in2(s_93_1721), .in1(c_92_1705) );
  Fadder_ A_93_1725( .carry(c_93_1725), .sum(s_93_1725), .in3(s_93_1722), .in2(s_93_1723), .in1(c_92_1706) );
  Fadder_ A_93_1726( .carry(c_93_1726), .sum(s_93_1726), .in3(c_92_1707), .in2(s_93_1724), .in1(s_93_1725) );
  Fadder_ A_93_1727( .carry(c[93]), .sum(s[93]), .in3(c_92_1708), .in2(c_92_1709), .in1(s_93_1726) );

  // ***** Bit 94 ***** //
  Hadder_ A_94_1728( .carry(c_94_1728), .sum(s_94_1728), .in2(sign_), .in1(P_31[32]) );
  Fadder_ A_94_1729( .carry(c_94_1729), .sum(s_94_1729), .in3(P_30[34]), .in2(P_29[36]), .in1(P_28[38]) );
  Fadder_ A_94_1730( .carry(c_94_1730), .sum(s_94_1730), .in3(P_27[40]), .in2(P_26[42]), .in1(P_25[44]) );
  Fadder_ A_94_1731( .carry(c_94_1731), .sum(s_94_1731), .in3(P_24[46]), .in2(P_23[48]), .in1(P_22[50]) );
  Fadder_ A_94_1732( .carry(c_94_1732), .sum(s_94_1732), .in3(P_21[52]), .in2(P_20[54]), .in1(P_19[56]) );
  Fadder_ A_94_1733( .carry(c_94_1733), .sum(s_94_1733), .in3(P_18[58]), .in2(P_17[60]), .in1(P_16[62]) );
  Fadder_ A_94_1734( .carry(c_94_1734), .sum(s_94_1734), .in3(P_15[64]), .in2(c_93_1716), .in1(c_93_1715) );
  Fadder_ A_94_1735( .carry(c_94_1735), .sum(s_94_1735), .in3(c_93_1714), .in2(c_93_1713), .in1(c_93_1712) );
  Fadder_ A_94_1736( .carry(c_94_1736), .sum(s_94_1736), .in3(c_93_1711), .in2(s_94_1728), .in1(s_94_1733) );
  Fadder_ A_94_1737( .carry(c_94_1737), .sum(s_94_1737), .in3(s_94_1732), .in2(s_94_1731), .in1(s_94_1730) );
  Fadder_ A_94_1738( .carry(c_94_1738), .sum(s_94_1738), .in3(s_94_1729), .in2(c_93_1718), .in1(c_93_1717) );
  Fadder_ A_94_1739( .carry(c_94_1739), .sum(s_94_1739), .in3(s_94_1734), .in2(s_94_1735), .in1(c_93_1720) );
  Fadder_ A_94_1740( .carry(c_94_1740), .sum(s_94_1740), .in3(c_93_1719), .in2(s_94_1736), .in1(s_94_1737) );
  Fadder_ A_94_1741( .carry(c_94_1741), .sum(s_94_1741), .in3(c_93_1721), .in2(s_94_1738), .in1(c_93_1722) );
  Fadder_ A_94_1742( .carry(c_94_1742), .sum(s_94_1742), .in3(s_94_1739), .in2(c_93_1723), .in1(s_94_1740) );
  Fadder_ A_94_1743( .carry(c_94_1743), .sum(s_94_1743), .in3(c_93_1724), .in2(s_94_1741), .in1(s_94_1742) );
  Fadder_ A_94_1744( .carry(c[94]), .sum(s[94]), .in3(c_93_1725), .in2(c_93_1726), .in1(s_94_1743) );

  // ***** Bit 95 ***** //
  Fadder_ A_95_1745( .carry(c_95_1745), .sum(s_95_1745), .in3(P_31[33]), .in2(P_30[35]), .in1(P_29[37]) );
  Fadder_ A_95_1746( .carry(c_95_1746), .sum(s_95_1746), .in3(P_28[39]), .in2(P_27[41]), .in1(P_26[43]) );
  Fadder_ A_95_1747( .carry(c_95_1747), .sum(s_95_1747), .in3(P_25[45]), .in2(P_24[47]), .in1(P_23[49]) );
  Fadder_ A_95_1748( .carry(c_95_1748), .sum(s_95_1748), .in3(P_22[51]), .in2(P_21[53]), .in1(P_20[55]) );
  Fadder_ A_95_1749( .carry(c_95_1749), .sum(s_95_1749), .in3(P_19[57]), .in2(P_18[59]), .in1(P_17[61]) );
  Fadder_ A_95_1750( .carry(c_95_1750), .sum(s_95_1750), .in3(P_16[63]), .in2(P_15[65]), .in1(c_94_1728) );
  Fadder_ A_95_1751( .carry(c_95_1751), .sum(s_95_1751), .in3(c_94_1733), .in2(c_94_1732), .in1(c_94_1731) );
  Fadder_ A_95_1752( .carry(c_95_1752), .sum(s_95_1752), .in3(c_94_1730), .in2(c_94_1729), .in1(s_95_1749) );
  Fadder_ A_95_1753( .carry(c_95_1753), .sum(s_95_1753), .in3(s_95_1748), .in2(s_95_1747), .in1(s_95_1746) );
  Fadder_ A_95_1754( .carry(c_95_1754), .sum(s_95_1754), .in3(s_95_1745), .in2(s_95_1750), .in1(c_94_1735) );
  Fadder_ A_95_1755( .carry(c_95_1755), .sum(s_95_1755), .in3(c_94_1734), .in2(c_94_1736), .in1(s_95_1751) );
  Fadder_ A_95_1756( .carry(c_95_1756), .sum(s_95_1756), .in3(c_94_1737), .in2(s_95_1752), .in1(s_95_1753) );
  Fadder_ A_95_1757( .carry(c_95_1757), .sum(s_95_1757), .in3(c_94_1738), .in2(s_95_1754), .in1(c_94_1739) );
  Fadder_ A_95_1758( .carry(c_95_1758), .sum(s_95_1758), .in3(s_95_1755), .in2(c_94_1740), .in1(s_95_1756) );
  Fadder_ A_95_1759( .carry(c_95_1759), .sum(s_95_1759), .in3(c_94_1741), .in2(s_95_1757), .in1(c_94_1742) );
  Fadder_ A_95_1760( .carry(c[95]), .sum(s[95]), .in3(s_95_1758), .in2(c_94_1743), .in1(s_95_1759) );

  // ***** Bit 96 ***** //
  Hadder_ A_96_1761( .carry(c_96_1761), .sum(s_96_1761), .in2(sign_), .in1(P_31[34]) );
  Fadder_ A_96_1762( .carry(c_96_1762), .sum(s_96_1762), .in3(P_30[36]), .in2(P_29[38]), .in1(P_28[40]) );
  Fadder_ A_96_1763( .carry(c_96_1763), .sum(s_96_1763), .in3(P_27[42]), .in2(P_26[44]), .in1(P_25[46]) );
  Fadder_ A_96_1764( .carry(c_96_1764), .sum(s_96_1764), .in3(P_24[48]), .in2(P_23[50]), .in1(P_22[52]) );
  Fadder_ A_96_1765( .carry(c_96_1765), .sum(s_96_1765), .in3(P_21[54]), .in2(P_20[56]), .in1(P_19[58]) );
  Fadder_ A_96_1766( .carry(c_96_1766), .sum(s_96_1766), .in3(P_18[60]), .in2(P_17[62]), .in1(P_16[64]) );
  Fadder_ A_96_1767( .carry(c_96_1767), .sum(s_96_1767), .in3(c_95_1749), .in2(c_95_1748), .in1(c_95_1747) );
  Fadder_ A_96_1768( .carry(c_96_1768), .sum(s_96_1768), .in3(c_95_1746), .in2(c_95_1745), .in1(s_96_1761) );
  Fadder_ A_96_1769( .carry(c_96_1769), .sum(s_96_1769), .in3(s_96_1766), .in2(s_96_1765), .in1(s_96_1764) );
  Fadder_ A_96_1770( .carry(c_96_1770), .sum(s_96_1770), .in3(s_96_1763), .in2(s_96_1762), .in1(c_95_1750) );
  Fadder_ A_96_1771( .carry(c_96_1771), .sum(s_96_1771), .in3(c_95_1751), .in2(c_95_1752), .in1(s_96_1767) );
  Fadder_ A_96_1772( .carry(c_96_1772), .sum(s_96_1772), .in3(c_95_1753), .in2(s_96_1768), .in1(s_96_1769) );
  Fadder_ A_96_1773( .carry(c_96_1773), .sum(s_96_1773), .in3(s_96_1770), .in2(c_95_1754), .in1(c_95_1755) );
  Fadder_ A_96_1774( .carry(c_96_1774), .sum(s_96_1774), .in3(s_96_1771), .in2(c_95_1756), .in1(s_96_1772) );
  Fadder_ A_96_1775( .carry(c_96_1775), .sum(s_96_1775), .in3(c_95_1757), .in2(s_96_1773), .in1(c_95_1758) );
  Fadder_ A_96_1776( .carry(c[96]), .sum(s[96]), .in3(s_96_1774), .in2(c_95_1759), .in1(s_96_1775) );

  // ***** Bit 97 ***** //
  Fadder_ A_97_1777( .carry(c_97_1777), .sum(s_97_1777), .in3(P_31[35]), .in2(P_30[37]), .in1(P_29[39]) );
  Fadder_ A_97_1778( .carry(c_97_1778), .sum(s_97_1778), .in3(P_28[41]), .in2(P_27[43]), .in1(P_26[45]) );
  Fadder_ A_97_1779( .carry(c_97_1779), .sum(s_97_1779), .in3(P_25[47]), .in2(P_24[49]), .in1(P_23[51]) );
  Fadder_ A_97_1780( .carry(c_97_1780), .sum(s_97_1780), .in3(P_22[53]), .in2(P_21[55]), .in1(P_20[57]) );
  Fadder_ A_97_1781( .carry(c_97_1781), .sum(s_97_1781), .in3(P_19[59]), .in2(P_18[61]), .in1(P_17[63]) );
  Fadder_ A_97_1782( .carry(c_97_1782), .sum(s_97_1782), .in3(P_16[65]), .in2(c_96_1761), .in1(c_96_1766) );
  Fadder_ A_97_1783( .carry(c_97_1783), .sum(s_97_1783), .in3(c_96_1765), .in2(c_96_1764), .in1(c_96_1763) );
  Fadder_ A_97_1784( .carry(c_97_1784), .sum(s_97_1784), .in3(c_96_1762), .in2(s_97_1781), .in1(s_97_1780) );
  Fadder_ A_97_1785( .carry(c_97_1785), .sum(s_97_1785), .in3(s_97_1779), .in2(s_97_1778), .in1(s_97_1777) );
  Fadder_ A_97_1786( .carry(c_97_1786), .sum(s_97_1786), .in3(c_96_1768), .in2(c_96_1767), .in1(s_97_1782) );
  Fadder_ A_97_1787( .carry(c_97_1787), .sum(s_97_1787), .in3(s_97_1783), .in2(c_96_1769), .in1(c_96_1770) );
  Fadder_ A_97_1788( .carry(c_97_1788), .sum(s_97_1788), .in3(s_97_1784), .in2(s_97_1785), .in1(c_96_1771) );
  Fadder_ A_97_1789( .carry(c_97_1789), .sum(s_97_1789), .in3(c_96_1772), .in2(s_97_1786), .in1(s_97_1787) );
  Fadder_ A_97_1790( .carry(c_97_1790), .sum(s_97_1790), .in3(c_96_1773), .in2(s_97_1788), .in1(c_96_1774) );
  Fadder_ A_97_1791( .carry(c[97]), .sum(s[97]), .in3(s_97_1789), .in2(c_96_1775), .in1(s_97_1790) );

  // ***** Bit 98 ***** //
  Hadder_ A_98_1792( .carry(c_98_1792), .sum(s_98_1792), .in2(sign_), .in1(P_31[36]) );
  Fadder_ A_98_1793( .carry(c_98_1793), .sum(s_98_1793), .in3(P_30[38]), .in2(P_29[40]), .in1(P_28[42]) );
  Fadder_ A_98_1794( .carry(c_98_1794), .sum(s_98_1794), .in3(P_27[44]), .in2(P_26[46]), .in1(P_25[48]) );
  Fadder_ A_98_1795( .carry(c_98_1795), .sum(s_98_1795), .in3(P_24[50]), .in2(P_23[52]), .in1(P_22[54]) );
  Fadder_ A_98_1796( .carry(c_98_1796), .sum(s_98_1796), .in3(P_21[56]), .in2(P_20[58]), .in1(P_19[60]) );
  Fadder_ A_98_1797( .carry(c_98_1797), .sum(s_98_1797), .in3(P_18[62]), .in2(P_17[64]), .in1(c_97_1781) );
  Fadder_ A_98_1798( .carry(c_98_1798), .sum(s_98_1798), .in3(c_97_1780), .in2(c_97_1779), .in1(c_97_1778) );
  Fadder_ A_98_1799( .carry(c_98_1799), .sum(s_98_1799), .in3(c_97_1777), .in2(s_98_1792), .in1(s_98_1796) );
  Fadder_ A_98_1800( .carry(c_98_1800), .sum(s_98_1800), .in3(s_98_1795), .in2(s_98_1794), .in1(s_98_1793) );
  Fadder_ A_98_1801( .carry(c_98_1801), .sum(s_98_1801), .in3(c_97_1782), .in2(c_97_1783), .in1(s_98_1797) );
  Fadder_ A_98_1802( .carry(c_98_1802), .sum(s_98_1802), .in3(s_98_1798), .in2(c_97_1785), .in1(c_97_1784) );
  Fadder_ A_98_1803( .carry(c_98_1803), .sum(s_98_1803), .in3(s_98_1799), .in2(s_98_1800), .in1(c_97_1786) );
  Fadder_ A_98_1804( .carry(c_98_1804), .sum(s_98_1804), .in3(c_97_1787), .in2(s_98_1801), .in1(s_98_1802) );
  Fadder_ A_98_1805( .carry(c_98_1805), .sum(s_98_1805), .in3(c_97_1788), .in2(s_98_1803), .in1(c_97_1789) );
  Fadder_ A_98_1806( .carry(c[98]), .sum(s[98]), .in3(s_98_1804), .in2(c_97_1790), .in1(s_98_1805) );

  // ***** Bit 99 ***** //
  Fadder_ A_99_1807( .carry(c_99_1807), .sum(s_99_1807), .in3(P_31[37]), .in2(P_30[39]), .in1(P_29[41]) );
  Fadder_ A_99_1808( .carry(c_99_1808), .sum(s_99_1808), .in3(P_28[43]), .in2(P_27[45]), .in1(P_26[47]) );
  Fadder_ A_99_1809( .carry(c_99_1809), .sum(s_99_1809), .in3(P_25[49]), .in2(P_24[51]), .in1(P_23[53]) );
  Fadder_ A_99_1810( .carry(c_99_1810), .sum(s_99_1810), .in3(P_22[55]), .in2(P_21[57]), .in1(P_20[59]) );
  Fadder_ A_99_1811( .carry(c_99_1811), .sum(s_99_1811), .in3(P_19[61]), .in2(P_18[63]), .in1(P_17[65]) );
  Fadder_ A_99_1812( .carry(c_99_1812), .sum(s_99_1812), .in3(c_98_1792), .in2(c_98_1796), .in1(c_98_1795) );
  Fadder_ A_99_1813( .carry(c_99_1813), .sum(s_99_1813), .in3(c_98_1794), .in2(c_98_1793), .in1(s_99_1811) );
  Fadder_ A_99_1814( .carry(c_99_1814), .sum(s_99_1814), .in3(s_99_1810), .in2(s_99_1809), .in1(s_99_1808) );
  Fadder_ A_99_1815( .carry(c_99_1815), .sum(s_99_1815), .in3(s_99_1807), .in2(c_98_1797), .in1(c_98_1798) );
  Fadder_ A_99_1816( .carry(c_99_1816), .sum(s_99_1816), .in3(c_98_1799), .in2(s_99_1812), .in1(c_98_1800) );
  Fadder_ A_99_1817( .carry(c_99_1817), .sum(s_99_1817), .in3(s_99_1813), .in2(s_99_1814), .in1(c_98_1801) );
  Fadder_ A_99_1818( .carry(c_99_1818), .sum(s_99_1818), .in3(s_99_1815), .in2(c_98_1802), .in1(s_99_1816) );
  Fadder_ A_99_1819( .carry(c_99_1819), .sum(s_99_1819), .in3(c_98_1803), .in2(s_99_1817), .in1(c_98_1804) );
  Fadder_ A_99_1820( .carry(c[99]), .sum(s[99]), .in3(s_99_1818), .in2(c_98_1805), .in1(s_99_1819) );

  // ***** Bit 100 ***** //
  Hadder_ A_100_1821( .carry(c_100_1821), .sum(s_100_1821), .in2(sign_), .in1(P_31[38]) );
  Fadder_ A_100_1822( .carry(c_100_1822), .sum(s_100_1822), .in3(P_30[40]), .in2(P_29[42]), .in1(P_28[44]) );
  Fadder_ A_100_1823( .carry(c_100_1823), .sum(s_100_1823), .in3(P_27[46]), .in2(P_26[48]), .in1(P_25[50]) );
  Fadder_ A_100_1824( .carry(c_100_1824), .sum(s_100_1824), .in3(P_24[52]), .in2(P_23[54]), .in1(P_22[56]) );
  Fadder_ A_100_1825( .carry(c_100_1825), .sum(s_100_1825), .in3(P_21[58]), .in2(P_20[60]), .in1(P_19[62]) );
  Fadder_ A_100_1826( .carry(c_100_1826), .sum(s_100_1826), .in3(P_18[64]), .in2(c_99_1811), .in1(c_99_1810) );
  Fadder_ A_100_1827( .carry(c_100_1827), .sum(s_100_1827), .in3(c_99_1809), .in2(c_99_1808), .in1(c_99_1807) );
  Fadder_ A_100_1828( .carry(c_100_1828), .sum(s_100_1828), .in3(s_100_1821), .in2(s_100_1825), .in1(s_100_1824) );
  Fadder_ A_100_1829( .carry(c_100_1829), .sum(s_100_1829), .in3(s_100_1823), .in2(s_100_1822), .in1(c_99_1812) );
  Fadder_ A_100_1830( .carry(c_100_1830), .sum(s_100_1830), .in3(c_99_1813), .in2(s_100_1826), .in1(s_100_1827) );
  Fadder_ A_100_1831( .carry(c_100_1831), .sum(s_100_1831), .in3(c_99_1814), .in2(s_100_1828), .in1(c_99_1815) );
  Fadder_ A_100_1832( .carry(c_100_1832), .sum(s_100_1832), .in3(s_100_1829), .in2(c_99_1816), .in1(s_100_1830) );
  Fadder_ A_100_1833( .carry(c_100_1833), .sum(s_100_1833), .in3(c_99_1817), .in2(s_100_1831), .in1(c_99_1818) );
  Fadder_ A_100_1834( .carry(c[100]), .sum(s[100]), .in3(s_100_1832), .in2(c_99_1819), .in1(s_100_1833) );

  // ***** Bit 101 ***** //
  Fadder_ A_101_1835( .carry(c_101_1835), .sum(s_101_1835), .in3(P_31[39]), .in2(P_30[41]), .in1(P_29[43]) );
  Fadder_ A_101_1836( .carry(c_101_1836), .sum(s_101_1836), .in3(P_28[45]), .in2(P_27[47]), .in1(P_26[49]) );
  Fadder_ A_101_1837( .carry(c_101_1837), .sum(s_101_1837), .in3(P_25[51]), .in2(P_24[53]), .in1(P_23[55]) );
  Fadder_ A_101_1838( .carry(c_101_1838), .sum(s_101_1838), .in3(P_22[57]), .in2(P_21[59]), .in1(P_20[61]) );
  Fadder_ A_101_1839( .carry(c_101_1839), .sum(s_101_1839), .in3(P_19[63]), .in2(P_18[65]), .in1(c_100_1821) );
  Fadder_ A_101_1840( .carry(c_101_1840), .sum(s_101_1840), .in3(c_100_1825), .in2(c_100_1824), .in1(c_100_1823) );
  Fadder_ A_101_1841( .carry(c_101_1841), .sum(s_101_1841), .in3(c_100_1822), .in2(s_101_1838), .in1(s_101_1837) );
  Fadder_ A_101_1842( .carry(c_101_1842), .sum(s_101_1842), .in3(s_101_1836), .in2(s_101_1835), .in1(s_101_1839) );
  Fadder_ A_101_1843( .carry(c_101_1843), .sum(s_101_1843), .in3(c_100_1827), .in2(c_100_1826), .in1(s_101_1840) );
  Fadder_ A_101_1844( .carry(c_101_1844), .sum(s_101_1844), .in3(c_100_1828), .in2(s_101_1841), .in1(s_101_1842) );
  Fadder_ A_101_1845( .carry(c_101_1845), .sum(s_101_1845), .in3(c_100_1829), .in2(c_100_1830), .in1(s_101_1843) );
  Fadder_ A_101_1846( .carry(c_101_1846), .sum(s_101_1846), .in3(c_100_1831), .in2(s_101_1844), .in1(c_100_1832) );
  Fadder_ A_101_1847( .carry(c[101]), .sum(s[101]), .in3(s_101_1845), .in2(c_100_1833), .in1(s_101_1846) );

  // ***** Bit 102 ***** //
  Hadder_ A_102_1848( .carry(c_102_1848), .sum(s_102_1848), .in2(sign_), .in1(P_31[40]) );
  Fadder_ A_102_1849( .carry(c_102_1849), .sum(s_102_1849), .in3(P_30[42]), .in2(P_29[44]), .in1(P_28[46]) );
  Fadder_ A_102_1850( .carry(c_102_1850), .sum(s_102_1850), .in3(P_27[48]), .in2(P_26[50]), .in1(P_25[52]) );
  Fadder_ A_102_1851( .carry(c_102_1851), .sum(s_102_1851), .in3(P_24[54]), .in2(P_23[56]), .in1(P_22[58]) );
  Fadder_ A_102_1852( .carry(c_102_1852), .sum(s_102_1852), .in3(P_21[60]), .in2(P_20[62]), .in1(P_19[64]) );
  Fadder_ A_102_1853( .carry(c_102_1853), .sum(s_102_1853), .in3(c_101_1838), .in2(c_101_1837), .in1(c_101_1836) );
  Fadder_ A_102_1854( .carry(c_102_1854), .sum(s_102_1854), .in3(c_101_1835), .in2(s_102_1848), .in1(s_102_1852) );
  Fadder_ A_102_1855( .carry(c_102_1855), .sum(s_102_1855), .in3(s_102_1851), .in2(s_102_1850), .in1(s_102_1849) );
  Fadder_ A_102_1856( .carry(c_102_1856), .sum(s_102_1856), .in3(c_101_1839), .in2(c_101_1840), .in1(s_102_1853) );
  Fadder_ A_102_1857( .carry(c_102_1857), .sum(s_102_1857), .in3(c_101_1841), .in2(s_102_1854), .in1(s_102_1855) );
  Fadder_ A_102_1858( .carry(c_102_1858), .sum(s_102_1858), .in3(c_101_1842), .in2(c_101_1843), .in1(s_102_1856) );
  Fadder_ A_102_1859( .carry(c_102_1859), .sum(s_102_1859), .in3(s_102_1857), .in2(c_101_1844), .in1(c_101_1845) );
  Fadder_ A_102_1860( .carry(c[102]), .sum(s[102]), .in3(s_102_1858), .in2(c_101_1846), .in1(s_102_1859) );

  // ***** Bit 103 ***** //
  Fadder_ A_103_1861( .carry(c_103_1861), .sum(s_103_1861), .in3(P_31[41]), .in2(P_30[43]), .in1(P_29[45]) );
  Fadder_ A_103_1862( .carry(c_103_1862), .sum(s_103_1862), .in3(P_28[47]), .in2(P_27[49]), .in1(P_26[51]) );
  Fadder_ A_103_1863( .carry(c_103_1863), .sum(s_103_1863), .in3(P_25[53]), .in2(P_24[55]), .in1(P_23[57]) );
  Fadder_ A_103_1864( .carry(c_103_1864), .sum(s_103_1864), .in3(P_22[59]), .in2(P_21[61]), .in1(P_20[63]) );
  Fadder_ A_103_1865( .carry(c_103_1865), .sum(s_103_1865), .in3(P_19[65]), .in2(c_102_1848), .in1(c_102_1852) );
  Fadder_ A_103_1866( .carry(c_103_1866), .sum(s_103_1866), .in3(c_102_1851), .in2(c_102_1850), .in1(c_102_1849) );
  Fadder_ A_103_1867( .carry(c_103_1867), .sum(s_103_1867), .in3(s_103_1864), .in2(s_103_1863), .in1(s_103_1862) );
  Fadder_ A_103_1868( .carry(c_103_1868), .sum(s_103_1868), .in3(s_103_1861), .in2(c_102_1853), .in1(c_102_1854) );
  Fadder_ A_103_1869( .carry(c_103_1869), .sum(s_103_1869), .in3(s_103_1865), .in2(s_103_1866), .in1(c_102_1855) );
  Fadder_ A_103_1870( .carry(c_103_1870), .sum(s_103_1870), .in3(s_103_1867), .in2(c_102_1856), .in1(s_103_1868) );
  Fadder_ A_103_1871( .carry(c_103_1871), .sum(s_103_1871), .in3(s_103_1869), .in2(c_102_1857), .in1(c_102_1858) );
  Fadder_ A_103_1872( .carry(c[103]), .sum(s[103]), .in3(s_103_1870), .in2(c_102_1859), .in1(s_103_1871) );

  // ***** Bit 104 ***** //
  Hadder_ A_104_1873( .carry(c_104_1873), .sum(s_104_1873), .in2(sign_), .in1(P_31[42]) );
  Fadder_ A_104_1874( .carry(c_104_1874), .sum(s_104_1874), .in3(P_30[44]), .in2(P_29[46]), .in1(P_28[48]) );
  Fadder_ A_104_1875( .carry(c_104_1875), .sum(s_104_1875), .in3(P_27[50]), .in2(P_26[52]), .in1(P_25[54]) );
  Fadder_ A_104_1876( .carry(c_104_1876), .sum(s_104_1876), .in3(P_24[56]), .in2(P_23[58]), .in1(P_22[60]) );
  Fadder_ A_104_1877( .carry(c_104_1877), .sum(s_104_1877), .in3(P_21[62]), .in2(P_20[64]), .in1(c_103_1864) );
  Fadder_ A_104_1878( .carry(c_104_1878), .sum(s_104_1878), .in3(c_103_1863), .in2(c_103_1862), .in1(c_103_1861) );
  Fadder_ A_104_1879( .carry(c_104_1879), .sum(s_104_1879), .in3(s_104_1873), .in2(s_104_1876), .in1(s_104_1875) );
  Fadder_ A_104_1880( .carry(c_104_1880), .sum(s_104_1880), .in3(s_104_1874), .in2(c_103_1865), .in1(c_103_1866) );
  Fadder_ A_104_1881( .carry(c_104_1881), .sum(s_104_1881), .in3(s_104_1877), .in2(s_104_1878), .in1(c_103_1867) );
  Fadder_ A_104_1882( .carry(c_104_1882), .sum(s_104_1882), .in3(s_104_1879), .in2(c_103_1868), .in1(s_104_1880) );
  Fadder_ A_104_1883( .carry(c_104_1883), .sum(s_104_1883), .in3(c_103_1869), .in2(s_104_1881), .in1(c_103_1870) );
  Fadder_ A_104_1884( .carry(c[104]), .sum(s[104]), .in3(s_104_1882), .in2(c_103_1871), .in1(s_104_1883) );

  // ***** Bit 105 ***** //
  Fadder_ A_105_1885( .carry(c_105_1885), .sum(s_105_1885), .in3(P_31[43]), .in2(P_30[45]), .in1(P_29[47]) );
  Fadder_ A_105_1886( .carry(c_105_1886), .sum(s_105_1886), .in3(P_28[49]), .in2(P_27[51]), .in1(P_26[53]) );
  Fadder_ A_105_1887( .carry(c_105_1887), .sum(s_105_1887), .in3(P_25[55]), .in2(P_24[57]), .in1(P_23[59]) );
  Fadder_ A_105_1888( .carry(c_105_1888), .sum(s_105_1888), .in3(P_22[61]), .in2(P_21[63]), .in1(P_20[65]) );
  Fadder_ A_105_1889( .carry(c_105_1889), .sum(s_105_1889), .in3(c_104_1873), .in2(c_104_1876), .in1(c_104_1875) );
  Fadder_ A_105_1890( .carry(c_105_1890), .sum(s_105_1890), .in3(c_104_1874), .in2(s_105_1888), .in1(s_105_1887) );
  Fadder_ A_105_1891( .carry(c_105_1891), .sum(s_105_1891), .in3(s_105_1886), .in2(s_105_1885), .in1(c_104_1877) );
  Fadder_ A_105_1892( .carry(c_105_1892), .sum(s_105_1892), .in3(c_104_1878), .in2(s_105_1889), .in1(c_104_1879) );
  Fadder_ A_105_1893( .carry(c_105_1893), .sum(s_105_1893), .in3(s_105_1890), .in2(c_104_1880), .in1(s_105_1891) );
  Fadder_ A_105_1894( .carry(c_105_1894), .sum(s_105_1894), .in3(c_104_1881), .in2(s_105_1892), .in1(c_104_1882) );
  Fadder_ A_105_1895( .carry(c[105]), .sum(s[105]), .in3(s_105_1893), .in2(c_104_1883), .in1(s_105_1894) );

  // ***** Bit 106 ***** //
  Hadder_ A_106_1896( .carry(c_106_1896), .sum(s_106_1896), .in2(sign_), .in1(P_31[44]) );
  Fadder_ A_106_1897( .carry(c_106_1897), .sum(s_106_1897), .in3(P_30[46]), .in2(P_29[48]), .in1(P_28[50]) );
  Fadder_ A_106_1898( .carry(c_106_1898), .sum(s_106_1898), .in3(P_27[52]), .in2(P_26[54]), .in1(P_25[56]) );
  Fadder_ A_106_1899( .carry(c_106_1899), .sum(s_106_1899), .in3(P_24[58]), .in2(P_23[60]), .in1(P_22[62]) );
  Fadder_ A_106_1900( .carry(c_106_1900), .sum(s_106_1900), .in3(P_21[64]), .in2(c_105_1888), .in1(c_105_1887) );
  Fadder_ A_106_1901( .carry(c_106_1901), .sum(s_106_1901), .in3(c_105_1886), .in2(c_105_1885), .in1(s_106_1896) );
  Fadder_ A_106_1902( .carry(c_106_1902), .sum(s_106_1902), .in3(s_106_1899), .in2(s_106_1898), .in1(s_106_1897) );
  Fadder_ A_106_1903( .carry(c_106_1903), .sum(s_106_1903), .in3(c_105_1889), .in2(s_106_1900), .in1(c_105_1890) );
  Fadder_ A_106_1904( .carry(c_106_1904), .sum(s_106_1904), .in3(s_106_1901), .in2(s_106_1902), .in1(c_105_1891) );
  Fadder_ A_106_1905( .carry(c_106_1905), .sum(s_106_1905), .in3(c_105_1892), .in2(s_106_1903), .in1(s_106_1904) );
  Fadder_ A_106_1906( .carry(c[106]), .sum(s[106]), .in3(c_105_1893), .in2(c_105_1894), .in1(s_106_1905) );

  // ***** Bit 107 ***** //
  Fadder_ A_107_1907( .carry(c_107_1907), .sum(s_107_1907), .in3(P_31[45]), .in2(P_30[47]), .in1(P_29[49]) );
  Fadder_ A_107_1908( .carry(c_107_1908), .sum(s_107_1908), .in3(P_28[51]), .in2(P_27[53]), .in1(P_26[55]) );
  Fadder_ A_107_1909( .carry(c_107_1909), .sum(s_107_1909), .in3(P_25[57]), .in2(P_24[59]), .in1(P_23[61]) );
  Fadder_ A_107_1910( .carry(c_107_1910), .sum(s_107_1910), .in3(P_22[63]), .in2(P_21[65]), .in1(c_106_1896) );
  Fadder_ A_107_1911( .carry(c_107_1911), .sum(s_107_1911), .in3(c_106_1899), .in2(c_106_1898), .in1(c_106_1897) );
  Fadder_ A_107_1912( .carry(c_107_1912), .sum(s_107_1912), .in3(s_107_1909), .in2(s_107_1908), .in1(s_107_1907) );
  Fadder_ A_107_1913( .carry(c_107_1913), .sum(s_107_1913), .in3(s_107_1910), .in2(c_106_1901), .in1(c_106_1900) );
  Fadder_ A_107_1914( .carry(c_107_1914), .sum(s_107_1914), .in3(s_107_1911), .in2(c_106_1902), .in1(s_107_1912) );
  Fadder_ A_107_1915( .carry(c_107_1915), .sum(s_107_1915), .in3(s_107_1913), .in2(c_106_1903), .in1(c_106_1904) );
  Fadder_ A_107_1916( .carry(c[107]), .sum(s[107]), .in3(s_107_1914), .in2(s_107_1915), .in1(c_106_1905) );

  // ***** Bit 108 ***** //
  Hadder_ A_108_1917( .carry(c_108_1917), .sum(s_108_1917), .in2(sign_), .in1(P_31[46]) );
  Fadder_ A_108_1918( .carry(c_108_1918), .sum(s_108_1918), .in3(P_30[48]), .in2(P_29[50]), .in1(P_28[52]) );
  Fadder_ A_108_1919( .carry(c_108_1919), .sum(s_108_1919), .in3(P_27[54]), .in2(P_26[56]), .in1(P_25[58]) );
  Fadder_ A_108_1920( .carry(c_108_1920), .sum(s_108_1920), .in3(P_24[60]), .in2(P_23[62]), .in1(P_22[64]) );
  Fadder_ A_108_1921( .carry(c_108_1921), .sum(s_108_1921), .in3(c_107_1909), .in2(c_107_1908), .in1(c_107_1907) );
  Fadder_ A_108_1922( .carry(c_108_1922), .sum(s_108_1922), .in3(s_108_1917), .in2(s_108_1920), .in1(s_108_1919) );
  Fadder_ A_108_1923( .carry(c_108_1923), .sum(s_108_1923), .in3(s_108_1918), .in2(c_107_1910), .in1(c_107_1911) );
  Fadder_ A_108_1924( .carry(c_108_1924), .sum(s_108_1924), .in3(s_108_1921), .in2(c_107_1912), .in1(s_108_1922) );
  Fadder_ A_108_1925( .carry(c_108_1925), .sum(s_108_1925), .in3(c_107_1913), .in2(s_108_1923), .in1(c_107_1914) );
  Fadder_ A_108_1926( .carry(c[108]), .sum(s[108]), .in3(s_108_1924), .in2(c_107_1915), .in1(s_108_1925) );

  // ***** Bit 109 ***** //
  Fadder_ A_109_1927( .carry(c_109_1927), .sum(s_109_1927), .in3(P_31[47]), .in2(P_30[49]), .in1(P_29[51]) );
  Fadder_ A_109_1928( .carry(c_109_1928), .sum(s_109_1928), .in3(P_28[53]), .in2(P_27[55]), .in1(P_26[57]) );
  Fadder_ A_109_1929( .carry(c_109_1929), .sum(s_109_1929), .in3(P_25[59]), .in2(P_24[61]), .in1(P_23[63]) );
  Fadder_ A_109_1930( .carry(c_109_1930), .sum(s_109_1930), .in3(P_22[65]), .in2(c_108_1917), .in1(c_108_1920) );
  Fadder_ A_109_1931( .carry(c_109_1931), .sum(s_109_1931), .in3(c_108_1919), .in2(c_108_1918), .in1(s_109_1929) );
  Fadder_ A_109_1932( .carry(c_109_1932), .sum(s_109_1932), .in3(s_109_1928), .in2(s_109_1927), .in1(c_108_1921) );
  Fadder_ A_109_1933( .carry(c_109_1933), .sum(s_109_1933), .in3(s_109_1930), .in2(c_108_1922), .in1(s_109_1931) );
  Fadder_ A_109_1934( .carry(c_109_1934), .sum(s_109_1934), .in3(c_108_1923), .in2(s_109_1932), .in1(c_108_1924) );
  Fadder_ A_109_1935( .carry(c[109]), .sum(s[109]), .in3(s_109_1933), .in2(c_108_1925), .in1(s_109_1934) );

  // ***** Bit 110 ***** //
  Hadder_ A_110_1936( .carry(c_110_1936), .sum(s_110_1936), .in2(sign_), .in1(P_31[48]) );
  Fadder_ A_110_1937( .carry(c_110_1937), .sum(s_110_1937), .in3(P_30[50]), .in2(P_29[52]), .in1(P_28[54]) );
  Fadder_ A_110_1938( .carry(c_110_1938), .sum(s_110_1938), .in3(P_27[56]), .in2(P_26[58]), .in1(P_25[60]) );
  Fadder_ A_110_1939( .carry(c_110_1939), .sum(s_110_1939), .in3(P_24[62]), .in2(P_23[64]), .in1(c_109_1929) );
  Fadder_ A_110_1940( .carry(c_110_1940), .sum(s_110_1940), .in3(c_109_1928), .in2(c_109_1927), .in1(s_110_1936) );
  Fadder_ A_110_1941( .carry(c_110_1941), .sum(s_110_1941), .in3(s_110_1938), .in2(s_110_1937), .in1(c_109_1930) );
  Fadder_ A_110_1942( .carry(c_110_1942), .sum(s_110_1942), .in3(c_109_1931), .in2(s_110_1939), .in1(s_110_1940) );
  Fadder_ A_110_1943( .carry(c_110_1943), .sum(s_110_1943), .in3(c_109_1932), .in2(s_110_1941), .in1(c_109_1933) );
  Fadder_ A_110_1944( .carry(c[110]), .sum(s[110]), .in3(s_110_1942), .in2(c_109_1934), .in1(s_110_1943) );

  // ***** Bit 111 ***** //
  Fadder_ A_111_1945( .carry(c_111_1945), .sum(s_111_1945), .in3(P_31[49]), .in2(P_30[51]), .in1(P_29[53]) );
  Fadder_ A_111_1946( .carry(c_111_1946), .sum(s_111_1946), .in3(P_28[55]), .in2(P_27[57]), .in1(P_26[59]) );
  Fadder_ A_111_1947( .carry(c_111_1947), .sum(s_111_1947), .in3(P_25[61]), .in2(P_24[63]), .in1(P_23[65]) );
  Fadder_ A_111_1948( .carry(c_111_1948), .sum(s_111_1948), .in3(c_110_1936), .in2(c_110_1938), .in1(c_110_1937) );
  Fadder_ A_111_1949( .carry(c_111_1949), .sum(s_111_1949), .in3(s_111_1947), .in2(s_111_1946), .in1(s_111_1945) );
  Fadder_ A_111_1950( .carry(c_111_1950), .sum(s_111_1950), .in3(c_110_1939), .in2(c_110_1940), .in1(s_111_1948) );
  Fadder_ A_111_1951( .carry(c_111_1951), .sum(s_111_1951), .in3(s_111_1949), .in2(c_110_1941), .in1(c_110_1942) );
  Fadder_ A_111_1952( .carry(c[111]), .sum(s[111]), .in3(s_111_1950), .in2(c_110_1943), .in1(s_111_1951) );

  // ***** Bit 112 ***** //
  Hadder_ A_112_1953( .carry(c_112_1953), .sum(s_112_1953), .in2(sign_), .in1(P_31[50]) );
  Fadder_ A_112_1954( .carry(c_112_1954), .sum(s_112_1954), .in3(P_30[52]), .in2(P_29[54]), .in1(P_28[56]) );
  Fadder_ A_112_1955( .carry(c_112_1955), .sum(s_112_1955), .in3(P_27[58]), .in2(P_26[60]), .in1(P_25[62]) );
  Fadder_ A_112_1956( .carry(c_112_1956), .sum(s_112_1956), .in3(P_24[64]), .in2(c_111_1947), .in1(c_111_1946) );
  Fadder_ A_112_1957( .carry(c_112_1957), .sum(s_112_1957), .in3(c_111_1945), .in2(s_112_1953), .in1(s_112_1955) );
  Fadder_ A_112_1958( .carry(c_112_1958), .sum(s_112_1958), .in3(s_112_1954), .in2(c_111_1948), .in1(s_112_1956) );
  Fadder_ A_112_1959( .carry(c_112_1959), .sum(s_112_1959), .in3(c_111_1949), .in2(s_112_1957), .in1(c_111_1950) );
  Fadder_ A_112_1960( .carry(c[112]), .sum(s[112]), .in3(s_112_1958), .in2(c_111_1951), .in1(s_112_1959) );

  // ***** Bit 113 ***** //
  Fadder_ A_113_1961( .carry(c_113_1961), .sum(s_113_1961), .in3(P_31[51]), .in2(P_30[53]), .in1(P_29[55]) );
  Fadder_ A_113_1962( .carry(c_113_1962), .sum(s_113_1962), .in3(P_28[57]), .in2(P_27[59]), .in1(P_26[61]) );
  Fadder_ A_113_1963( .carry(c_113_1963), .sum(s_113_1963), .in3(P_25[63]), .in2(P_24[65]), .in1(c_112_1953) );
  Fadder_ A_113_1964( .carry(c_113_1964), .sum(s_113_1964), .in3(c_112_1955), .in2(c_112_1954), .in1(s_113_1962) );
  Fadder_ A_113_1965( .carry(c_113_1965), .sum(s_113_1965), .in3(s_113_1961), .in2(s_113_1963), .in1(c_112_1956) );
  Fadder_ A_113_1966( .carry(c_113_1966), .sum(s_113_1966), .in3(c_112_1957), .in2(s_113_1964), .in1(c_112_1958) );
  Fadder_ A_113_1967( .carry(c[113]), .sum(s[113]), .in3(s_113_1965), .in2(c_112_1959), .in1(s_113_1966) );

  // ***** Bit 114 ***** //
  Hadder_ A_114_1968( .carry(c_114_1968), .sum(s_114_1968), .in2(sign_), .in1(P_31[52]) );
  Fadder_ A_114_1969( .carry(c_114_1969), .sum(s_114_1969), .in3(P_30[54]), .in2(P_29[56]), .in1(P_28[58]) );
  Fadder_ A_114_1970( .carry(c_114_1970), .sum(s_114_1970), .in3(P_27[60]), .in2(P_26[62]), .in1(P_25[64]) );
  Fadder_ A_114_1971( .carry(c_114_1971), .sum(s_114_1971), .in3(c_113_1962), .in2(c_113_1961), .in1(s_114_1968) );
  Fadder_ A_114_1972( .carry(c_114_1972), .sum(s_114_1972), .in3(s_114_1970), .in2(s_114_1969), .in1(c_113_1963) );
  Fadder_ A_114_1973( .carry(c_114_1973), .sum(s_114_1973), .in3(c_113_1964), .in2(s_114_1971), .in1(s_114_1972) );
  Fadder_ A_114_1974( .carry(c[114]), .sum(s[114]), .in3(c_113_1965), .in2(s_114_1973), .in1(c_113_1966) );

  // ***** Bit 115 ***** //
  Fadder_ A_115_1975( .carry(c_115_1975), .sum(s_115_1975), .in3(P_31[53]), .in2(P_30[55]), .in1(P_29[57]) );
  Fadder_ A_115_1976( .carry(c_115_1976), .sum(s_115_1976), .in3(P_28[59]), .in2(P_27[61]), .in1(P_26[63]) );
  Fadder_ A_115_1977( .carry(c_115_1977), .sum(s_115_1977), .in3(P_25[65]), .in2(c_114_1968), .in1(c_114_1970) );
  Fadder_ A_115_1978( .carry(c_115_1978), .sum(s_115_1978), .in3(c_114_1969), .in2(s_115_1976), .in1(s_115_1975) );
  Fadder_ A_115_1979( .carry(c_115_1979), .sum(s_115_1979), .in3(c_114_1971), .in2(s_115_1977), .in1(c_114_1972) );
  Fadder_ A_115_1980( .carry(c[115]), .sum(s[115]), .in3(s_115_1978), .in2(s_115_1979), .in1(c_114_1973) );

  // ***** Bit 116 ***** //
  Hadder_ A_116_1981( .carry(c_116_1981), .sum(s_116_1981), .in2(sign_), .in1(P_31[54]) );
  Fadder_ A_116_1982( .carry(c_116_1982), .sum(s_116_1982), .in3(P_30[56]), .in2(P_29[58]), .in1(P_28[60]) );
  Fadder_ A_116_1983( .carry(c_116_1983), .sum(s_116_1983), .in3(P_27[62]), .in2(P_26[64]), .in1(c_115_1976) );
  Fadder_ A_116_1984( .carry(c_116_1984), .sum(s_116_1984), .in3(c_115_1975), .in2(s_116_1981), .in1(s_116_1982) );
  Fadder_ A_116_1985( .carry(c_116_1985), .sum(s_116_1985), .in3(c_115_1977), .in2(s_116_1983), .in1(c_115_1978) );
  Fadder_ A_116_1986( .carry(c[116]), .sum(s[116]), .in3(s_116_1984), .in2(c_115_1979), .in1(s_116_1985) );

  // ***** Bit 117 ***** //
  Fadder_ A_117_1987( .carry(c_117_1987), .sum(s_117_1987), .in3(P_31[55]), .in2(P_30[57]), .in1(P_29[59]) );
  Fadder_ A_117_1988( .carry(c_117_1988), .sum(s_117_1988), .in3(P_28[61]), .in2(P_27[63]), .in1(P_26[65]) );
  Fadder_ A_117_1989( .carry(c_117_1989), .sum(s_117_1989), .in3(c_116_1981), .in2(c_116_1982), .in1(s_117_1988) );
  Fadder_ A_117_1990( .carry(c_117_1990), .sum(s_117_1990), .in3(s_117_1987), .in2(c_116_1983), .in1(c_116_1984) );
  Fadder_ A_117_1991( .carry(c[117]), .sum(s[117]), .in3(s_117_1989), .in2(c_116_1985), .in1(s_117_1990) );

  // ***** Bit 118 ***** //
  Hadder_ A_118_1992( .carry(c_118_1992), .sum(s_118_1992), .in2(sign_), .in1(P_31[56]) );
  Fadder_ A_118_1993( .carry(c_118_1993), .sum(s_118_1993), .in3(P_30[58]), .in2(P_29[60]), .in1(P_28[62]) );
  Fadder_ A_118_1994( .carry(c_118_1994), .sum(s_118_1994), .in3(P_27[64]), .in2(c_117_1988), .in1(c_117_1987) );
  Fadder_ A_118_1995( .carry(c_118_1995), .sum(s_118_1995), .in3(s_118_1992), .in2(s_118_1993), .in1(c_117_1989) );
  Fadder_ A_118_1996( .carry(c[118]), .sum(s[118]), .in3(s_118_1994), .in2(c_117_1990), .in1(s_118_1995) );

  // ***** Bit 119 ***** //
  Fadder_ A_119_1997( .carry(c_119_1997), .sum(s_119_1997), .in3(P_31[57]), .in2(P_30[59]), .in1(P_29[61]) );
  Fadder_ A_119_1998( .carry(c_119_1998), .sum(s_119_1998), .in3(P_28[63]), .in2(P_27[65]), .in1(c_118_1992) );
  Fadder_ A_119_1999( .carry(c_119_1999), .sum(s_119_1999), .in3(c_118_1993), .in2(s_119_1997), .in1(s_119_1998) );
  Fadder_ A_119_2000( .carry(c[119]), .sum(s[119]), .in3(c_118_1994), .in2(s_119_1999), .in1(c_118_1995) );

  // ***** Bit 120 ***** //
  Hadder_ A_120_2001( .carry(c_120_2001), .sum(s_120_2001), .in2(sign_), .in1(P_31[58]) );
  Fadder_ A_120_2002( .carry(c_120_2002), .sum(s_120_2002), .in3(P_30[60]), .in2(P_29[62]), .in1(P_28[64]) );
  Fadder_ A_120_2003( .carry(c_120_2003), .sum(s_120_2003), .in3(c_119_1997), .in2(s_120_2001), .in1(s_120_2002) );
  Fadder_ A_120_2004( .carry(c[120]), .sum(s[120]), .in3(c_119_1998), .in2(s_120_2003), .in1(c_119_1999) );

  // ***** Bit 121 ***** //
  Fadder_ A_121_2005( .carry(c_121_2005), .sum(s_121_2005), .in3(P_31[59]), .in2(P_30[61]), .in1(P_29[63]) );
  Fadder_ A_121_2006( .carry(c_121_2006), .sum(s_121_2006), .in3(P_28[65]), .in2(c_120_2001), .in1(c_120_2002) );
  Fadder_ A_121_2007( .carry(c[121]), .sum(s[121]), .in3(s_121_2005), .in2(c_120_2003), .in1(s_121_2006) );

  // ***** Bit 122 ***** //
  Hadder_ A_122_2008( .carry(c_122_2008), .sum(s_122_2008), .in2(sign_), .in1(P_31[60]) );
  Fadder_ A_122_2009( .carry(c_122_2009), .sum(s_122_2009), .in3(P_30[62]), .in2(P_29[64]), .in1(c_121_2005) );
  Fadder_ A_122_2010( .carry(c[122]), .sum(s[122]), .in3(s_122_2008), .in2(c_121_2006), .in1(s_122_2009) );

  // ***** Bit 123 ***** //
  Fadder_ A_123_2011( .carry(c_123_2011), .sum(s_123_2011), .in3(P_31[61]), .in2(P_30[63]), .in1(P_29[65]) );
  Fadder_ A_123_2012( .carry(c[123]), .sum(s[123]), .in3(c_122_2008), .in2(s_123_2011), .in1(c_122_2009) );

  // ***** Bit 124 ***** //
  Hadder_ A_124_2013( .carry(c_124_2013), .sum(s_124_2013), .in2(sign_), .in1(P_31[62]) );
  Fadder_ A_124_2014( .carry(c[124]), .sum(s[124]), .in3(P_30[64]), .in2(c_123_2011), .in1(s_124_2013) );

  // ***** Bit 125 ***** //
  Fadder_ A_125_2015( .carry(c[125]), .sum(s[125]), .in3(P_31[63]), .in2(P_30[65]), .in1(c_124_2013) );

  // ***** Bit 126 ***** //
  Hadder_ A_126_2016( .carry(c[126]), .sum(s[126]), .in2(sign_), .in1(P_31[64]) );

  // ***** Bit 127 ***** //
  assign s[127] = P_31[65] ;

endmodule

module add_csa140(
  add_sub,
  in_sum,
  in_carry,
  product,
  out_sum,
  out_carry);

  input add_sub;
  input [139:0] in_sum;
  input [138:0] in_carry;
  input [139:0] product;
  output [139:0] out_sum, out_carry;

  wire inc;
  wire [139:0] comp_sum;
  wire [138:0] comp_carry;

  assign inc = (add_sub==1'b1)? 1'b0 : 1'b1;
  assign comp_sum = (add_sub==1'b1)? in_sum : (~in_sum);
  assign comp_carry = (add_sub==1'b1)? in_carry : (~in_carry);

  Fadder_ u0( .in3(comp_sum[0]), .in2(product[0]), .in1(inc), .sum(out_sum[0]), .carry(out_carry[0]) );
  Fadder_ u1( .in3(comp_sum[1]), .in2(comp_carry[0]), .in1(product[1]), .sum(out_sum[1]), .carry(out_carry[1]) );
  Fadder_ u2( .in3(comp_sum[2]), .in2(comp_carry[1]), .in1(product[2]), .sum(out_sum[2]), .carry(out_carry[2]) );
  Fadder_ u3( .in3(comp_sum[3]), .in2(comp_carry[2]), .in1(product[3]), .sum(out_sum[3]), .carry(out_carry[3]) );
  Fadder_ u4( .in3(comp_sum[4]), .in2(comp_carry[3]), .in1(product[4]), .sum(out_sum[4]), .carry(out_carry[4]) );
  Fadder_ u5( .in3(comp_sum[5]), .in2(comp_carry[4]), .in1(product[5]), .sum(out_sum[5]), .carry(out_carry[5]) );
  Fadder_ u6( .in3(comp_sum[6]), .in2(comp_carry[5]), .in1(product[6]), .sum(out_sum[6]), .carry(out_carry[6]) );
  Fadder_ u7( .in3(comp_sum[7]), .in2(comp_carry[6]), .in1(product[7]), .sum(out_sum[7]), .carry(out_carry[7]) );
  Fadder_ u8( .in3(comp_sum[8]), .in2(comp_carry[7]), .in1(product[8]), .sum(out_sum[8]), .carry(out_carry[8]) );
  Fadder_ u9( .in3(comp_sum[9]), .in2(comp_carry[8]), .in1(product[9]), .sum(out_sum[9]), .carry(out_carry[9]) );
  Fadder_ u10( .in3(comp_sum[10]), .in2(comp_carry[9]), .in1(product[10]), .sum(out_sum[10]), .carry(out_carry[10]) );
  Fadder_ u11( .in3(comp_sum[11]), .in2(comp_carry[10]), .in1(product[11]), .sum(out_sum[11]), .carry(out_carry[11]) );
  Fadder_ u12( .in3(comp_sum[12]), .in2(comp_carry[11]), .in1(product[12]), .sum(out_sum[12]), .carry(out_carry[12]) );
  Fadder_ u13( .in3(comp_sum[13]), .in2(comp_carry[12]), .in1(product[13]), .sum(out_sum[13]), .carry(out_carry[13]) );
  Fadder_ u14( .in3(comp_sum[14]), .in2(comp_carry[13]), .in1(product[14]), .sum(out_sum[14]), .carry(out_carry[14]) );
  Fadder_ u15( .in3(comp_sum[15]), .in2(comp_carry[14]), .in1(product[15]), .sum(out_sum[15]), .carry(out_carry[15]) );
  Fadder_ u16( .in3(comp_sum[16]), .in2(comp_carry[15]), .in1(product[16]), .sum(out_sum[16]), .carry(out_carry[16]) );
  Fadder_ u17( .in3(comp_sum[17]), .in2(comp_carry[16]), .in1(product[17]), .sum(out_sum[17]), .carry(out_carry[17]) );
  Fadder_ u18( .in3(comp_sum[18]), .in2(comp_carry[17]), .in1(product[18]), .sum(out_sum[18]), .carry(out_carry[18]) );
  Fadder_ u19( .in3(comp_sum[19]), .in2(comp_carry[18]), .in1(product[19]), .sum(out_sum[19]), .carry(out_carry[19]) );
  Fadder_ u20( .in3(comp_sum[20]), .in2(comp_carry[19]), .in1(product[20]), .sum(out_sum[20]), .carry(out_carry[20]) );
  Fadder_ u21( .in3(comp_sum[21]), .in2(comp_carry[20]), .in1(product[21]), .sum(out_sum[21]), .carry(out_carry[21]) );
  Fadder_ u22( .in3(comp_sum[22]), .in2(comp_carry[21]), .in1(product[22]), .sum(out_sum[22]), .carry(out_carry[22]) );
  Fadder_ u23( .in3(comp_sum[23]), .in2(comp_carry[22]), .in1(product[23]), .sum(out_sum[23]), .carry(out_carry[23]) );
  Fadder_ u24( .in3(comp_sum[24]), .in2(comp_carry[23]), .in1(product[24]), .sum(out_sum[24]), .carry(out_carry[24]) );
  Fadder_ u25( .in3(comp_sum[25]), .in2(comp_carry[24]), .in1(product[25]), .sum(out_sum[25]), .carry(out_carry[25]) );
  Fadder_ u26( .in3(comp_sum[26]), .in2(comp_carry[25]), .in1(product[26]), .sum(out_sum[26]), .carry(out_carry[26]) );
  Fadder_ u27( .in3(comp_sum[27]), .in2(comp_carry[26]), .in1(product[27]), .sum(out_sum[27]), .carry(out_carry[27]) );
  Fadder_ u28( .in3(comp_sum[28]), .in2(comp_carry[27]), .in1(product[28]), .sum(out_sum[28]), .carry(out_carry[28]) );
  Fadder_ u29( .in3(comp_sum[29]), .in2(comp_carry[28]), .in1(product[29]), .sum(out_sum[29]), .carry(out_carry[29]) );
  Fadder_ u30( .in3(comp_sum[30]), .in2(comp_carry[29]), .in1(product[30]), .sum(out_sum[30]), .carry(out_carry[30]) );
  Fadder_ u31( .in3(comp_sum[31]), .in2(comp_carry[30]), .in1(product[31]), .sum(out_sum[31]), .carry(out_carry[31]) );
  Fadder_ u32( .in3(comp_sum[32]), .in2(comp_carry[31]), .in1(product[32]), .sum(out_sum[32]), .carry(out_carry[32]) );
  Fadder_ u33( .in3(comp_sum[33]), .in2(comp_carry[32]), .in1(product[33]), .sum(out_sum[33]), .carry(out_carry[33]) );
  Fadder_ u34( .in3(comp_sum[34]), .in2(comp_carry[33]), .in1(product[34]), .sum(out_sum[34]), .carry(out_carry[34]) );
  Fadder_ u35( .in3(comp_sum[35]), .in2(comp_carry[34]), .in1(product[35]), .sum(out_sum[35]), .carry(out_carry[35]) );
  Fadder_ u36( .in3(comp_sum[36]), .in2(comp_carry[35]), .in1(product[36]), .sum(out_sum[36]), .carry(out_carry[36]) );
  Fadder_ u37( .in3(comp_sum[37]), .in2(comp_carry[36]), .in1(product[37]), .sum(out_sum[37]), .carry(out_carry[37]) );
  Fadder_ u38( .in3(comp_sum[38]), .in2(comp_carry[37]), .in1(product[38]), .sum(out_sum[38]), .carry(out_carry[38]) );
  Fadder_ u39( .in3(comp_sum[39]), .in2(comp_carry[38]), .in1(product[39]), .sum(out_sum[39]), .carry(out_carry[39]) );
  Fadder_ u40( .in3(comp_sum[40]), .in2(comp_carry[39]), .in1(product[40]), .sum(out_sum[40]), .carry(out_carry[40]) );
  Fadder_ u41( .in3(comp_sum[41]), .in2(comp_carry[40]), .in1(product[41]), .sum(out_sum[41]), .carry(out_carry[41]) );
  Fadder_ u42( .in3(comp_sum[42]), .in2(comp_carry[41]), .in1(product[42]), .sum(out_sum[42]), .carry(out_carry[42]) );
  Fadder_ u43( .in3(comp_sum[43]), .in2(comp_carry[42]), .in1(product[43]), .sum(out_sum[43]), .carry(out_carry[43]) );
  Fadder_ u44( .in3(comp_sum[44]), .in2(comp_carry[43]), .in1(product[44]), .sum(out_sum[44]), .carry(out_carry[44]) );
  Fadder_ u45( .in3(comp_sum[45]), .in2(comp_carry[44]), .in1(product[45]), .sum(out_sum[45]), .carry(out_carry[45]) );
  Fadder_ u46( .in3(comp_sum[46]), .in2(comp_carry[45]), .in1(product[46]), .sum(out_sum[46]), .carry(out_carry[46]) );
  Fadder_ u47( .in3(comp_sum[47]), .in2(comp_carry[46]), .in1(product[47]), .sum(out_sum[47]), .carry(out_carry[47]) );
  Fadder_ u48( .in3(comp_sum[48]), .in2(comp_carry[47]), .in1(product[48]), .sum(out_sum[48]), .carry(out_carry[48]) );
  Fadder_ u49( .in3(comp_sum[49]), .in2(comp_carry[48]), .in1(product[49]), .sum(out_sum[49]), .carry(out_carry[49]) );
  Fadder_ u50( .in3(comp_sum[50]), .in2(comp_carry[49]), .in1(product[50]), .sum(out_sum[50]), .carry(out_carry[50]) );
  Fadder_ u51( .in3(comp_sum[51]), .in2(comp_carry[50]), .in1(product[51]), .sum(out_sum[51]), .carry(out_carry[51]) );
  Fadder_ u52( .in3(comp_sum[52]), .in2(comp_carry[51]), .in1(product[52]), .sum(out_sum[52]), .carry(out_carry[52]) );
  Fadder_ u53( .in3(comp_sum[53]), .in2(comp_carry[52]), .in1(product[53]), .sum(out_sum[53]), .carry(out_carry[53]) );
  Fadder_ u54( .in3(comp_sum[54]), .in2(comp_carry[53]), .in1(product[54]), .sum(out_sum[54]), .carry(out_carry[54]) );
  Fadder_ u55( .in3(comp_sum[55]), .in2(comp_carry[54]), .in1(product[55]), .sum(out_sum[55]), .carry(out_carry[55]) );
  Fadder_ u56( .in3(comp_sum[56]), .in2(comp_carry[55]), .in1(product[56]), .sum(out_sum[56]), .carry(out_carry[56]) );
  Fadder_ u57( .in3(comp_sum[57]), .in2(comp_carry[56]), .in1(product[57]), .sum(out_sum[57]), .carry(out_carry[57]) );
  Fadder_ u58( .in3(comp_sum[58]), .in2(comp_carry[57]), .in1(product[58]), .sum(out_sum[58]), .carry(out_carry[58]) );
  Fadder_ u59( .in3(comp_sum[59]), .in2(comp_carry[58]), .in1(product[59]), .sum(out_sum[59]), .carry(out_carry[59]) );
  Fadder_ u60( .in3(comp_sum[60]), .in2(comp_carry[59]), .in1(product[60]), .sum(out_sum[60]), .carry(out_carry[60]) );
  Fadder_ u61( .in3(comp_sum[61]), .in2(comp_carry[60]), .in1(product[61]), .sum(out_sum[61]), .carry(out_carry[61]) );
  Fadder_ u62( .in3(comp_sum[62]), .in2(comp_carry[61]), .in1(product[62]), .sum(out_sum[62]), .carry(out_carry[62]) );
  Fadder_ u63( .in3(comp_sum[63]), .in2(comp_carry[62]), .in1(product[63]), .sum(out_sum[63]), .carry(out_carry[63]) );
  Fadder_ u64( .in3(comp_sum[64]), .in2(comp_carry[63]), .in1(product[64]), .sum(out_sum[64]), .carry(out_carry[64]) );
  Fadder_ u65( .in3(comp_sum[65]), .in2(comp_carry[64]), .in1(product[65]), .sum(out_sum[65]), .carry(out_carry[65]) );
  Fadder_ u66( .in3(comp_sum[66]), .in2(comp_carry[65]), .in1(product[66]), .sum(out_sum[66]), .carry(out_carry[66]) );
  Fadder_ u67( .in3(comp_sum[67]), .in2(comp_carry[66]), .in1(product[67]), .sum(out_sum[67]), .carry(out_carry[67]) );
  Fadder_ u68( .in3(comp_sum[68]), .in2(comp_carry[67]), .in1(product[68]), .sum(out_sum[68]), .carry(out_carry[68]) );
  Fadder_ u69( .in3(comp_sum[69]), .in2(comp_carry[68]), .in1(product[69]), .sum(out_sum[69]), .carry(out_carry[69]) );
  Fadder_ u70( .in3(comp_sum[70]), .in2(comp_carry[69]), .in1(product[70]), .sum(out_sum[70]), .carry(out_carry[70]) );
  Fadder_ u71( .in3(comp_sum[71]), .in2(comp_carry[70]), .in1(product[71]), .sum(out_sum[71]), .carry(out_carry[71]) );
  Fadder_ u72( .in3(comp_sum[72]), .in2(comp_carry[71]), .in1(product[72]), .sum(out_sum[72]), .carry(out_carry[72]) );
  Fadder_ u73( .in3(comp_sum[73]), .in2(comp_carry[72]), .in1(product[73]), .sum(out_sum[73]), .carry(out_carry[73]) );
  Fadder_ u74( .in3(comp_sum[74]), .in2(comp_carry[73]), .in1(product[74]), .sum(out_sum[74]), .carry(out_carry[74]) );
  Fadder_ u75( .in3(comp_sum[75]), .in2(comp_carry[74]), .in1(product[75]), .sum(out_sum[75]), .carry(out_carry[75]) );
  Fadder_ u76( .in3(comp_sum[76]), .in2(comp_carry[75]), .in1(product[76]), .sum(out_sum[76]), .carry(out_carry[76]) );
  Fadder_ u77( .in3(comp_sum[77]), .in2(comp_carry[76]), .in1(product[77]), .sum(out_sum[77]), .carry(out_carry[77]) );
  Fadder_ u78( .in3(comp_sum[78]), .in2(comp_carry[77]), .in1(product[78]), .sum(out_sum[78]), .carry(out_carry[78]) );
  Fadder_ u79( .in3(comp_sum[79]), .in2(comp_carry[78]), .in1(product[79]), .sum(out_sum[79]), .carry(out_carry[79]) );
  Fadder_ u80( .in3(comp_sum[80]), .in2(comp_carry[79]), .in1(product[80]), .sum(out_sum[80]), .carry(out_carry[80]) );
  Fadder_ u81( .in3(comp_sum[81]), .in2(comp_carry[80]), .in1(product[81]), .sum(out_sum[81]), .carry(out_carry[81]) );
  Fadder_ u82( .in3(comp_sum[82]), .in2(comp_carry[81]), .in1(product[82]), .sum(out_sum[82]), .carry(out_carry[82]) );
  Fadder_ u83( .in3(comp_sum[83]), .in2(comp_carry[82]), .in1(product[83]), .sum(out_sum[83]), .carry(out_carry[83]) );
  Fadder_ u84( .in3(comp_sum[84]), .in2(comp_carry[83]), .in1(product[84]), .sum(out_sum[84]), .carry(out_carry[84]) );
  Fadder_ u85( .in3(comp_sum[85]), .in2(comp_carry[84]), .in1(product[85]), .sum(out_sum[85]), .carry(out_carry[85]) );
  Fadder_ u86( .in3(comp_sum[86]), .in2(comp_carry[85]), .in1(product[86]), .sum(out_sum[86]), .carry(out_carry[86]) );
  Fadder_ u87( .in3(comp_sum[87]), .in2(comp_carry[86]), .in1(product[87]), .sum(out_sum[87]), .carry(out_carry[87]) );
  Fadder_ u88( .in3(comp_sum[88]), .in2(comp_carry[87]), .in1(product[88]), .sum(out_sum[88]), .carry(out_carry[88]) );
  Fadder_ u89( .in3(comp_sum[89]), .in2(comp_carry[88]), .in1(product[89]), .sum(out_sum[89]), .carry(out_carry[89]) );
  Fadder_ u90( .in3(comp_sum[90]), .in2(comp_carry[89]), .in1(product[90]), .sum(out_sum[90]), .carry(out_carry[90]) );
  Fadder_ u91( .in3(comp_sum[91]), .in2(comp_carry[90]), .in1(product[91]), .sum(out_sum[91]), .carry(out_carry[91]) );
  Fadder_ u92( .in3(comp_sum[92]), .in2(comp_carry[91]), .in1(product[92]), .sum(out_sum[92]), .carry(out_carry[92]) );
  Fadder_ u93( .in3(comp_sum[93]), .in2(comp_carry[92]), .in1(product[93]), .sum(out_sum[93]), .carry(out_carry[93]) );
  Fadder_ u94( .in3(comp_sum[94]), .in2(comp_carry[93]), .in1(product[94]), .sum(out_sum[94]), .carry(out_carry[94]) );
  Fadder_ u95( .in3(comp_sum[95]), .in2(comp_carry[94]), .in1(product[95]), .sum(out_sum[95]), .carry(out_carry[95]) );
  Fadder_ u96( .in3(comp_sum[96]), .in2(comp_carry[95]), .in1(product[96]), .sum(out_sum[96]), .carry(out_carry[96]) );
  Fadder_ u97( .in3(comp_sum[97]), .in2(comp_carry[96]), .in1(product[97]), .sum(out_sum[97]), .carry(out_carry[97]) );
  Fadder_ u98( .in3(comp_sum[98]), .in2(comp_carry[97]), .in1(product[98]), .sum(out_sum[98]), .carry(out_carry[98]) );
  Fadder_ u99( .in3(comp_sum[99]), .in2(comp_carry[98]), .in1(product[99]), .sum(out_sum[99]), .carry(out_carry[99]) );
  Fadder_ u100( .in3(comp_sum[100]), .in2(comp_carry[99]), .in1(product[100]), .sum(out_sum[100]), .carry(out_carry[100]) );
  Fadder_ u101( .in3(comp_sum[101]), .in2(comp_carry[100]), .in1(product[101]), .sum(out_sum[101]), .carry(out_carry[101]) );
  Fadder_ u102( .in3(comp_sum[102]), .in2(comp_carry[101]), .in1(product[102]), .sum(out_sum[102]), .carry(out_carry[102]) );
  Fadder_ u103( .in3(comp_sum[103]), .in2(comp_carry[102]), .in1(product[103]), .sum(out_sum[103]), .carry(out_carry[103]) );
  Fadder_ u104( .in3(comp_sum[104]), .in2(comp_carry[103]), .in1(product[104]), .sum(out_sum[104]), .carry(out_carry[104]) );
  Fadder_ u105( .in3(comp_sum[105]), .in2(comp_carry[104]), .in1(product[105]), .sum(out_sum[105]), .carry(out_carry[105]) );
  Fadder_ u106( .in3(comp_sum[106]), .in2(comp_carry[105]), .in1(product[106]), .sum(out_sum[106]), .carry(out_carry[106]) );
  Fadder_ u107( .in3(comp_sum[107]), .in2(comp_carry[106]), .in1(product[107]), .sum(out_sum[107]), .carry(out_carry[107]) );
  Fadder_ u108( .in3(comp_sum[108]), .in2(comp_carry[107]), .in1(product[108]), .sum(out_sum[108]), .carry(out_carry[108]) );
  Fadder_ u109( .in3(comp_sum[109]), .in2(comp_carry[108]), .in1(product[109]), .sum(out_sum[109]), .carry(out_carry[109]) );
  Fadder_ u110( .in3(comp_sum[110]), .in2(comp_carry[109]), .in1(product[110]), .sum(out_sum[110]), .carry(out_carry[110]) );
  Fadder_ u111( .in3(comp_sum[111]), .in2(comp_carry[110]), .in1(product[111]), .sum(out_sum[111]), .carry(out_carry[111]) );
  Fadder_ u112( .in3(comp_sum[112]), .in2(comp_carry[111]), .in1(product[112]), .sum(out_sum[112]), .carry(out_carry[112]) );
  Fadder_ u113( .in3(comp_sum[113]), .in2(comp_carry[112]), .in1(product[113]), .sum(out_sum[113]), .carry(out_carry[113]) );
  Fadder_ u114( .in3(comp_sum[114]), .in2(comp_carry[113]), .in1(product[114]), .sum(out_sum[114]), .carry(out_carry[114]) );
  Fadder_ u115( .in3(comp_sum[115]), .in2(comp_carry[114]), .in1(product[115]), .sum(out_sum[115]), .carry(out_carry[115]) );
  Fadder_ u116( .in3(comp_sum[116]), .in2(comp_carry[115]), .in1(product[116]), .sum(out_sum[116]), .carry(out_carry[116]) );
  Fadder_ u117( .in3(comp_sum[117]), .in2(comp_carry[116]), .in1(product[117]), .sum(out_sum[117]), .carry(out_carry[117]) );
  Fadder_ u118( .in3(comp_sum[118]), .in2(comp_carry[117]), .in1(product[118]), .sum(out_sum[118]), .carry(out_carry[118]) );
  Fadder_ u119( .in3(comp_sum[119]), .in2(comp_carry[118]), .in1(product[119]), .sum(out_sum[119]), .carry(out_carry[119]) );
  Fadder_ u120( .in3(comp_sum[120]), .in2(comp_carry[119]), .in1(product[120]), .sum(out_sum[120]), .carry(out_carry[120]) );
  Fadder_ u121( .in3(comp_sum[121]), .in2(comp_carry[120]), .in1(product[121]), .sum(out_sum[121]), .carry(out_carry[121]) );
  Fadder_ u122( .in3(comp_sum[122]), .in2(comp_carry[121]), .in1(product[122]), .sum(out_sum[122]), .carry(out_carry[122]) );
  Fadder_ u123( .in3(comp_sum[123]), .in2(comp_carry[122]), .in1(product[123]), .sum(out_sum[123]), .carry(out_carry[123]) );
  Fadder_ u124( .in3(comp_sum[124]), .in2(comp_carry[123]), .in1(product[124]), .sum(out_sum[124]), .carry(out_carry[124]) );
  Fadder_ u125( .in3(comp_sum[125]), .in2(comp_carry[124]), .in1(product[125]), .sum(out_sum[125]), .carry(out_carry[125]) );
  Fadder_ u126( .in3(comp_sum[126]), .in2(comp_carry[125]), .in1(product[126]), .sum(out_sum[126]), .carry(out_carry[126]) );
  Fadder_ u127( .in3(comp_sum[127]), .in2(comp_carry[126]), .in1(product[127]), .sum(out_sum[127]), .carry(out_carry[127]) );
  Fadder_ u128( .in3(comp_sum[128]), .in2(comp_carry[127]), .in1(product[128]), .sum(out_sum[128]), .carry(out_carry[128]) );
  Fadder_ u129( .in3(comp_sum[129]), .in2(comp_carry[128]), .in1(product[129]), .sum(out_sum[129]), .carry(out_carry[129]) );
  Fadder_ u130( .in3(comp_sum[130]), .in2(comp_carry[129]), .in1(product[130]), .sum(out_sum[130]), .carry(out_carry[130]) );
  Fadder_ u131( .in3(comp_sum[131]), .in2(comp_carry[130]), .in1(product[131]), .sum(out_sum[131]), .carry(out_carry[131]) );
  Fadder_ u132( .in3(comp_sum[132]), .in2(comp_carry[131]), .in1(product[132]), .sum(out_sum[132]), .carry(out_carry[132]) );
  Fadder_ u133( .in3(comp_sum[133]), .in2(comp_carry[132]), .in1(product[133]), .sum(out_sum[133]), .carry(out_carry[133]) );
  Fadder_ u134( .in3(comp_sum[134]), .in2(comp_carry[133]), .in1(product[134]), .sum(out_sum[134]), .carry(out_carry[134]) );
  Fadder_ u135( .in3(comp_sum[135]), .in2(comp_carry[134]), .in1(product[135]), .sum(out_sum[135]), .carry(out_carry[135]) );
  Fadder_ u136( .in3(comp_sum[136]), .in2(comp_carry[135]), .in1(product[136]), .sum(out_sum[136]), .carry(out_carry[136]) );
  Fadder_ u137( .in3(comp_sum[137]), .in2(comp_carry[136]), .in1(product[137]), .sum(out_sum[137]), .carry(out_carry[137]) );
  Fadder_ u138( .in3(comp_sum[138]), .in2(comp_carry[137]), .in1(product[138]), .sum(out_sum[138]), .carry(out_carry[138]) );
  Fadder_ u139( .in3(comp_sum[139]), .in2(comp_carry[138]), .in1(product[139]), .sum(out_sum[139]), .carry(out_carry[139]) );

endmodule

module DW01_add2 (A,B,CI,SUM,CO);

  parameter width=71;

  output [width-1 : 0] SUM;
  output CO;
  input [width-1 : 0] A,B;
  input CI;

  wire [width-1 : 0] SUM;
  reg [width-2 : 0] sum_temp;
  reg CO;

  assign SUM = {CO, sum_temp};

always @(A or B or CI)
  begin
    {CO, sum_temp} = A+B+CI;
  end
endmodule

module DW01_add1 (A,B,CI,SUM,CO);

  parameter width=70;

  output [width-1 : 0] SUM;
  output CO;
  input [width-1 : 0] A,B;
  input CI;

  wire [width-1 : 0] SUM;
  reg [width-2 : 0] sum_temp;
  reg CO;
  reg c_out;

	assign SUM = {CO, sum_temp};

always @(A or B or CI)
  begin
    {CO, sum_temp} = A+B+CI;
//	sum_out = A + B;
//    plus(sum_out,c_out,A,B,CI);
//    SUM = sum_out;
//    CO =  c_out;
  end

/*
  task plus;
    output  [width-1 : 0] sumout;
    output CO;
    input [width-1 : 0] A,B;
    input CI;
    reg [width-1 : 0] sumout,SUM;
    reg CO;
    reg carry;
    reg [width-1 : 0] A,B;
    integer i;

    begin
      carry = CI;
      for (i = 0; i <= width-1; i = i + 1) begin
        sumout[i] = A[i] ^ B[i] ^ carry;
        carry = (A[i] & B[i]) | (A[i] & carry) | (carry & B[i]);
      end
      SUM = sumout;
      CO = carry;
    end
  endtask
*/
endmodule

module Adder141(
  a,
  b,
  cin,
  sum,
  cout);

  input [140:0]a, b;
  input cin;
  output [140:0]sum;
  output cout;

  wire [69:0] temp1, result1;
  wire [70:0] temp2_1, temp2_2, result2;
  wire co1, co2_1, co2_2;

  assign result1= temp1;
  assign result2= (co1==1'b0) ? temp2_1 : temp2_2;
  assign sum={result2,result1};
  assign cout=(co1==1'b0) ? co2_1 : co2_2;

  DW01_add1  u1_1(.A(a[69:0]), .B(b[69:0]), .CI(cin), .SUM(temp1), .CO(co1));
  DW01_add2  u2_1(.A(a[140:70]), .B(b[140:70]), .CI(1'b0), .SUM(temp2_1), .CO(co2_1));
  DW01_add2  u2_2(.A(a[140:70]), .B(b[140:70]), .CI(1'b1), .SUM(temp2_2), .CO(co2_2));

endmodule

module cla_csa140(
  sum,
  carry,
  add_sub,
  result,
  overflow);

  input [139:0] sum;
  input [139:0] carry;
  input add_sub;
  output [139:0] result;
  output overflow;

  reg [139:0] result;
  reg overflow;
  wire [140:0] temp;
  wire inc1, inc2;

  assign inc1=(add_sub==1'b1)? 1'b0 : 1'b1;
  assign inc2=(add_sub==1'b1)? 1'b0 : 1'b1;

  Adder141 U(.a({sum[139],sum}), .b({carry,inc1}), .cin(inc2), .sum(temp));

  always @( temp )
    begin
      result = temp[139:0];
      if (temp[140]^temp[139]==1'b1)
        overflow = 1'b1;
      else
        overflow = 1'b0;
    end

endmodule


module mac2(
  clk,
  reset,
  stall,
  add_sub,
  mode,
  mulcand,
  mulier,
  init_value,
  cnt_overflow,
  answer,
  overflow);

  input clk;
  input reset;
  input stall;
  input add_sub;
  input mode;
  input [139:0] init_value;
  input [63:0] mulcand;
  input [63:0] mulier;
  input cnt_overflow;
  output [139:0] answer;
  output overflow;

  reg [63:0] in1;
  reg [63:0] in2;
  wire [127:0] wire_s;
  wire [126:0] wire_c;
  reg [127:0] temp_s;
  reg [126:0] temp_c;
  wire [139:0] operand_answer;
  wire [139:0] operand_s;
  wire [138:0] operand_c;
  wire [139:0] final_sum;
  wire [139:0] final_carry;
  wire [139:0] wire_answer;
  reg [139:0] answer;
  wire [139:0] final_answer;
  wire wire_overflow;
  reg overflow;

  assign operand_answer = mode==1'b0 ? answer : 'b0; 
  assign final_answer=((wire_overflow&cnt_overflow)==1'b1) ? 140'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111 : wire_answer;
  assign operand_s ={ temp_s[127],temp_s[127],temp_s[127],temp_s[127],temp_s[127],temp_s[127],temp_s[127],temp_s[127],temp_s[127],temp_s[127],temp_s[127],temp_s[127],temp_s };
  assign operand_c ={ temp_c[126],temp_c[126],temp_c[126],temp_c[126],temp_c[126],temp_c[126],temp_c[126],temp_c[126],temp_c[126],temp_c[126],temp_c[126],temp_c[126],temp_c };

  mult_ u1(.a(in1), .b(in2), .s(wire_s), .c(wire_c));

  add_csa140 u2( .add_sub(add_sub), .in_sum(operand_s), .in_carry(operand_c), .product(operand_answer), .out_sum(final_sum), .out_carry(final_carry) );

  cla_csa140 u3( .add_sub(add_sub), .sum(final_sum), .carry(final_carry), .result(wire_answer), .overflow(wire_overflow) );

  always @(posedge clk)
    begin
    if( reset==1'b1 )
      begin
      in1<='b0;
      in2<='b0;
      temp_s<='b0;
      temp_c<='b0;
      answer<=init_value;
      overflow<='b0;
      end
    else
      begin
      if (stall==1'b0)
        begin
        in1<=mulcand;
        in2<=mulier;
        temp_s<=wire_s;
        temp_c<=wire_c;
        overflow<=wire_overflow;
        answer<=final_answer;
        end
      end
    end

endmodule
