`define BINARY_OP(out,a,b) xnor(out, a, b);
`include "../.generic/wire_test.v"