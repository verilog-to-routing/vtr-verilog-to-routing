`define BINARY_OP(out,a,b) xnor(out, a, b);
`include "wire_test.v"