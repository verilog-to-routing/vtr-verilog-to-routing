module test4(input [2:0] a, output [2:0] b);
    wire [2:0] c;
    assign c = a;
    assign b = c;
endmodule