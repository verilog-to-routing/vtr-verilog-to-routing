module test2(input [2:0] a, output [2:0] b);
    assign b = a;
endmodule