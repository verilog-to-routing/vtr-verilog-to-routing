/*

Copyright (c) 2020 Alex Forencich

Permission is hereby granted, free of charge, to any person obtaining a copy
of this software and associated documentation files (the "Software"), to deal
in the Software without restriction, including without limitation the rights
to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
copies of the Software, and to permit persons to whom the Software is
furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in
all copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY
FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
THE SOFTWARE.

*/

// Language: Verilog 2001

`resetall
`timescale 1ns / 1ps
`default_nettype none

/*
 * AXI4 lite 1x24 interconnect (wrapper)
 */
module axil_interconnect_wrap_1x24 #
(
    parameter DATA_WIDTH = 32,
    parameter ADDR_WIDTH = 16,
    parameter STRB_WIDTH = (DATA_WIDTH/8),
    parameter M_REGIONS = 1,
    parameter M00_BASE_ADDR = 0,
    parameter M00_ADDR_WIDTH = {M_REGIONS{32'd24}},
    parameter M00_CONNECT_READ = 1'b1,
    parameter M00_CONNECT_WRITE = 1'b1,
    parameter M00_SECURE = 1'b0,
    parameter M01_BASE_ADDR = 0,
    parameter M01_ADDR_WIDTH = {M_REGIONS{32'd24}},
    parameter M01_CONNECT_READ = 1'b1,
    parameter M01_CONNECT_WRITE = 1'b1,
    parameter M01_SECURE = 1'b0,
    parameter M02_BASE_ADDR = 0,
    parameter M02_ADDR_WIDTH = {M_REGIONS{32'd24}},
    parameter M02_CONNECT_READ = 1'b1,
    parameter M02_CONNECT_WRITE = 1'b1,
    parameter M02_SECURE = 1'b0,
    parameter M03_BASE_ADDR = 0,
    parameter M03_ADDR_WIDTH = {M_REGIONS{32'd24}},
    parameter M03_CONNECT_READ = 1'b1,
    parameter M03_CONNECT_WRITE = 1'b1,
    parameter M03_SECURE = 1'b0,
    parameter M04_BASE_ADDR = 0,
    parameter M04_ADDR_WIDTH = {M_REGIONS{32'd24}},
    parameter M04_CONNECT_READ = 1'b1,
    parameter M04_CONNECT_WRITE = 1'b1,
    parameter M04_SECURE = 1'b0,
    parameter M05_BASE_ADDR = 0,
    parameter M05_ADDR_WIDTH = {M_REGIONS{32'd24}},
    parameter M05_CONNECT_READ = 1'b1,
    parameter M05_CONNECT_WRITE = 1'b1,
    parameter M05_SECURE = 1'b0,
    parameter M06_BASE_ADDR = 0,
    parameter M06_ADDR_WIDTH = {M_REGIONS{32'd24}},
    parameter M06_CONNECT_READ = 1'b1,
    parameter M06_CONNECT_WRITE = 1'b1,
    parameter M06_SECURE = 1'b0,
    parameter M07_BASE_ADDR = 0,
    parameter M07_ADDR_WIDTH = {M_REGIONS{32'd24}},
    parameter M07_CONNECT_READ = 1'b1,
    parameter M07_CONNECT_WRITE = 1'b1,
    parameter M07_SECURE = 1'b0,
    parameter M08_BASE_ADDR = 0,
    parameter M08_ADDR_WIDTH = {M_REGIONS{32'd24}},
    parameter M08_CONNECT_READ = 1'b1,
    parameter M08_CONNECT_WRITE = 1'b1,
    parameter M08_SECURE = 1'b0,
    parameter M09_BASE_ADDR = 0,
    parameter M09_ADDR_WIDTH = {M_REGIONS{32'd24}},
    parameter M09_CONNECT_READ = 1'b1,
    parameter M09_CONNECT_WRITE = 1'b1,
    parameter M09_SECURE = 1'b0,
    parameter M10_BASE_ADDR = 0,
    parameter M10_ADDR_WIDTH = {M_REGIONS{32'd24}},
    parameter M10_CONNECT_READ = 1'b1,
    parameter M10_CONNECT_WRITE = 1'b1,
    parameter M10_SECURE = 1'b0,
    parameter M11_BASE_ADDR = 0,
    parameter M11_ADDR_WIDTH = {M_REGIONS{32'd24}},
    parameter M11_CONNECT_READ = 1'b1,
    parameter M11_CONNECT_WRITE = 1'b1,
    parameter M11_SECURE = 1'b0,
    parameter M12_BASE_ADDR = 0,
    parameter M12_ADDR_WIDTH = {M_REGIONS{32'd24}},
    parameter M12_CONNECT_READ = 1'b1,
    parameter M12_CONNECT_WRITE = 1'b1,
    parameter M12_SECURE = 1'b0,
    parameter M13_BASE_ADDR = 0,
    parameter M13_ADDR_WIDTH = {M_REGIONS{32'd24}},
    parameter M13_CONNECT_READ = 1'b1,
    parameter M13_CONNECT_WRITE = 1'b1,
    parameter M13_SECURE = 1'b0,
    parameter M14_BASE_ADDR = 0,
    parameter M14_ADDR_WIDTH = {M_REGIONS{32'd24}},
    parameter M14_CONNECT_READ = 1'b1,
    parameter M14_CONNECT_WRITE = 1'b1,
    parameter M14_SECURE = 1'b0,
    parameter M15_BASE_ADDR = 0,
    parameter M15_ADDR_WIDTH = {M_REGIONS{32'd24}},
    parameter M15_CONNECT_READ = 1'b1,
    parameter M15_CONNECT_WRITE = 1'b1,
    parameter M15_SECURE = 1'b0,
    parameter M16_BASE_ADDR = 0,
    parameter M16_ADDR_WIDTH = {M_REGIONS{32'd24}},
    parameter M16_CONNECT_READ = 1'b1,
    parameter M16_CONNECT_WRITE = 1'b1,
    parameter M16_SECURE = 1'b0,
    parameter M17_BASE_ADDR = 0,
    parameter M17_ADDR_WIDTH = {M_REGIONS{32'd24}},
    parameter M17_CONNECT_READ = 1'b1,
    parameter M17_CONNECT_WRITE = 1'b1,
    parameter M17_SECURE = 1'b0,
    parameter M18_BASE_ADDR = 0,
    parameter M18_ADDR_WIDTH = {M_REGIONS{32'd24}},
    parameter M18_CONNECT_READ = 1'b1,
    parameter M18_CONNECT_WRITE = 1'b1,
    parameter M18_SECURE = 1'b0,
    parameter M19_BASE_ADDR = 0,
    parameter M19_ADDR_WIDTH = {M_REGIONS{32'd24}},
    parameter M19_CONNECT_READ = 1'b1,
    parameter M19_CONNECT_WRITE = 1'b1,
    parameter M19_SECURE = 1'b0,
    parameter M20_BASE_ADDR = 0,
    parameter M20_ADDR_WIDTH = {M_REGIONS{32'd24}},
    parameter M20_CONNECT_READ = 1'b1,
    parameter M20_CONNECT_WRITE = 1'b1,
    parameter M20_SECURE = 1'b0,
    parameter M21_BASE_ADDR = 0,
    parameter M21_ADDR_WIDTH = {M_REGIONS{32'd24}},
    parameter M21_CONNECT_READ = 1'b1,
    parameter M21_CONNECT_WRITE = 1'b1,
    parameter M21_SECURE = 1'b0,
    parameter M22_BASE_ADDR = 0,
    parameter M22_ADDR_WIDTH = {M_REGIONS{32'd24}},
    parameter M22_CONNECT_READ = 1'b1,
    parameter M22_CONNECT_WRITE = 1'b1,
    parameter M22_SECURE = 1'b0,
    parameter M23_BASE_ADDR = 0,
    parameter M23_ADDR_WIDTH = {M_REGIONS{32'd24}},
    parameter M23_CONNECT_READ = 1'b1,
    parameter M23_CONNECT_WRITE = 1'b1,
    parameter M23_SECURE = 1'b0
)
(
    input  wire                     clk,
    input  wire                     rst,

    /*
     * AXI lite slave interfaces
     */
    input  wire [ADDR_WIDTH-1:0]    s00_axil_awaddr,
    input  wire [2:0]               s00_axil_awprot,
    input  wire                     s00_axil_awvalid,
    output wire                     s00_axil_awready,
    input  wire [DATA_WIDTH-1:0]    s00_axil_wdata,
    input  wire [STRB_WIDTH-1:0]    s00_axil_wstrb,
    input  wire                     s00_axil_wvalid,
    output wire                     s00_axil_wready,
    output wire [1:0]               s00_axil_bresp,
    output wire                     s00_axil_bvalid,
    input  wire                     s00_axil_bready,
    input  wire [ADDR_WIDTH-1:0]    s00_axil_araddr,
    input  wire [2:0]               s00_axil_arprot,
    input  wire                     s00_axil_arvalid,
    output wire                     s00_axil_arready,
    output wire [DATA_WIDTH-1:0]    s00_axil_rdata,
    output wire [1:0]               s00_axil_rresp,
    output wire                     s00_axil_rvalid,
    input  wire                     s00_axil_rready,

    /*
     * AXI lite master interfaces
     */
    output wire [ADDR_WIDTH-1:0]    m00_axil_awaddr,
    output wire [2:0]               m00_axil_awprot,
    output wire                     m00_axil_awvalid,
    input  wire                     m00_axil_awready,
    output wire [DATA_WIDTH-1:0]    m00_axil_wdata,
    output wire [STRB_WIDTH-1:0]    m00_axil_wstrb,
    output wire                     m00_axil_wvalid,
    input  wire                     m00_axil_wready,
    input  wire [1:0]               m00_axil_bresp,
    input  wire                     m00_axil_bvalid,
    output wire                     m00_axil_bready,
    output wire [ADDR_WIDTH-1:0]    m00_axil_araddr,
    output wire [2:0]               m00_axil_arprot,
    output wire                     m00_axil_arvalid,
    input  wire                     m00_axil_arready,
    input  wire [DATA_WIDTH-1:0]    m00_axil_rdata,
    input  wire [1:0]               m00_axil_rresp,
    input  wire                     m00_axil_rvalid,
    output wire                     m00_axil_rready,

    output wire [ADDR_WIDTH-1:0]    m01_axil_awaddr,
    output wire [2:0]               m01_axil_awprot,
    output wire                     m01_axil_awvalid,
    input  wire                     m01_axil_awready,
    output wire [DATA_WIDTH-1:0]    m01_axil_wdata,
    output wire [STRB_WIDTH-1:0]    m01_axil_wstrb,
    output wire                     m01_axil_wvalid,
    input  wire                     m01_axil_wready,
    input  wire [1:0]               m01_axil_bresp,
    input  wire                     m01_axil_bvalid,
    output wire                     m01_axil_bready,
    output wire [ADDR_WIDTH-1:0]    m01_axil_araddr,
    output wire [2:0]               m01_axil_arprot,
    output wire                     m01_axil_arvalid,
    input  wire                     m01_axil_arready,
    input  wire [DATA_WIDTH-1:0]    m01_axil_rdata,
    input  wire [1:0]               m01_axil_rresp,
    input  wire                     m01_axil_rvalid,
    output wire                     m01_axil_rready,

    output wire [ADDR_WIDTH-1:0]    m02_axil_awaddr,
    output wire [2:0]               m02_axil_awprot,
    output wire                     m02_axil_awvalid,
    input  wire                     m02_axil_awready,
    output wire [DATA_WIDTH-1:0]    m02_axil_wdata,
    output wire [STRB_WIDTH-1:0]    m02_axil_wstrb,
    output wire                     m02_axil_wvalid,
    input  wire                     m02_axil_wready,
    input  wire [1:0]               m02_axil_bresp,
    input  wire                     m02_axil_bvalid,
    output wire                     m02_axil_bready,
    output wire [ADDR_WIDTH-1:0]    m02_axil_araddr,
    output wire [2:0]               m02_axil_arprot,
    output wire                     m02_axil_arvalid,
    input  wire                     m02_axil_arready,
    input  wire [DATA_WIDTH-1:0]    m02_axil_rdata,
    input  wire [1:0]               m02_axil_rresp,
    input  wire                     m02_axil_rvalid,
    output wire                     m02_axil_rready,

    output wire [ADDR_WIDTH-1:0]    m03_axil_awaddr,
    output wire [2:0]               m03_axil_awprot,
    output wire                     m03_axil_awvalid,
    input  wire                     m03_axil_awready,
    output wire [DATA_WIDTH-1:0]    m03_axil_wdata,
    output wire [STRB_WIDTH-1:0]    m03_axil_wstrb,
    output wire                     m03_axil_wvalid,
    input  wire                     m03_axil_wready,
    input  wire [1:0]               m03_axil_bresp,
    input  wire                     m03_axil_bvalid,
    output wire                     m03_axil_bready,
    output wire [ADDR_WIDTH-1:0]    m03_axil_araddr,
    output wire [2:0]               m03_axil_arprot,
    output wire                     m03_axil_arvalid,
    input  wire                     m03_axil_arready,
    input  wire [DATA_WIDTH-1:0]    m03_axil_rdata,
    input  wire [1:0]               m03_axil_rresp,
    input  wire                     m03_axil_rvalid,
    output wire                     m03_axil_rready,

    output wire [ADDR_WIDTH-1:0]    m04_axil_awaddr,
    output wire [2:0]               m04_axil_awprot,
    output wire                     m04_axil_awvalid,
    input  wire                     m04_axil_awready,
    output wire [DATA_WIDTH-1:0]    m04_axil_wdata,
    output wire [STRB_WIDTH-1:0]    m04_axil_wstrb,
    output wire                     m04_axil_wvalid,
    input  wire                     m04_axil_wready,
    input  wire [1:0]               m04_axil_bresp,
    input  wire                     m04_axil_bvalid,
    output wire                     m04_axil_bready,
    output wire [ADDR_WIDTH-1:0]    m04_axil_araddr,
    output wire [2:0]               m04_axil_arprot,
    output wire                     m04_axil_arvalid,
    input  wire                     m04_axil_arready,
    input  wire [DATA_WIDTH-1:0]    m04_axil_rdata,
    input  wire [1:0]               m04_axil_rresp,
    input  wire                     m04_axil_rvalid,
    output wire                     m04_axil_rready,

    output wire [ADDR_WIDTH-1:0]    m05_axil_awaddr,
    output wire [2:0]               m05_axil_awprot,
    output wire                     m05_axil_awvalid,
    input  wire                     m05_axil_awready,
    output wire [DATA_WIDTH-1:0]    m05_axil_wdata,
    output wire [STRB_WIDTH-1:0]    m05_axil_wstrb,
    output wire                     m05_axil_wvalid,
    input  wire                     m05_axil_wready,
    input  wire [1:0]               m05_axil_bresp,
    input  wire                     m05_axil_bvalid,
    output wire                     m05_axil_bready,
    output wire [ADDR_WIDTH-1:0]    m05_axil_araddr,
    output wire [2:0]               m05_axil_arprot,
    output wire                     m05_axil_arvalid,
    input  wire                     m05_axil_arready,
    input  wire [DATA_WIDTH-1:0]    m05_axil_rdata,
    input  wire [1:0]               m05_axil_rresp,
    input  wire                     m05_axil_rvalid,
    output wire                     m05_axil_rready,

    output wire [ADDR_WIDTH-1:0]    m06_axil_awaddr,
    output wire [2:0]               m06_axil_awprot,
    output wire                     m06_axil_awvalid,
    input  wire                     m06_axil_awready,
    output wire [DATA_WIDTH-1:0]    m06_axil_wdata,
    output wire [STRB_WIDTH-1:0]    m06_axil_wstrb,
    output wire                     m06_axil_wvalid,
    input  wire                     m06_axil_wready,
    input  wire [1:0]               m06_axil_bresp,
    input  wire                     m06_axil_bvalid,
    output wire                     m06_axil_bready,
    output wire [ADDR_WIDTH-1:0]    m06_axil_araddr,
    output wire [2:0]               m06_axil_arprot,
    output wire                     m06_axil_arvalid,
    input  wire                     m06_axil_arready,
    input  wire [DATA_WIDTH-1:0]    m06_axil_rdata,
    input  wire [1:0]               m06_axil_rresp,
    input  wire                     m06_axil_rvalid,
    output wire                     m06_axil_rready,

    output wire [ADDR_WIDTH-1:0]    m07_axil_awaddr,
    output wire [2:0]               m07_axil_awprot,
    output wire                     m07_axil_awvalid,
    input  wire                     m07_axil_awready,
    output wire [DATA_WIDTH-1:0]    m07_axil_wdata,
    output wire [STRB_WIDTH-1:0]    m07_axil_wstrb,
    output wire                     m07_axil_wvalid,
    input  wire                     m07_axil_wready,
    input  wire [1:0]               m07_axil_bresp,
    input  wire                     m07_axil_bvalid,
    output wire                     m07_axil_bready,
    output wire [ADDR_WIDTH-1:0]    m07_axil_araddr,
    output wire [2:0]               m07_axil_arprot,
    output wire                     m07_axil_arvalid,
    input  wire                     m07_axil_arready,
    input  wire [DATA_WIDTH-1:0]    m07_axil_rdata,
    input  wire [1:0]               m07_axil_rresp,
    input  wire                     m07_axil_rvalid,
    output wire                     m07_axil_rready,

    output wire [ADDR_WIDTH-1:0]    m08_axil_awaddr,
    output wire [2:0]               m08_axil_awprot,
    output wire                     m08_axil_awvalid,
    input  wire                     m08_axil_awready,
    output wire [DATA_WIDTH-1:0]    m08_axil_wdata,
    output wire [STRB_WIDTH-1:0]    m08_axil_wstrb,
    output wire                     m08_axil_wvalid,
    input  wire                     m08_axil_wready,
    input  wire [1:0]               m08_axil_bresp,
    input  wire                     m08_axil_bvalid,
    output wire                     m08_axil_bready,
    output wire [ADDR_WIDTH-1:0]    m08_axil_araddr,
    output wire [2:0]               m08_axil_arprot,
    output wire                     m08_axil_arvalid,
    input  wire                     m08_axil_arready,
    input  wire [DATA_WIDTH-1:0]    m08_axil_rdata,
    input  wire [1:0]               m08_axil_rresp,
    input  wire                     m08_axil_rvalid,
    output wire                     m08_axil_rready,

    output wire [ADDR_WIDTH-1:0]    m09_axil_awaddr,
    output wire [2:0]               m09_axil_awprot,
    output wire                     m09_axil_awvalid,
    input  wire                     m09_axil_awready,
    output wire [DATA_WIDTH-1:0]    m09_axil_wdata,
    output wire [STRB_WIDTH-1:0]    m09_axil_wstrb,
    output wire                     m09_axil_wvalid,
    input  wire                     m09_axil_wready,
    input  wire [1:0]               m09_axil_bresp,
    input  wire                     m09_axil_bvalid,
    output wire                     m09_axil_bready,
    output wire [ADDR_WIDTH-1:0]    m09_axil_araddr,
    output wire [2:0]               m09_axil_arprot,
    output wire                     m09_axil_arvalid,
    input  wire                     m09_axil_arready,
    input  wire [DATA_WIDTH-1:0]    m09_axil_rdata,
    input  wire [1:0]               m09_axil_rresp,
    input  wire                     m09_axil_rvalid,
    output wire                     m09_axil_rready,

    output wire [ADDR_WIDTH-1:0]    m10_axil_awaddr,
    output wire [2:0]               m10_axil_awprot,
    output wire                     m10_axil_awvalid,
    input  wire                     m10_axil_awready,
    output wire [DATA_WIDTH-1:0]    m10_axil_wdata,
    output wire [STRB_WIDTH-1:0]    m10_axil_wstrb,
    output wire                     m10_axil_wvalid,
    input  wire                     m10_axil_wready,
    input  wire [1:0]               m10_axil_bresp,
    input  wire                     m10_axil_bvalid,
    output wire                     m10_axil_bready,
    output wire [ADDR_WIDTH-1:0]    m10_axil_araddr,
    output wire [2:0]               m10_axil_arprot,
    output wire                     m10_axil_arvalid,
    input  wire                     m10_axil_arready,
    input  wire [DATA_WIDTH-1:0]    m10_axil_rdata,
    input  wire [1:0]               m10_axil_rresp,
    input  wire                     m10_axil_rvalid,
    output wire                     m10_axil_rready,

    output wire [ADDR_WIDTH-1:0]    m11_axil_awaddr,
    output wire [2:0]               m11_axil_awprot,
    output wire                     m11_axil_awvalid,
    input  wire                     m11_axil_awready,
    output wire [DATA_WIDTH-1:0]    m11_axil_wdata,
    output wire [STRB_WIDTH-1:0]    m11_axil_wstrb,
    output wire                     m11_axil_wvalid,
    input  wire                     m11_axil_wready,
    input  wire [1:0]               m11_axil_bresp,
    input  wire                     m11_axil_bvalid,
    output wire                     m11_axil_bready,
    output wire [ADDR_WIDTH-1:0]    m11_axil_araddr,
    output wire [2:0]               m11_axil_arprot,
    output wire                     m11_axil_arvalid,
    input  wire                     m11_axil_arready,
    input  wire [DATA_WIDTH-1:0]    m11_axil_rdata,
    input  wire [1:0]               m11_axil_rresp,
    input  wire                     m11_axil_rvalid,
    output wire                     m11_axil_rready,

    output wire [ADDR_WIDTH-1:0]    m12_axil_awaddr,
    output wire [2:0]               m12_axil_awprot,
    output wire                     m12_axil_awvalid,
    input  wire                     m12_axil_awready,
    output wire [DATA_WIDTH-1:0]    m12_axil_wdata,
    output wire [STRB_WIDTH-1:0]    m12_axil_wstrb,
    output wire                     m12_axil_wvalid,
    input  wire                     m12_axil_wready,
    input  wire [1:0]               m12_axil_bresp,
    input  wire                     m12_axil_bvalid,
    output wire                     m12_axil_bready,
    output wire [ADDR_WIDTH-1:0]    m12_axil_araddr,
    output wire [2:0]               m12_axil_arprot,
    output wire                     m12_axil_arvalid,
    input  wire                     m12_axil_arready,
    input  wire [DATA_WIDTH-1:0]    m12_axil_rdata,
    input  wire [1:0]               m12_axil_rresp,
    input  wire                     m12_axil_rvalid,
    output wire                     m12_axil_rready,

    output wire [ADDR_WIDTH-1:0]    m13_axil_awaddr,
    output wire [2:0]               m13_axil_awprot,
    output wire                     m13_axil_awvalid,
    input  wire                     m13_axil_awready,
    output wire [DATA_WIDTH-1:0]    m13_axil_wdata,
    output wire [STRB_WIDTH-1:0]    m13_axil_wstrb,
    output wire                     m13_axil_wvalid,
    input  wire                     m13_axil_wready,
    input  wire [1:0]               m13_axil_bresp,
    input  wire                     m13_axil_bvalid,
    output wire                     m13_axil_bready,
    output wire [ADDR_WIDTH-1:0]    m13_axil_araddr,
    output wire [2:0]               m13_axil_arprot,
    output wire                     m13_axil_arvalid,
    input  wire                     m13_axil_arready,
    input  wire [DATA_WIDTH-1:0]    m13_axil_rdata,
    input  wire [1:0]               m13_axil_rresp,
    input  wire                     m13_axil_rvalid,
    output wire                     m13_axil_rready,

    output wire [ADDR_WIDTH-1:0]    m14_axil_awaddr,
    output wire [2:0]               m14_axil_awprot,
    output wire                     m14_axil_awvalid,
    input  wire                     m14_axil_awready,
    output wire [DATA_WIDTH-1:0]    m14_axil_wdata,
    output wire [STRB_WIDTH-1:0]    m14_axil_wstrb,
    output wire                     m14_axil_wvalid,
    input  wire                     m14_axil_wready,
    input  wire [1:0]               m14_axil_bresp,
    input  wire                     m14_axil_bvalid,
    output wire                     m14_axil_bready,
    output wire [ADDR_WIDTH-1:0]    m14_axil_araddr,
    output wire [2:0]               m14_axil_arprot,
    output wire                     m14_axil_arvalid,
    input  wire                     m14_axil_arready,
    input  wire [DATA_WIDTH-1:0]    m14_axil_rdata,
    input  wire [1:0]               m14_axil_rresp,
    input  wire                     m14_axil_rvalid,
    output wire                     m14_axil_rready,

    output wire [ADDR_WIDTH-1:0]    m15_axil_awaddr,
    output wire [2:0]               m15_axil_awprot,
    output wire                     m15_axil_awvalid,
    input  wire                     m15_axil_awready,
    output wire [DATA_WIDTH-1:0]    m15_axil_wdata,
    output wire [STRB_WIDTH-1:0]    m15_axil_wstrb,
    output wire                     m15_axil_wvalid,
    input  wire                     m15_axil_wready,
    input  wire [1:0]               m15_axil_bresp,
    input  wire                     m15_axil_bvalid,
    output wire                     m15_axil_bready,
    output wire [ADDR_WIDTH-1:0]    m15_axil_araddr,
    output wire [2:0]               m15_axil_arprot,
    output wire                     m15_axil_arvalid,
    input  wire                     m15_axil_arready,
    input  wire [DATA_WIDTH-1:0]    m15_axil_rdata,
    input  wire [1:0]               m15_axil_rresp,
    input  wire                     m15_axil_rvalid,
    output wire                     m15_axil_rready,

    output wire [ADDR_WIDTH-1:0]    m16_axil_awaddr,
    output wire [2:0]               m16_axil_awprot,
    output wire                     m16_axil_awvalid,
    input  wire                     m16_axil_awready,
    output wire [DATA_WIDTH-1:0]    m16_axil_wdata,
    output wire [STRB_WIDTH-1:0]    m16_axil_wstrb,
    output wire                     m16_axil_wvalid,
    input  wire                     m16_axil_wready,
    input  wire [1:0]               m16_axil_bresp,
    input  wire                     m16_axil_bvalid,
    output wire                     m16_axil_bready,
    output wire [ADDR_WIDTH-1:0]    m16_axil_araddr,
    output wire [2:0]               m16_axil_arprot,
    output wire                     m16_axil_arvalid,
    input  wire                     m16_axil_arready,
    input  wire [DATA_WIDTH-1:0]    m16_axil_rdata,
    input  wire [1:0]               m16_axil_rresp,
    input  wire                     m16_axil_rvalid,
    output wire                     m16_axil_rready,

    output wire [ADDR_WIDTH-1:0]    m17_axil_awaddr,
    output wire [2:0]               m17_axil_awprot,
    output wire                     m17_axil_awvalid,
    input  wire                     m17_axil_awready,
    output wire [DATA_WIDTH-1:0]    m17_axil_wdata,
    output wire [STRB_WIDTH-1:0]    m17_axil_wstrb,
    output wire                     m17_axil_wvalid,
    input  wire                     m17_axil_wready,
    input  wire [1:0]               m17_axil_bresp,
    input  wire                     m17_axil_bvalid,
    output wire                     m17_axil_bready,
    output wire [ADDR_WIDTH-1:0]    m17_axil_araddr,
    output wire [2:0]               m17_axil_arprot,
    output wire                     m17_axil_arvalid,
    input  wire                     m17_axil_arready,
    input  wire [DATA_WIDTH-1:0]    m17_axil_rdata,
    input  wire [1:0]               m17_axil_rresp,
    input  wire                     m17_axil_rvalid,
    output wire                     m17_axil_rready,

    output wire [ADDR_WIDTH-1:0]    m18_axil_awaddr,
    output wire [2:0]               m18_axil_awprot,
    output wire                     m18_axil_awvalid,
    input  wire                     m18_axil_awready,
    output wire [DATA_WIDTH-1:0]    m18_axil_wdata,
    output wire [STRB_WIDTH-1:0]    m18_axil_wstrb,
    output wire                     m18_axil_wvalid,
    input  wire                     m18_axil_wready,
    input  wire [1:0]               m18_axil_bresp,
    input  wire                     m18_axil_bvalid,
    output wire                     m18_axil_bready,
    output wire [ADDR_WIDTH-1:0]    m18_axil_araddr,
    output wire [2:0]               m18_axil_arprot,
    output wire                     m18_axil_arvalid,
    input  wire                     m18_axil_arready,
    input  wire [DATA_WIDTH-1:0]    m18_axil_rdata,
    input  wire [1:0]               m18_axil_rresp,
    input  wire                     m18_axil_rvalid,
    output wire                     m18_axil_rready,

    output wire [ADDR_WIDTH-1:0]    m19_axil_awaddr,
    output wire [2:0]               m19_axil_awprot,
    output wire                     m19_axil_awvalid,
    input  wire                     m19_axil_awready,
    output wire [DATA_WIDTH-1:0]    m19_axil_wdata,
    output wire [STRB_WIDTH-1:0]    m19_axil_wstrb,
    output wire                     m19_axil_wvalid,
    input  wire                     m19_axil_wready,
    input  wire [1:0]               m19_axil_bresp,
    input  wire                     m19_axil_bvalid,
    output wire                     m19_axil_bready,
    output wire [ADDR_WIDTH-1:0]    m19_axil_araddr,
    output wire [2:0]               m19_axil_arprot,
    output wire                     m19_axil_arvalid,
    input  wire                     m19_axil_arready,
    input  wire [DATA_WIDTH-1:0]    m19_axil_rdata,
    input  wire [1:0]               m19_axil_rresp,
    input  wire                     m19_axil_rvalid,
    output wire                     m19_axil_rready,

    output wire [ADDR_WIDTH-1:0]    m20_axil_awaddr,
    output wire [2:0]               m20_axil_awprot,
    output wire                     m20_axil_awvalid,
    input  wire                     m20_axil_awready,
    output wire [DATA_WIDTH-1:0]    m20_axil_wdata,
    output wire [STRB_WIDTH-1:0]    m20_axil_wstrb,
    output wire                     m20_axil_wvalid,
    input  wire                     m20_axil_wready,
    input  wire [1:0]               m20_axil_bresp,
    input  wire                     m20_axil_bvalid,
    output wire                     m20_axil_bready,
    output wire [ADDR_WIDTH-1:0]    m20_axil_araddr,
    output wire [2:0]               m20_axil_arprot,
    output wire                     m20_axil_arvalid,
    input  wire                     m20_axil_arready,
    input  wire [DATA_WIDTH-1:0]    m20_axil_rdata,
    input  wire [1:0]               m20_axil_rresp,
    input  wire                     m20_axil_rvalid,
    output wire                     m20_axil_rready,

    output wire [ADDR_WIDTH-1:0]    m21_axil_awaddr,
    output wire [2:0]               m21_axil_awprot,
    output wire                     m21_axil_awvalid,
    input  wire                     m21_axil_awready,
    output wire [DATA_WIDTH-1:0]    m21_axil_wdata,
    output wire [STRB_WIDTH-1:0]    m21_axil_wstrb,
    output wire                     m21_axil_wvalid,
    input  wire                     m21_axil_wready,
    input  wire [1:0]               m21_axil_bresp,
    input  wire                     m21_axil_bvalid,
    output wire                     m21_axil_bready,
    output wire [ADDR_WIDTH-1:0]    m21_axil_araddr,
    output wire [2:0]               m21_axil_arprot,
    output wire                     m21_axil_arvalid,
    input  wire                     m21_axil_arready,
    input  wire [DATA_WIDTH-1:0]    m21_axil_rdata,
    input  wire [1:0]               m21_axil_rresp,
    input  wire                     m21_axil_rvalid,
    output wire                     m21_axil_rready,

    output wire [ADDR_WIDTH-1:0]    m22_axil_awaddr,
    output wire [2:0]               m22_axil_awprot,
    output wire                     m22_axil_awvalid,
    input  wire                     m22_axil_awready,
    output wire [DATA_WIDTH-1:0]    m22_axil_wdata,
    output wire [STRB_WIDTH-1:0]    m22_axil_wstrb,
    output wire                     m22_axil_wvalid,
    input  wire                     m22_axil_wready,
    input  wire [1:0]               m22_axil_bresp,
    input  wire                     m22_axil_bvalid,
    output wire                     m22_axil_bready,
    output wire [ADDR_WIDTH-1:0]    m22_axil_araddr,
    output wire [2:0]               m22_axil_arprot,
    output wire                     m22_axil_arvalid,
    input  wire                     m22_axil_arready,
    input  wire [DATA_WIDTH-1:0]    m22_axil_rdata,
    input  wire [1:0]               m22_axil_rresp,
    input  wire                     m22_axil_rvalid,
    output wire                     m22_axil_rready,

    output wire [ADDR_WIDTH-1:0]    m23_axil_awaddr,
    output wire [2:0]               m23_axil_awprot,
    output wire                     m23_axil_awvalid,
    input  wire                     m23_axil_awready,
    output wire [DATA_WIDTH-1:0]    m23_axil_wdata,
    output wire [STRB_WIDTH-1:0]    m23_axil_wstrb,
    output wire                     m23_axil_wvalid,
    input  wire                     m23_axil_wready,
    input  wire [1:0]               m23_axil_bresp,
    input  wire                     m23_axil_bvalid,
    output wire                     m23_axil_bready,
    output wire [ADDR_WIDTH-1:0]    m23_axil_araddr,
    output wire [2:0]               m23_axil_arprot,
    output wire                     m23_axil_arvalid,
    input  wire                     m23_axil_arready,
    input  wire [DATA_WIDTH-1:0]    m23_axil_rdata,
    input  wire [1:0]               m23_axil_rresp,
    input  wire                     m23_axil_rvalid,
    output wire                     m23_axil_rready
);

localparam S_COUNT = 1;
localparam M_COUNT = 24;

// parameter sizing helpers
function [ADDR_WIDTH*M_REGIONS-1:0] w_a_r(input [ADDR_WIDTH*M_REGIONS-1:0] val);
    w_a_r = val;
endfunction

function [32*M_REGIONS-1:0] w_32_r(input [32*M_REGIONS-1:0] val);
    w_32_r = val;
endfunction

function [S_COUNT-1:0] w_s(input [S_COUNT-1:0] val);
    w_s = val;
endfunction

function w_1(input val);
    w_1 = val;
endfunction

axil_interconnect #(
    .S_COUNT(S_COUNT),
    .M_COUNT(M_COUNT),
    .DATA_WIDTH(DATA_WIDTH),
    .ADDR_WIDTH(ADDR_WIDTH),
    .STRB_WIDTH(STRB_WIDTH),
    .M_REGIONS(M_REGIONS),
    .M_BASE_ADDR({ w_a_r(M23_BASE_ADDR), w_a_r(M22_BASE_ADDR), w_a_r(M21_BASE_ADDR), w_a_r(M20_BASE_ADDR), w_a_r(M19_BASE_ADDR), w_a_r(M18_BASE_ADDR), w_a_r(M17_BASE_ADDR), w_a_r(M16_BASE_ADDR), w_a_r(M15_BASE_ADDR), w_a_r(M14_BASE_ADDR), w_a_r(M13_BASE_ADDR), w_a_r(M12_BASE_ADDR), w_a_r(M11_BASE_ADDR), w_a_r(M10_BASE_ADDR), w_a_r(M09_BASE_ADDR), w_a_r(M08_BASE_ADDR), w_a_r(M07_BASE_ADDR), w_a_r(M06_BASE_ADDR), w_a_r(M05_BASE_ADDR), w_a_r(M04_BASE_ADDR), w_a_r(M03_BASE_ADDR), w_a_r(M02_BASE_ADDR), w_a_r(M01_BASE_ADDR), w_a_r(M00_BASE_ADDR) }),
    .M_ADDR_WIDTH({ w_32_r(M23_ADDR_WIDTH), w_32_r(M22_ADDR_WIDTH), w_32_r(M21_ADDR_WIDTH), w_32_r(M20_ADDR_WIDTH), w_32_r(M19_ADDR_WIDTH), w_32_r(M18_ADDR_WIDTH), w_32_r(M17_ADDR_WIDTH), w_32_r(M16_ADDR_WIDTH), w_32_r(M15_ADDR_WIDTH), w_32_r(M14_ADDR_WIDTH), w_32_r(M13_ADDR_WIDTH), w_32_r(M12_ADDR_WIDTH), w_32_r(M11_ADDR_WIDTH), w_32_r(M10_ADDR_WIDTH), w_32_r(M09_ADDR_WIDTH), w_32_r(M08_ADDR_WIDTH), w_32_r(M07_ADDR_WIDTH), w_32_r(M06_ADDR_WIDTH), w_32_r(M05_ADDR_WIDTH), w_32_r(M04_ADDR_WIDTH), w_32_r(M03_ADDR_WIDTH), w_32_r(M02_ADDR_WIDTH), w_32_r(M01_ADDR_WIDTH), w_32_r(M00_ADDR_WIDTH) }),
    .M_CONNECT_READ({ w_s(M23_CONNECT_READ), w_s(M22_CONNECT_READ), w_s(M21_CONNECT_READ), w_s(M20_CONNECT_READ), w_s(M19_CONNECT_READ), w_s(M18_CONNECT_READ), w_s(M17_CONNECT_READ), w_s(M16_CONNECT_READ), w_s(M15_CONNECT_READ), w_s(M14_CONNECT_READ), w_s(M13_CONNECT_READ), w_s(M12_CONNECT_READ), w_s(M11_CONNECT_READ), w_s(M10_CONNECT_READ), w_s(M09_CONNECT_READ), w_s(M08_CONNECT_READ), w_s(M07_CONNECT_READ), w_s(M06_CONNECT_READ), w_s(M05_CONNECT_READ), w_s(M04_CONNECT_READ), w_s(M03_CONNECT_READ), w_s(M02_CONNECT_READ), w_s(M01_CONNECT_READ), w_s(M00_CONNECT_READ) }),
    .M_CONNECT_WRITE({ w_s(M23_CONNECT_WRITE), w_s(M22_CONNECT_WRITE), w_s(M21_CONNECT_WRITE), w_s(M20_CONNECT_WRITE), w_s(M19_CONNECT_WRITE), w_s(M18_CONNECT_WRITE), w_s(M17_CONNECT_WRITE), w_s(M16_CONNECT_WRITE), w_s(M15_CONNECT_WRITE), w_s(M14_CONNECT_WRITE), w_s(M13_CONNECT_WRITE), w_s(M12_CONNECT_WRITE), w_s(M11_CONNECT_WRITE), w_s(M10_CONNECT_WRITE), w_s(M09_CONNECT_WRITE), w_s(M08_CONNECT_WRITE), w_s(M07_CONNECT_WRITE), w_s(M06_CONNECT_WRITE), w_s(M05_CONNECT_WRITE), w_s(M04_CONNECT_WRITE), w_s(M03_CONNECT_WRITE), w_s(M02_CONNECT_WRITE), w_s(M01_CONNECT_WRITE), w_s(M00_CONNECT_WRITE) }),
    .M_SECURE({ w_1(M23_SECURE), w_1(M22_SECURE), w_1(M21_SECURE), w_1(M20_SECURE), w_1(M19_SECURE), w_1(M18_SECURE), w_1(M17_SECURE), w_1(M16_SECURE), w_1(M15_SECURE), w_1(M14_SECURE), w_1(M13_SECURE), w_1(M12_SECURE), w_1(M11_SECURE), w_1(M10_SECURE), w_1(M09_SECURE), w_1(M08_SECURE), w_1(M07_SECURE), w_1(M06_SECURE), w_1(M05_SECURE), w_1(M04_SECURE), w_1(M03_SECURE), w_1(M02_SECURE), w_1(M01_SECURE), w_1(M00_SECURE) })
)
axil_interconnect_inst (
    .clk(clk),
    .rst(rst),
    .s_axil_awaddr({ s00_axil_awaddr }),
    .s_axil_awprot({ s00_axil_awprot }),
    .s_axil_awvalid({ s00_axil_awvalid }),
    .s_axil_awready({ s00_axil_awready }),
    .s_axil_wdata({ s00_axil_wdata }),
    .s_axil_wstrb({ s00_axil_wstrb }),
    .s_axil_wvalid({ s00_axil_wvalid }),
    .s_axil_wready({ s00_axil_wready }),
    .s_axil_bresp({ s00_axil_bresp }),
    .s_axil_bvalid({ s00_axil_bvalid }),
    .s_axil_bready({ s00_axil_bready }),
    .s_axil_araddr({ s00_axil_araddr }),
    .s_axil_arprot({ s00_axil_arprot }),
    .s_axil_arvalid({ s00_axil_arvalid }),
    .s_axil_arready({ s00_axil_arready }),
    .s_axil_rdata({ s00_axil_rdata }),
    .s_axil_rresp({ s00_axil_rresp }),
    .s_axil_rvalid({ s00_axil_rvalid }),
    .s_axil_rready({ s00_axil_rready }),
    .m_axil_awaddr({ m23_axil_awaddr, m22_axil_awaddr, m21_axil_awaddr, m20_axil_awaddr, m19_axil_awaddr, m18_axil_awaddr, m17_axil_awaddr, m16_axil_awaddr, m15_axil_awaddr, m14_axil_awaddr, m13_axil_awaddr, m12_axil_awaddr, m11_axil_awaddr, m10_axil_awaddr, m09_axil_awaddr, m08_axil_awaddr, m07_axil_awaddr, m06_axil_awaddr, m05_axil_awaddr, m04_axil_awaddr, m03_axil_awaddr, m02_axil_awaddr, m01_axil_awaddr, m00_axil_awaddr }),
    .m_axil_awprot({ m23_axil_awprot, m22_axil_awprot, m21_axil_awprot, m20_axil_awprot, m19_axil_awprot, m18_axil_awprot, m17_axil_awprot, m16_axil_awprot, m15_axil_awprot, m14_axil_awprot, m13_axil_awprot, m12_axil_awprot, m11_axil_awprot, m10_axil_awprot, m09_axil_awprot, m08_axil_awprot, m07_axil_awprot, m06_axil_awprot, m05_axil_awprot, m04_axil_awprot, m03_axil_awprot, m02_axil_awprot, m01_axil_awprot, m00_axil_awprot }),
    .m_axil_awvalid({ m23_axil_awvalid, m22_axil_awvalid, m21_axil_awvalid, m20_axil_awvalid, m19_axil_awvalid, m18_axil_awvalid, m17_axil_awvalid, m16_axil_awvalid, m15_axil_awvalid, m14_axil_awvalid, m13_axil_awvalid, m12_axil_awvalid, m11_axil_awvalid, m10_axil_awvalid, m09_axil_awvalid, m08_axil_awvalid, m07_axil_awvalid, m06_axil_awvalid, m05_axil_awvalid, m04_axil_awvalid, m03_axil_awvalid, m02_axil_awvalid, m01_axil_awvalid, m00_axil_awvalid }),
    .m_axil_awready({ m23_axil_awready, m22_axil_awready, m21_axil_awready, m20_axil_awready, m19_axil_awready, m18_axil_awready, m17_axil_awready, m16_axil_awready, m15_axil_awready, m14_axil_awready, m13_axil_awready, m12_axil_awready, m11_axil_awready, m10_axil_awready, m09_axil_awready, m08_axil_awready, m07_axil_awready, m06_axil_awready, m05_axil_awready, m04_axil_awready, m03_axil_awready, m02_axil_awready, m01_axil_awready, m00_axil_awready }),
    .m_axil_wdata({ m23_axil_wdata, m22_axil_wdata, m21_axil_wdata, m20_axil_wdata, m19_axil_wdata, m18_axil_wdata, m17_axil_wdata, m16_axil_wdata, m15_axil_wdata, m14_axil_wdata, m13_axil_wdata, m12_axil_wdata, m11_axil_wdata, m10_axil_wdata, m09_axil_wdata, m08_axil_wdata, m07_axil_wdata, m06_axil_wdata, m05_axil_wdata, m04_axil_wdata, m03_axil_wdata, m02_axil_wdata, m01_axil_wdata, m00_axil_wdata }),
    .m_axil_wstrb({ m23_axil_wstrb, m22_axil_wstrb, m21_axil_wstrb, m20_axil_wstrb, m19_axil_wstrb, m18_axil_wstrb, m17_axil_wstrb, m16_axil_wstrb, m15_axil_wstrb, m14_axil_wstrb, m13_axil_wstrb, m12_axil_wstrb, m11_axil_wstrb, m10_axil_wstrb, m09_axil_wstrb, m08_axil_wstrb, m07_axil_wstrb, m06_axil_wstrb, m05_axil_wstrb, m04_axil_wstrb, m03_axil_wstrb, m02_axil_wstrb, m01_axil_wstrb, m00_axil_wstrb }),
    .m_axil_wvalid({ m23_axil_wvalid, m22_axil_wvalid, m21_axil_wvalid, m20_axil_wvalid, m19_axil_wvalid, m18_axil_wvalid, m17_axil_wvalid, m16_axil_wvalid, m15_axil_wvalid, m14_axil_wvalid, m13_axil_wvalid, m12_axil_wvalid, m11_axil_wvalid, m10_axil_wvalid, m09_axil_wvalid, m08_axil_wvalid, m07_axil_wvalid, m06_axil_wvalid, m05_axil_wvalid, m04_axil_wvalid, m03_axil_wvalid, m02_axil_wvalid, m01_axil_wvalid, m00_axil_wvalid }),
    .m_axil_wready({ m23_axil_wready, m22_axil_wready, m21_axil_wready, m20_axil_wready, m19_axil_wready, m18_axil_wready, m17_axil_wready, m16_axil_wready, m15_axil_wready, m14_axil_wready, m13_axil_wready, m12_axil_wready, m11_axil_wready, m10_axil_wready, m09_axil_wready, m08_axil_wready, m07_axil_wready, m06_axil_wready, m05_axil_wready, m04_axil_wready, m03_axil_wready, m02_axil_wready, m01_axil_wready, m00_axil_wready }),
    .m_axil_bresp({ m23_axil_bresp, m22_axil_bresp, m21_axil_bresp, m20_axil_bresp, m19_axil_bresp, m18_axil_bresp, m17_axil_bresp, m16_axil_bresp, m15_axil_bresp, m14_axil_bresp, m13_axil_bresp, m12_axil_bresp, m11_axil_bresp, m10_axil_bresp, m09_axil_bresp, m08_axil_bresp, m07_axil_bresp, m06_axil_bresp, m05_axil_bresp, m04_axil_bresp, m03_axil_bresp, m02_axil_bresp, m01_axil_bresp, m00_axil_bresp }),
    .m_axil_bvalid({ m23_axil_bvalid, m22_axil_bvalid, m21_axil_bvalid, m20_axil_bvalid, m19_axil_bvalid, m18_axil_bvalid, m17_axil_bvalid, m16_axil_bvalid, m15_axil_bvalid, m14_axil_bvalid, m13_axil_bvalid, m12_axil_bvalid, m11_axil_bvalid, m10_axil_bvalid, m09_axil_bvalid, m08_axil_bvalid, m07_axil_bvalid, m06_axil_bvalid, m05_axil_bvalid, m04_axil_bvalid, m03_axil_bvalid, m02_axil_bvalid, m01_axil_bvalid, m00_axil_bvalid }),
    .m_axil_bready({ m23_axil_bready, m22_axil_bready, m21_axil_bready, m20_axil_bready, m19_axil_bready, m18_axil_bready, m17_axil_bready, m16_axil_bready, m15_axil_bready, m14_axil_bready, m13_axil_bready, m12_axil_bready, m11_axil_bready, m10_axil_bready, m09_axil_bready, m08_axil_bready, m07_axil_bready, m06_axil_bready, m05_axil_bready, m04_axil_bready, m03_axil_bready, m02_axil_bready, m01_axil_bready, m00_axil_bready }),
    .m_axil_araddr({ m23_axil_araddr, m22_axil_araddr, m21_axil_araddr, m20_axil_araddr, m19_axil_araddr, m18_axil_araddr, m17_axil_araddr, m16_axil_araddr, m15_axil_araddr, m14_axil_araddr, m13_axil_araddr, m12_axil_araddr, m11_axil_araddr, m10_axil_araddr, m09_axil_araddr, m08_axil_araddr, m07_axil_araddr, m06_axil_araddr, m05_axil_araddr, m04_axil_araddr, m03_axil_araddr, m02_axil_araddr, m01_axil_araddr, m00_axil_araddr }),
    .m_axil_arprot({ m23_axil_arprot, m22_axil_arprot, m21_axil_arprot, m20_axil_arprot, m19_axil_arprot, m18_axil_arprot, m17_axil_arprot, m16_axil_arprot, m15_axil_arprot, m14_axil_arprot, m13_axil_arprot, m12_axil_arprot, m11_axil_arprot, m10_axil_arprot, m09_axil_arprot, m08_axil_arprot, m07_axil_arprot, m06_axil_arprot, m05_axil_arprot, m04_axil_arprot, m03_axil_arprot, m02_axil_arprot, m01_axil_arprot, m00_axil_arprot }),
    .m_axil_arvalid({ m23_axil_arvalid, m22_axil_arvalid, m21_axil_arvalid, m20_axil_arvalid, m19_axil_arvalid, m18_axil_arvalid, m17_axil_arvalid, m16_axil_arvalid, m15_axil_arvalid, m14_axil_arvalid, m13_axil_arvalid, m12_axil_arvalid, m11_axil_arvalid, m10_axil_arvalid, m09_axil_arvalid, m08_axil_arvalid, m07_axil_arvalid, m06_axil_arvalid, m05_axil_arvalid, m04_axil_arvalid, m03_axil_arvalid, m02_axil_arvalid, m01_axil_arvalid, m00_axil_arvalid }),
    .m_axil_arready({ m23_axil_arready, m22_axil_arready, m21_axil_arready, m20_axil_arready, m19_axil_arready, m18_axil_arready, m17_axil_arready, m16_axil_arready, m15_axil_arready, m14_axil_arready, m13_axil_arready, m12_axil_arready, m11_axil_arready, m10_axil_arready, m09_axil_arready, m08_axil_arready, m07_axil_arready, m06_axil_arready, m05_axil_arready, m04_axil_arready, m03_axil_arready, m02_axil_arready, m01_axil_arready, m00_axil_arready }),
    .m_axil_rdata({ m23_axil_rdata, m22_axil_rdata, m21_axil_rdata, m20_axil_rdata, m19_axil_rdata, m18_axil_rdata, m17_axil_rdata, m16_axil_rdata, m15_axil_rdata, m14_axil_rdata, m13_axil_rdata, m12_axil_rdata, m11_axil_rdata, m10_axil_rdata, m09_axil_rdata, m08_axil_rdata, m07_axil_rdata, m06_axil_rdata, m05_axil_rdata, m04_axil_rdata, m03_axil_rdata, m02_axil_rdata, m01_axil_rdata, m00_axil_rdata }),
    .m_axil_rresp({ m23_axil_rresp, m22_axil_rresp, m21_axil_rresp, m20_axil_rresp, m19_axil_rresp, m18_axil_rresp, m17_axil_rresp, m16_axil_rresp, m15_axil_rresp, m14_axil_rresp, m13_axil_rresp, m12_axil_rresp, m11_axil_rresp, m10_axil_rresp, m09_axil_rresp, m08_axil_rresp, m07_axil_rresp, m06_axil_rresp, m05_axil_rresp, m04_axil_rresp, m03_axil_rresp, m02_axil_rresp, m01_axil_rresp, m00_axil_rresp }),
    .m_axil_rvalid({ m23_axil_rvalid, m22_axil_rvalid, m21_axil_rvalid, m20_axil_rvalid, m19_axil_rvalid, m18_axil_rvalid, m17_axil_rvalid, m16_axil_rvalid, m15_axil_rvalid, m14_axil_rvalid, m13_axil_rvalid, m12_axil_rvalid, m11_axil_rvalid, m10_axil_rvalid, m09_axil_rvalid, m08_axil_rvalid, m07_axil_rvalid, m06_axil_rvalid, m05_axil_rvalid, m04_axil_rvalid, m03_axil_rvalid, m02_axil_rvalid, m01_axil_rvalid, m00_axil_rvalid }),
    .m_axil_rready({ m23_axil_rready, m22_axil_rready, m21_axil_rready, m20_axil_rready, m19_axil_rready, m18_axil_rready, m17_axil_rready, m16_axil_rready, m15_axil_rready, m14_axil_rready, m13_axil_rready, m12_axil_rready, m11_axil_rready, m10_axil_rready, m09_axil_rready, m08_axil_rready, m07_axil_rready, m06_axil_rready, m05_axil_rready, m04_axil_rready, m03_axil_rready, m02_axil_rready, m01_axil_rready, m00_axil_rready })
);

endmodule

`resetall
