`define complex_dsp
`define hard_mem
`include "../../../../../vtr_flow/benchmarks/system_verilog/koios_sv/deepfreeze.style3.sv"
