/*
 * Ultra wide range test
*/

`define WIDTH 256
`define operator xnor
`include "../.generic/range_any_width_binary_test.v"