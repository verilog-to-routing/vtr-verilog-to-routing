module simple_op(in,out);
    input  [`WIDTH-1:0] in;
    output [`WIDTH-1:0] out;

    assign out = in;
endmodule