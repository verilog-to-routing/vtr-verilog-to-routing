module top(input in, output reg out);
	always @(*)
		out <= in;
endmodule
