`define BINARY_OP(out,a,b) nand(out, a, b);
`include "../.generic/wire_test.v"